// Benchmark "adder" written by ABC on Wed Jul 17 17:31:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n149,
    new_n150, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n179, new_n180, new_n181,
    new_n182, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n323, new_n326,
    new_n327, new_n329, new_n331, new_n332, new_n333;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n08x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nand22aa1n03x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  norp02aa1n04x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  tech160nm_fiao0012aa1n02p5x5 g006(.a(new_n99), .b(new_n101), .c(new_n100), .o(new_n102));
  inv000aa1d42x5               g007(.a(\a[2] ), .o1(new_n103));
  inv000aa1d42x5               g008(.a(\b[1] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  tech160nm_fioaoi03aa1n03p5x5 g010(.a(new_n103), .b(new_n104), .c(new_n105), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n02x4               g012(.a(new_n107), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n108));
  oabi12aa1n06x5               g013(.a(new_n102), .b(new_n108), .c(new_n106), .out0(new_n109));
  xorc02aa1n12x5               g014(.a(\a[7] ), .b(\b[6] ), .out0(new_n110));
  tech160nm_fixorc02aa1n05x5   g015(.a(\a[6] ), .b(\b[5] ), .out0(new_n111));
  nanp02aa1n02x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  xorc02aa1n02x5               g017(.a(\a[5] ), .b(\b[4] ), .out0(new_n113));
  xorc02aa1n02x5               g018(.a(\a[8] ), .b(\b[7] ), .out0(new_n114));
  nano22aa1n03x7               g019(.a(new_n112), .b(new_n113), .c(new_n114), .out0(new_n115));
  oai022aa1n02x5               g020(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n116));
  aoi022aa1n02x5               g021(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n116), .b(new_n117), .o1(new_n118));
  oa0022aa1n06x5               g023(.a(\a[8] ), .b(\b[7] ), .c(\a[7] ), .d(\b[6] ), .o(new_n119));
  aoi022aa1n06x5               g024(.a(new_n118), .b(new_n119), .c(\b[7] ), .d(\a[8] ), .o1(new_n120));
  xorc02aa1n02x5               g025(.a(\a[9] ), .b(\b[8] ), .out0(new_n121));
  aoai13aa1n03x5               g026(.a(new_n121), .b(new_n120), .c(new_n115), .d(new_n109), .o1(new_n122));
  nor042aa1n04x5               g027(.a(\b[9] ), .b(\a[10] ), .o1(new_n123));
  nand42aa1n04x5               g028(.a(\b[9] ), .b(\a[10] ), .o1(new_n124));
  norb02aa1n12x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n125), .b(new_n122), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g031(.a(new_n125), .o1(new_n127));
  oai012aa1n12x5               g032(.a(new_n124), .b(new_n123), .c(new_n97), .o1(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n122), .d(new_n98), .o1(new_n129));
  nand02aa1n06x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor002aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  norb02aa1n02x5               g037(.a(new_n128), .b(new_n132), .out0(new_n133));
  aoai13aa1n03x5               g038(.a(new_n133), .b(new_n127), .c(new_n122), .d(new_n98), .o1(new_n134));
  aob012aa1n02x5               g039(.a(new_n134), .b(new_n129), .c(new_n132), .out0(\s[11] ));
  nor022aa1n12x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1d06x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanb02aa1n02x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n134), .c(new_n130), .out0(\s[12] ));
  nona23aa1n09x5               g044(.a(new_n130), .b(new_n137), .c(new_n136), .d(new_n131), .out0(new_n140));
  nano22aa1n02x4               g045(.a(new_n140), .b(new_n121), .c(new_n125), .out0(new_n141));
  aoai13aa1n06x5               g046(.a(new_n141), .b(new_n120), .c(new_n115), .d(new_n109), .o1(new_n142));
  aoi012aa1n06x5               g047(.a(new_n136), .b(new_n131), .c(new_n137), .o1(new_n143));
  oai012aa1n12x5               g048(.a(new_n143), .b(new_n140), .c(new_n128), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n144), .o1(new_n145));
  nanp02aa1n02x5               g050(.a(new_n142), .b(new_n145), .o1(new_n146));
  xorb03aa1n02x5               g051(.a(new_n146), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g052(.a(\a[13] ), .o1(new_n148));
  inv000aa1d42x5               g053(.a(\b[12] ), .o1(new_n149));
  oaoi03aa1n02x5               g054(.a(new_n148), .b(new_n149), .c(new_n146), .o1(new_n150));
  xnrb03aa1n03x5               g055(.a(new_n150), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nand42aa1n08x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nor022aa1n04x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nor042aa1n04x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nand42aa1n06x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nona23aa1n06x5               g060(.a(new_n152), .b(new_n155), .c(new_n154), .d(new_n153), .out0(new_n156));
  aoai13aa1n02x5               g061(.a(new_n155), .b(new_n154), .c(new_n148), .d(new_n149), .o1(new_n157));
  aoai13aa1n04x5               g062(.a(new_n157), .b(new_n156), .c(new_n142), .d(new_n145), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand42aa1n06x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nor042aa1n03x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nor042aa1n02x5               g066(.a(\b[15] ), .b(\a[16] ), .o1(new_n162));
  nand02aa1n06x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n161), .c(new_n158), .d(new_n160), .o1(new_n165));
  aoi112aa1n02x7               g070(.a(new_n164), .b(new_n161), .c(new_n158), .d(new_n160), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(\s[16] ));
  nano23aa1n03x7               g072(.a(new_n136), .b(new_n131), .c(new_n137), .d(new_n130), .out0(new_n168));
  nano23aa1n06x5               g073(.a(new_n154), .b(new_n153), .c(new_n155), .d(new_n152), .out0(new_n169));
  nano23aa1n09x5               g074(.a(new_n162), .b(new_n161), .c(new_n163), .d(new_n160), .out0(new_n170));
  nand22aa1n03x5               g075(.a(new_n170), .b(new_n169), .o1(new_n171));
  nano32aa1n03x7               g076(.a(new_n171), .b(new_n168), .c(new_n125), .d(new_n121), .out0(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n120), .c(new_n115), .d(new_n109), .o1(new_n173));
  inv000aa1n02x5               g078(.a(new_n157), .o1(new_n174));
  aoai13aa1n06x5               g079(.a(new_n170), .b(new_n174), .c(new_n144), .d(new_n169), .o1(new_n175));
  tech160nm_fiaoi012aa1n04x5   g080(.a(new_n162), .b(new_n161), .c(new_n163), .o1(new_n176));
  nand23aa1n06x5               g081(.a(new_n173), .b(new_n175), .c(new_n176), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g083(.a(\a[18] ), .o1(new_n179));
  inv040aa1d32x5               g084(.a(\a[17] ), .o1(new_n180));
  inv030aa1d32x5               g085(.a(\b[16] ), .o1(new_n181));
  oaoi03aa1n03x5               g086(.a(new_n180), .b(new_n181), .c(new_n177), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[17] ), .c(new_n179), .out0(\s[18] ));
  oaoi13aa1n04x5               g088(.a(new_n156), .b(new_n143), .c(new_n140), .d(new_n128), .o1(new_n184));
  inv000aa1n02x5               g089(.a(new_n176), .o1(new_n185));
  oaoi13aa1n09x5               g090(.a(new_n185), .b(new_n170), .c(new_n184), .d(new_n174), .o1(new_n186));
  xroi22aa1d06x4               g091(.a(new_n180), .b(\b[16] ), .c(new_n179), .d(\b[17] ), .out0(new_n187));
  inv000aa1n02x5               g092(.a(new_n187), .o1(new_n188));
  oai022aa1n02x5               g093(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n189));
  oaib12aa1n02x5               g094(.a(new_n189), .b(new_n179), .c(\b[17] ), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n188), .c(new_n186), .d(new_n173), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g097(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n12x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand42aa1d28x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nanb02aa1n02x5               g100(.a(new_n194), .b(new_n195), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  nor042aa1n06x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nand42aa1d28x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  aoai13aa1n02x5               g105(.a(new_n200), .b(new_n194), .c(new_n191), .d(new_n197), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(new_n181), .b(new_n180), .o1(new_n202));
  oaoi03aa1n09x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n197), .b(new_n203), .c(new_n177), .d(new_n187), .o1(new_n204));
  nona22aa1n03x5               g109(.a(new_n204), .b(new_n200), .c(new_n194), .out0(new_n205));
  nanp02aa1n03x5               g110(.a(new_n201), .b(new_n205), .o1(\s[20] ));
  nano23aa1d15x5               g111(.a(new_n198), .b(new_n194), .c(new_n199), .d(new_n195), .out0(new_n207));
  nand22aa1n12x5               g112(.a(new_n187), .b(new_n207), .o1(new_n208));
  nona23aa1n02x4               g113(.a(new_n195), .b(new_n199), .c(new_n198), .d(new_n194), .out0(new_n209));
  tech160nm_fiaoi012aa1n03p5x5 g114(.a(new_n198), .b(new_n194), .c(new_n199), .o1(new_n210));
  oai012aa1n02x5               g115(.a(new_n210), .b(new_n209), .c(new_n190), .o1(new_n211));
  inv000aa1n02x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n02x7               g117(.a(new_n212), .b(new_n208), .c(new_n186), .d(new_n173), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  xnrc02aa1n12x5               g120(.a(\b[20] ), .b(\a[21] ), .out0(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  tech160nm_fixnrc02aa1n04x5   g122(.a(\b[21] ), .b(\a[22] ), .out0(new_n218));
  aoai13aa1n02x5               g123(.a(new_n218), .b(new_n215), .c(new_n213), .d(new_n217), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n208), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n217), .b(new_n211), .c(new_n177), .d(new_n220), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n218), .c(new_n215), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n219), .b(new_n222), .o1(\s[22] ));
  oao003aa1n02x5               g128(.a(new_n103), .b(new_n104), .c(new_n105), .carry(new_n224));
  nano23aa1n02x4               g129(.a(new_n99), .b(new_n101), .c(new_n107), .d(new_n100), .out0(new_n225));
  aoi012aa1n02x5               g130(.a(new_n102), .b(new_n225), .c(new_n224), .o1(new_n226));
  xnrc02aa1n02x5               g131(.a(\b[6] ), .b(\a[7] ), .out0(new_n227));
  xnrc02aa1n02x5               g132(.a(\b[7] ), .b(\a[8] ), .out0(new_n228));
  nona23aa1n02x4               g133(.a(new_n113), .b(new_n111), .c(new_n228), .d(new_n227), .out0(new_n229));
  inv000aa1n02x5               g134(.a(new_n120), .o1(new_n230));
  tech160nm_fioai012aa1n03p5x5 g135(.a(new_n230), .b(new_n229), .c(new_n226), .o1(new_n231));
  nona23aa1n02x4               g136(.a(new_n160), .b(new_n163), .c(new_n162), .d(new_n161), .out0(new_n232));
  inv040aa1n03x5               g137(.a(new_n128), .o1(new_n233));
  inv020aa1n02x5               g138(.a(new_n143), .o1(new_n234));
  aoai13aa1n02x7               g139(.a(new_n169), .b(new_n234), .c(new_n168), .d(new_n233), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n176), .b(new_n232), .c(new_n235), .d(new_n157), .o1(new_n236));
  nor042aa1n06x5               g141(.a(new_n218), .b(new_n216), .o1(new_n237));
  nano22aa1n02x4               g142(.a(new_n188), .b(new_n237), .c(new_n207), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n236), .c(new_n231), .d(new_n172), .o1(new_n239));
  inv030aa1n03x5               g144(.a(new_n210), .o1(new_n240));
  aoai13aa1n12x5               g145(.a(new_n237), .b(new_n240), .c(new_n207), .d(new_n203), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  inv000aa1d42x5               g147(.a(\a[22] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(\b[21] ), .o1(new_n244));
  oaoi03aa1n12x5               g149(.a(new_n243), .b(new_n244), .c(new_n215), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  nona22aa1n02x5               g151(.a(new_n239), .b(new_n242), .c(new_n246), .out0(new_n247));
  nor042aa1n03x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  and002aa1n12x5               g153(.a(\b[22] ), .b(\a[23] ), .o(new_n249));
  nor042aa1n03x5               g154(.a(new_n249), .b(new_n248), .o1(new_n250));
  nona32aa1n02x4               g155(.a(new_n239), .b(new_n250), .c(new_n246), .d(new_n242), .out0(new_n251));
  aobi12aa1n02x5               g156(.a(new_n251), .b(new_n250), .c(new_n247), .out0(\s[23] ));
  norb02aa1n02x5               g157(.a(new_n245), .b(new_n248), .out0(new_n253));
  aoi013aa1n02x4               g158(.a(new_n249), .b(new_n239), .c(new_n241), .d(new_n253), .o1(new_n254));
  tech160nm_fixnrc02aa1n05x5   g159(.a(\b[23] ), .b(\a[24] ), .out0(new_n255));
  nona32aa1n02x5               g160(.a(new_n239), .b(new_n248), .c(new_n246), .d(new_n242), .out0(new_n256));
  nanb03aa1n03x5               g161(.a(new_n249), .b(new_n256), .c(new_n255), .out0(new_n257));
  oai012aa1n03x5               g162(.a(new_n257), .b(new_n254), .c(new_n255), .o1(\s[24] ));
  norb02aa1n02x5               g163(.a(new_n250), .b(new_n255), .out0(new_n259));
  nano22aa1n03x7               g164(.a(new_n208), .b(new_n237), .c(new_n259), .out0(new_n260));
  inv020aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n259), .o1(new_n262));
  orn002aa1n02x5               g167(.a(\a[23] ), .b(\b[22] ), .o(new_n263));
  oao003aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .c(new_n263), .carry(new_n264));
  aoai13aa1n12x5               g169(.a(new_n264), .b(new_n262), .c(new_n241), .d(new_n245), .o1(new_n265));
  inv020aa1n03x5               g170(.a(new_n265), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n266), .b(new_n261), .c(new_n186), .d(new_n173), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  tech160nm_fixorc02aa1n03p5x5 g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[25] ), .b(\a[26] ), .out0(new_n271));
  aoai13aa1n03x5               g176(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n270), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n270), .b(new_n265), .c(new_n177), .d(new_n260), .o1(new_n273));
  nona22aa1n02x5               g178(.a(new_n273), .b(new_n271), .c(new_n269), .out0(new_n274));
  nanp02aa1n03x5               g179(.a(new_n272), .b(new_n274), .o1(\s[26] ));
  nor042aa1n04x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  and002aa1n18x5               g181(.a(\b[26] ), .b(\a[27] ), .o(new_n277));
  norp02aa1n06x5               g182(.a(new_n277), .b(new_n276), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n270), .b(new_n271), .out0(new_n279));
  nano32aa1n06x5               g184(.a(new_n208), .b(new_n279), .c(new_n237), .d(new_n259), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n236), .c(new_n231), .d(new_n172), .o1(new_n281));
  orn002aa1n02x5               g186(.a(\a[25] ), .b(\b[24] ), .o(new_n282));
  oao003aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .c(new_n282), .carry(new_n283));
  aobi12aa1n06x5               g188(.a(new_n283), .b(new_n265), .c(new_n279), .out0(new_n284));
  xnbna2aa1n06x5               g189(.a(new_n278), .b(new_n281), .c(new_n284), .out0(\s[27] ));
  inv000aa1d42x5               g190(.a(new_n277), .o1(new_n286));
  nanp02aa1n03x5               g191(.a(new_n265), .b(new_n279), .o1(new_n287));
  tech160nm_finand02aa1n03p5x5 g192(.a(new_n287), .b(new_n283), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n286), .b(new_n288), .c(new_n177), .d(new_n280), .o1(new_n289));
  xorc02aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .out0(new_n290));
  norp02aa1n02x5               g195(.a(new_n290), .b(new_n276), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n276), .o1(new_n292));
  aoai13aa1n02x7               g197(.a(new_n292), .b(new_n277), .c(new_n281), .d(new_n284), .o1(new_n293));
  aoi022aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n289), .d(new_n291), .o1(\s[28] ));
  and002aa1n06x5               g199(.a(new_n290), .b(new_n278), .o(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n288), .c(new_n177), .d(new_n280), .o1(new_n296));
  inv000aa1n02x5               g201(.a(new_n295), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .carry(new_n298));
  aoai13aa1n02x7               g203(.a(new_n298), .b(new_n297), .c(new_n281), .d(new_n284), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n298), .b(new_n300), .out0(new_n301));
  aoi022aa1n03x5               g206(.a(new_n299), .b(new_n300), .c(new_n296), .d(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g208(.a(new_n290), .b(new_n300), .c(new_n278), .o(new_n304));
  aoai13aa1n06x5               g209(.a(new_n304), .b(new_n288), .c(new_n177), .d(new_n280), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n307));
  aoai13aa1n02x7               g212(.a(new_n307), .b(new_n306), .c(new_n281), .d(new_n284), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n307), .b(new_n309), .out0(new_n310));
  aoi022aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n305), .d(new_n310), .o1(\s[30] ));
  nano22aa1n06x5               g216(.a(new_n297), .b(new_n300), .c(new_n309), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n288), .c(new_n177), .d(new_n280), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n312), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n315));
  aoai13aa1n02x7               g220(.a(new_n315), .b(new_n314), .c(new_n281), .d(new_n284), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[31] ), .b(\b[30] ), .out0(new_n317));
  and002aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .o(new_n318));
  oabi12aa1n02x5               g223(.a(new_n317), .b(\a[30] ), .c(\b[29] ), .out0(new_n319));
  oab012aa1n02x4               g224(.a(new_n319), .b(new_n307), .c(new_n318), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n316), .b(new_n317), .c(new_n313), .d(new_n320), .o1(\s[31] ));
  xnrb03aa1n02x5               g226(.a(new_n106), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g227(.a(\a[3] ), .b(\b[2] ), .c(new_n106), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g229(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanp02aa1n02x5               g230(.a(\b[4] ), .b(\a[5] ), .o1(new_n326));
  oaib12aa1n06x5               g231(.a(new_n326), .b(new_n109), .c(new_n113), .out0(new_n327));
  xnrc02aa1n02x5               g232(.a(new_n327), .b(new_n111), .out0(\s[6] ));
  oao003aa1n03x5               g233(.a(\a[6] ), .b(\b[5] ), .c(new_n327), .carry(new_n329));
  xnrc02aa1n02x5               g234(.a(new_n329), .b(new_n110), .out0(\s[7] ));
  and002aa1n02x5               g235(.a(\b[6] ), .b(\a[7] ), .o(new_n331));
  aoai13aa1n03x5               g236(.a(new_n228), .b(new_n331), .c(new_n329), .d(new_n110), .o1(new_n332));
  aoi112aa1n02x5               g237(.a(new_n228), .b(new_n331), .c(new_n329), .d(new_n110), .o1(new_n333));
  norb02aa1n03x4               g238(.a(new_n332), .b(new_n333), .out0(\s[8] ));
  xorb03aa1n02x5               g239(.a(new_n231), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


