// Benchmark "adder" written by ABC on Wed Jul 17 14:51:38 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n156, new_n157, new_n158, new_n159, new_n160, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n355, new_n356, new_n358, new_n359,
    new_n362, new_n363, new_n366, new_n368, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1n16x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  aob012aa1n06x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .out0(new_n107));
  nor042aa1n03x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand42aa1n03x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nano23aa1n03x5               g016(.a(new_n108), .b(new_n110), .c(new_n111), .d(new_n109), .out0(new_n112));
  nand42aa1n02x5               g017(.a(new_n112), .b(new_n107), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\a[3] ), .o1(new_n114));
  inv000aa1d42x5               g019(.a(\b[2] ), .o1(new_n115));
  aoai13aa1n03x5               g020(.a(new_n109), .b(new_n108), .c(new_n114), .d(new_n115), .o1(new_n116));
  nand02aa1n04x5               g021(.a(new_n113), .b(new_n116), .o1(new_n117));
  norp02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanp02aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  norb02aa1n02x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  norp02aa1n04x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nand42aa1n06x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  norb02aa1n02x7               g027(.a(new_n122), .b(new_n121), .out0(new_n123));
  xorc02aa1n12x5               g028(.a(\a[8] ), .b(\b[7] ), .out0(new_n124));
  inv000aa1d42x5               g029(.a(new_n124), .o1(new_n125));
  nor042aa1n03x5               g030(.a(\b[6] ), .b(\a[7] ), .o1(new_n126));
  nand42aa1n03x5               g031(.a(\b[6] ), .b(\a[7] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  nano32aa1n03x7               g033(.a(new_n125), .b(new_n128), .c(new_n120), .d(new_n123), .out0(new_n129));
  nona22aa1n06x5               g034(.a(new_n119), .b(new_n121), .c(new_n118), .out0(new_n130));
  nano22aa1n03x7               g035(.a(new_n126), .b(new_n119), .c(new_n127), .out0(new_n131));
  nanp03aa1n02x5               g036(.a(new_n130), .b(new_n131), .c(new_n124), .o1(new_n132));
  inv000aa1n03x5               g037(.a(new_n126), .o1(new_n133));
  oao003aa1n09x5               g038(.a(\a[8] ), .b(\b[7] ), .c(new_n133), .carry(new_n134));
  nand22aa1n02x5               g039(.a(new_n132), .b(new_n134), .o1(new_n135));
  nand42aa1n02x5               g040(.a(\b[8] ), .b(\a[9] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n100), .out0(new_n137));
  aoai13aa1n02x5               g042(.a(new_n137), .b(new_n135), .c(new_n117), .d(new_n129), .o1(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n99), .b(new_n138), .c(new_n101), .out0(\s[10] ));
  aobi12aa1n02x5               g044(.a(new_n116), .b(new_n112), .c(new_n107), .out0(new_n140));
  nano23aa1n02x4               g045(.a(new_n118), .b(new_n121), .c(new_n122), .d(new_n119), .out0(new_n141));
  nand23aa1n03x5               g046(.a(new_n141), .b(new_n124), .c(new_n128), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n134), .o1(new_n143));
  aoi013aa1n06x4               g048(.a(new_n143), .b(new_n131), .c(new_n130), .d(new_n124), .o1(new_n144));
  oai012aa1n02x5               g049(.a(new_n144), .b(new_n140), .c(new_n142), .o1(new_n145));
  nona23aa1d18x5               g050(.a(new_n136), .b(new_n98), .c(new_n97), .d(new_n100), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  aoi012aa1d24x5               g052(.a(new_n97), .b(new_n100), .c(new_n98), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nor002aa1d24x5               g054(.a(\b[10] ), .b(\a[11] ), .o1(new_n150));
  nand02aa1n03x5               g055(.a(\b[10] ), .b(\a[11] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n149), .c(new_n145), .d(new_n147), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n152), .b(new_n149), .c(new_n145), .d(new_n147), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(\s[11] ));
  inv040aa1n03x5               g060(.a(new_n150), .o1(new_n156));
  norp02aa1n04x5               g061(.a(\b[11] ), .b(\a[12] ), .o1(new_n157));
  nand42aa1n02x5               g062(.a(\b[11] ), .b(\a[12] ), .o1(new_n158));
  norb02aa1n02x5               g063(.a(new_n158), .b(new_n157), .out0(new_n159));
  nona23aa1n02x4               g064(.a(new_n153), .b(new_n158), .c(new_n157), .d(new_n150), .out0(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n159), .c(new_n156), .d(new_n153), .o1(\s[12] ));
  nona23aa1d18x5               g066(.a(new_n158), .b(new_n151), .c(new_n150), .d(new_n157), .out0(new_n162));
  nor042aa1n03x5               g067(.a(new_n162), .b(new_n146), .o1(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n135), .c(new_n117), .d(new_n129), .o1(new_n164));
  tech160nm_fioaoi03aa1n03p5x5 g069(.a(\a[12] ), .b(\b[11] ), .c(new_n156), .o1(new_n165));
  oabi12aa1n18x5               g070(.a(new_n165), .b(new_n162), .c(new_n148), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  nand42aa1n04x5               g072(.a(new_n164), .b(new_n167), .o1(new_n168));
  norp02aa1n04x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nand42aa1n03x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  nanb02aa1n12x5               g075(.a(new_n169), .b(new_n170), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  nano23aa1n06x5               g077(.a(new_n150), .b(new_n157), .c(new_n158), .d(new_n151), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(new_n165), .b(new_n172), .c(new_n173), .d(new_n149), .o1(new_n174));
  aoi022aa1n02x5               g079(.a(new_n168), .b(new_n172), .c(new_n164), .d(new_n174), .o1(\s[13] ));
  nor042aa1n02x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  nand42aa1n03x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n169), .c(new_n168), .d(new_n170), .o1(new_n179));
  nona22aa1n02x4               g084(.a(new_n177), .b(new_n176), .c(new_n169), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n179), .b(new_n180), .c(new_n172), .d(new_n168), .o1(\s[14] ));
  nano23aa1n09x5               g086(.a(new_n169), .b(new_n176), .c(new_n177), .d(new_n170), .out0(new_n182));
  tech160nm_fiaoi012aa1n04x5   g087(.a(new_n176), .b(new_n169), .c(new_n177), .o1(new_n183));
  inv000aa1n02x5               g088(.a(new_n183), .o1(new_n184));
  nor002aa1n06x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nanp02aa1n02x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  nanb02aa1n02x5               g091(.a(new_n185), .b(new_n186), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  aoai13aa1n03x5               g093(.a(new_n188), .b(new_n184), .c(new_n168), .d(new_n182), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(new_n188), .b(new_n184), .c(new_n168), .d(new_n182), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n189), .b(new_n190), .out0(\s[15] ));
  inv000aa1d42x5               g096(.a(new_n185), .o1(new_n192));
  nor002aa1n02x5               g097(.a(\b[15] ), .b(\a[16] ), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(\b[15] ), .b(\a[16] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  norb03aa1n02x5               g101(.a(new_n194), .b(new_n185), .c(new_n193), .out0(new_n197));
  nand02aa1n03x5               g102(.a(new_n189), .b(new_n197), .o1(new_n198));
  aoai13aa1n02x5               g103(.a(new_n198), .b(new_n196), .c(new_n192), .d(new_n189), .o1(\s[16] ));
  nano23aa1n06x5               g104(.a(new_n185), .b(new_n193), .c(new_n194), .d(new_n186), .out0(new_n200));
  nano32aa1n03x7               g105(.a(new_n146), .b(new_n200), .c(new_n173), .d(new_n182), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n135), .c(new_n117), .d(new_n129), .o1(new_n202));
  aoai13aa1n12x5               g107(.a(new_n200), .b(new_n184), .c(new_n166), .d(new_n182), .o1(new_n203));
  oai012aa1n02x5               g108(.a(new_n194), .b(new_n193), .c(new_n185), .o1(new_n204));
  nanp03aa1d12x5               g109(.a(new_n202), .b(new_n203), .c(new_n204), .o1(new_n205));
  tech160nm_fixorc02aa1n04x5   g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  nano22aa1n02x4               g111(.a(new_n206), .b(new_n203), .c(new_n204), .out0(new_n207));
  aoi022aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n205), .d(new_n206), .o1(\s[17] ));
  nor042aa1d18x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nona23aa1n09x5               g115(.a(new_n194), .b(new_n186), .c(new_n185), .d(new_n193), .out0(new_n211));
  nona32aa1n03x5               g116(.a(new_n163), .b(new_n211), .c(new_n178), .d(new_n171), .out0(new_n212));
  oaoi13aa1n09x5               g117(.a(new_n212), .b(new_n144), .c(new_n140), .d(new_n142), .o1(new_n213));
  aoai13aa1n06x5               g118(.a(new_n182), .b(new_n165), .c(new_n173), .d(new_n149), .o1(new_n214));
  aoai13aa1n06x5               g119(.a(new_n204), .b(new_n211), .c(new_n214), .d(new_n183), .o1(new_n215));
  oaih12aa1n02x5               g120(.a(new_n206), .b(new_n215), .c(new_n213), .o1(new_n216));
  nor042aa1n06x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  nand02aa1d12x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  norb02aa1n06x4               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  nona23aa1n02x4               g124(.a(new_n216), .b(new_n218), .c(new_n217), .d(new_n209), .out0(new_n220));
  aoai13aa1n02x5               g125(.a(new_n220), .b(new_n219), .c(new_n210), .d(new_n216), .o1(\s[18] ));
  and002aa1n02x5               g126(.a(new_n206), .b(new_n219), .o(new_n222));
  oaih12aa1n02x5               g127(.a(new_n222), .b(new_n215), .c(new_n213), .o1(new_n223));
  aoi012aa1d24x5               g128(.a(new_n217), .b(new_n209), .c(new_n218), .o1(new_n224));
  nor042aa1n06x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  nand22aa1n04x5               g130(.a(\b[18] ), .b(\a[19] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  xnbna2aa1n03x5               g132(.a(new_n227), .b(new_n223), .c(new_n224), .out0(\s[19] ));
  xnrc02aa1n02x5               g133(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g134(.a(new_n225), .o1(new_n230));
  inv030aa1n06x5               g135(.a(new_n224), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n227), .b(new_n231), .c(new_n205), .d(new_n222), .o1(new_n232));
  nor022aa1n06x5               g137(.a(\b[19] ), .b(\a[20] ), .o1(new_n233));
  nand22aa1n04x5               g138(.a(\b[19] ), .b(\a[20] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n227), .o1(new_n236));
  norb03aa1n02x5               g141(.a(new_n234), .b(new_n225), .c(new_n233), .out0(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n236), .c(new_n223), .d(new_n224), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n235), .c(new_n232), .d(new_n230), .o1(\s[20] ));
  nona23aa1d18x5               g144(.a(new_n234), .b(new_n226), .c(new_n225), .d(new_n233), .out0(new_n240));
  nano22aa1d15x5               g145(.a(new_n240), .b(new_n206), .c(new_n219), .out0(new_n241));
  tech160nm_fioai012aa1n04x5   g146(.a(new_n241), .b(new_n215), .c(new_n213), .o1(new_n242));
  oaoi03aa1n12x5               g147(.a(\a[20] ), .b(\b[19] ), .c(new_n230), .o1(new_n243));
  inv030aa1n02x5               g148(.a(new_n243), .o1(new_n244));
  oai012aa1d24x5               g149(.a(new_n244), .b(new_n240), .c(new_n224), .o1(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[20] ), .b(\a[21] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n245), .c(new_n205), .d(new_n241), .o1(new_n248));
  nano23aa1n06x5               g153(.a(new_n225), .b(new_n233), .c(new_n234), .d(new_n226), .out0(new_n249));
  aoi112aa1n02x5               g154(.a(new_n243), .b(new_n247), .c(new_n249), .d(new_n231), .o1(new_n250));
  aobi12aa1n03x7               g155(.a(new_n248), .b(new_n250), .c(new_n242), .out0(\s[21] ));
  nor042aa1n06x5               g156(.a(\b[20] ), .b(\a[21] ), .o1(new_n252));
  inv020aa1n04x5               g157(.a(new_n252), .o1(new_n253));
  xnrc02aa1n12x5               g158(.a(\b[21] ), .b(\a[22] ), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n245), .o1(new_n256));
  oai022aa1n02x5               g161(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n257));
  aoi012aa1n02x5               g162(.a(new_n257), .b(\a[22] ), .c(\b[21] ), .o1(new_n258));
  aoai13aa1n02x7               g163(.a(new_n258), .b(new_n246), .c(new_n242), .d(new_n256), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n255), .c(new_n248), .d(new_n253), .o1(\s[22] ));
  nor042aa1n06x5               g165(.a(new_n254), .b(new_n246), .o1(new_n261));
  nano32aa1n02x4               g166(.a(new_n240), .b(new_n261), .c(new_n206), .d(new_n219), .out0(new_n262));
  oaih12aa1n02x5               g167(.a(new_n262), .b(new_n215), .c(new_n213), .o1(new_n263));
  aoai13aa1n09x5               g168(.a(new_n261), .b(new_n243), .c(new_n249), .d(new_n231), .o1(new_n264));
  oaoi03aa1n02x5               g169(.a(\a[22] ), .b(\b[21] ), .c(new_n253), .o1(new_n265));
  inv000aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  nand22aa1n03x5               g171(.a(new_n264), .b(new_n266), .o1(new_n267));
  xorc02aa1n12x5               g172(.a(\a[23] ), .b(\b[22] ), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n267), .c(new_n205), .d(new_n262), .o1(new_n269));
  aoi112aa1n02x5               g174(.a(new_n268), .b(new_n265), .c(new_n245), .d(new_n261), .o1(new_n270));
  aobi12aa1n03x7               g175(.a(new_n269), .b(new_n270), .c(new_n263), .out0(\s[23] ));
  norp02aa1n02x5               g176(.a(\b[22] ), .b(\a[23] ), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[24] ), .b(\b[23] ), .out0(new_n274));
  inv000aa1d42x5               g179(.a(new_n267), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n268), .o1(new_n276));
  oai022aa1n02x5               g181(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n277));
  aoi012aa1n02x5               g182(.a(new_n277), .b(\a[24] ), .c(\b[23] ), .o1(new_n278));
  aoai13aa1n02x7               g183(.a(new_n278), .b(new_n276), .c(new_n263), .d(new_n275), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n274), .c(new_n269), .d(new_n273), .o1(\s[24] ));
  inv000aa1d42x5               g185(.a(new_n241), .o1(new_n281));
  and002aa1n02x7               g186(.a(new_n274), .b(new_n268), .o(new_n282));
  nano22aa1n02x4               g187(.a(new_n281), .b(new_n282), .c(new_n261), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n283), .b(new_n215), .c(new_n213), .o1(new_n284));
  inv000aa1n03x5               g189(.a(new_n282), .o1(new_n285));
  aob012aa1n02x5               g190(.a(new_n277), .b(\b[23] ), .c(\a[24] ), .out0(new_n286));
  aoai13aa1n12x5               g191(.a(new_n286), .b(new_n285), .c(new_n264), .d(new_n266), .o1(new_n287));
  xorc02aa1n12x5               g192(.a(\a[25] ), .b(\b[24] ), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n287), .c(new_n205), .d(new_n283), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n282), .b(new_n265), .c(new_n245), .d(new_n261), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n288), .o1(new_n291));
  and003aa1n02x5               g196(.a(new_n290), .b(new_n291), .c(new_n286), .o(new_n292));
  aobi12aa1n03x7               g197(.a(new_n289), .b(new_n292), .c(new_n284), .out0(\s[25] ));
  norp02aa1n02x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[26] ), .b(\b[25] ), .out0(new_n296));
  inv000aa1d42x5               g201(.a(new_n287), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(\b[25] ), .b(\a[26] ), .o1(new_n298));
  oai022aa1n02x5               g203(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n299));
  norb02aa1n02x5               g204(.a(new_n298), .b(new_n299), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n291), .c(new_n284), .d(new_n297), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n296), .c(new_n289), .d(new_n295), .o1(\s[26] ));
  and002aa1n02x5               g207(.a(new_n296), .b(new_n288), .o(new_n303));
  inv000aa1n02x5               g208(.a(new_n303), .o1(new_n304));
  nano32aa1n03x7               g209(.a(new_n304), .b(new_n241), .c(new_n282), .d(new_n261), .out0(new_n305));
  oai012aa1n06x5               g210(.a(new_n305), .b(new_n215), .c(new_n213), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(new_n299), .b(new_n298), .o1(new_n307));
  aoai13aa1n04x5               g212(.a(new_n307), .b(new_n304), .c(new_n290), .d(new_n286), .o1(new_n308));
  tech160nm_fixorc02aa1n03p5x5 g213(.a(\a[27] ), .b(\b[26] ), .out0(new_n309));
  aoai13aa1n06x5               g214(.a(new_n309), .b(new_n308), .c(new_n205), .d(new_n305), .o1(new_n310));
  aoi122aa1n02x5               g215(.a(new_n309), .b(new_n298), .c(new_n299), .d(new_n287), .e(new_n303), .o1(new_n311));
  aobi12aa1n03x7               g216(.a(new_n310), .b(new_n311), .c(new_n306), .out0(\s[27] ));
  nor042aa1n02x5               g217(.a(\b[26] ), .b(\a[27] ), .o1(new_n313));
  inv020aa1n02x5               g218(.a(new_n313), .o1(new_n314));
  nor002aa1n03x5               g219(.a(\b[27] ), .b(\a[28] ), .o1(new_n315));
  and002aa1n03x5               g220(.a(\b[27] ), .b(\a[28] ), .o(new_n316));
  nor042aa1n03x5               g221(.a(new_n316), .b(new_n315), .o1(new_n317));
  aoi022aa1n12x5               g222(.a(new_n287), .b(new_n303), .c(new_n298), .d(new_n299), .o1(new_n318));
  inv000aa1n02x5               g223(.a(new_n309), .o1(new_n319));
  norp03aa1n02x5               g224(.a(new_n316), .b(new_n315), .c(new_n313), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n306), .d(new_n318), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n310), .d(new_n314), .o1(\s[28] ));
  and002aa1n02x5               g227(.a(new_n309), .b(new_n317), .o(new_n323));
  aoai13aa1n06x5               g228(.a(new_n323), .b(new_n308), .c(new_n205), .d(new_n305), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  oab012aa1n06x5               g230(.a(new_n315), .b(new_n314), .c(new_n316), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n325), .c(new_n306), .d(new_n318), .o1(new_n327));
  tech160nm_fixorc02aa1n03p5x5 g232(.a(\a[29] ), .b(\b[28] ), .out0(new_n328));
  norb02aa1n02x5               g233(.a(new_n326), .b(new_n328), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n324), .d(new_n329), .o1(\s[29] ));
  xorb03aa1n02x5               g235(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g236(.a(new_n319), .b(new_n328), .c(new_n317), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n308), .c(new_n205), .d(new_n305), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n332), .o1(new_n334));
  tech160nm_fioaoi03aa1n02p5x5 g239(.a(\a[29] ), .b(\b[28] ), .c(new_n326), .o1(new_n335));
  inv000aa1d42x5               g240(.a(new_n335), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n334), .c(new_n306), .d(new_n318), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[30] ), .b(\b[29] ), .out0(new_n338));
  and002aa1n02x5               g243(.a(\b[28] ), .b(\a[29] ), .o(new_n339));
  oabi12aa1n02x5               g244(.a(new_n338), .b(\a[29] ), .c(\b[28] ), .out0(new_n340));
  oab012aa1n02x4               g245(.a(new_n340), .b(new_n326), .c(new_n339), .out0(new_n341));
  aoi022aa1n02x7               g246(.a(new_n337), .b(new_n338), .c(new_n333), .d(new_n341), .o1(\s[30] ));
  nano32aa1n02x4               g247(.a(new_n319), .b(new_n338), .c(new_n317), .d(new_n328), .out0(new_n343));
  aoai13aa1n06x5               g248(.a(new_n343), .b(new_n308), .c(new_n205), .d(new_n305), .o1(new_n344));
  inv000aa1n02x5               g249(.a(new_n343), .o1(new_n345));
  inv000aa1d42x5               g250(.a(\a[30] ), .o1(new_n346));
  inv000aa1d42x5               g251(.a(\b[29] ), .o1(new_n347));
  oaoi03aa1n02x5               g252(.a(new_n346), .b(new_n347), .c(new_n335), .o1(new_n348));
  aoai13aa1n03x5               g253(.a(new_n348), .b(new_n345), .c(new_n306), .d(new_n318), .o1(new_n349));
  xorc02aa1n02x5               g254(.a(\a[31] ), .b(\b[30] ), .out0(new_n350));
  oabi12aa1n02x5               g255(.a(new_n350), .b(\a[30] ), .c(\b[29] ), .out0(new_n351));
  oaoi13aa1n02x5               g256(.a(new_n351), .b(new_n335), .c(new_n346), .d(new_n347), .o1(new_n352));
  aoi022aa1n02x7               g257(.a(new_n349), .b(new_n350), .c(new_n344), .d(new_n352), .o1(\s[31] ));
  nanp03aa1n02x5               g258(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n354));
  nanb02aa1n02x5               g259(.a(new_n110), .b(new_n111), .out0(new_n355));
  inv000aa1d42x5               g260(.a(new_n355), .o1(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n356), .b(new_n354), .c(new_n104), .out0(\s[3] ));
  obai22aa1n02x7               g262(.a(new_n109), .b(new_n108), .c(\a[3] ), .d(\b[2] ), .out0(new_n358));
  aoi012aa1n02x5               g263(.a(new_n358), .b(new_n356), .c(new_n107), .o1(new_n359));
  oaoi13aa1n02x5               g264(.a(new_n359), .b(new_n117), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g265(.a(new_n123), .b(new_n113), .c(new_n116), .out0(\s[5] ));
  aoi012aa1n02x5               g266(.a(new_n121), .b(new_n117), .c(new_n122), .o1(new_n362));
  tech160nm_fiao0012aa1n02p5x5 g267(.a(new_n130), .b(new_n117), .c(new_n123), .o(new_n363));
  oai012aa1n02x5               g268(.a(new_n363), .b(new_n362), .c(new_n120), .o1(\s[6] ));
  xobna2aa1n03x5               g269(.a(new_n128), .b(new_n363), .c(new_n119), .out0(\s[7] ));
  aoai13aa1n02x5               g270(.a(new_n131), .b(new_n130), .c(new_n117), .d(new_n123), .o1(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n124), .b(new_n366), .c(new_n133), .out0(\s[8] ));
  nanp02aa1n02x5               g272(.a(new_n117), .b(new_n129), .o1(new_n368));
  aoi113aa1n02x5               g273(.a(new_n143), .b(new_n137), .c(new_n124), .d(new_n130), .e(new_n131), .o1(new_n369));
  aoi022aa1n02x5               g274(.a(new_n145), .b(new_n137), .c(new_n368), .d(new_n369), .o1(\s[9] ));
endmodule


