// Benchmark "adder" written by ABC on Wed Jul 17 14:59:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n319, new_n322, new_n323, new_n324, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor002aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand22aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n09x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  xnrc02aa1n12x5               g007(.a(\b[3] ), .b(\a[4] ), .out0(new_n103));
  nor042aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n03x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb02aa1n06x5               g010(.a(new_n104), .b(new_n105), .out0(new_n106));
  inv000aa1n02x5               g011(.a(new_n104), .o1(new_n107));
  oao003aa1n02x5               g012(.a(\a[4] ), .b(\b[3] ), .c(new_n107), .carry(new_n108));
  oai013aa1d12x5               g013(.a(new_n108), .b(new_n103), .c(new_n102), .d(new_n106), .o1(new_n109));
  xnrc02aa1n12x5               g014(.a(\b[7] ), .b(\a[8] ), .out0(new_n110));
  xnrc02aa1n12x5               g015(.a(\b[6] ), .b(\a[7] ), .out0(new_n111));
  nor002aa1n20x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nor022aa1n16x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand22aa1n09x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nona23aa1n09x5               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  nor043aa1n03x5               g021(.a(new_n116), .b(new_n111), .c(new_n110), .o1(new_n117));
  aoi012aa1n06x5               g022(.a(new_n114), .b(new_n112), .c(new_n115), .o1(new_n118));
  nor002aa1d32x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n119), .o1(new_n120));
  oao003aa1n03x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .carry(new_n121));
  oai013aa1d12x5               g026(.a(new_n121), .b(new_n111), .c(new_n110), .d(new_n118), .o1(new_n122));
  tech160nm_fixorc02aa1n03p5x5 g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  aoai13aa1n02x5               g028(.a(new_n123), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n124));
  tech160nm_fixorc02aa1n03p5x5 g029(.a(\a[10] ), .b(\b[9] ), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n125), .b(new_n124), .c(new_n98), .out0(\s[10] ));
  nand22aa1n03x5               g031(.a(new_n109), .b(new_n117), .o1(new_n127));
  inv000aa1d42x5               g032(.a(new_n122), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(new_n125), .b(new_n123), .o1(new_n129));
  nor002aa1n02x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  oai012aa1n09x5               g036(.a(new_n131), .b(new_n130), .c(new_n97), .o1(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n129), .c(new_n127), .d(new_n128), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1d18x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nanp02aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n135), .out0(new_n138));
  nanp02aa1n03x5               g043(.a(new_n133), .b(new_n138), .o1(new_n139));
  nor042aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n139), .c(new_n136), .out0(\s[12] ));
  nona23aa1d18x5               g048(.a(new_n141), .b(new_n137), .c(new_n135), .d(new_n140), .out0(new_n144));
  nano22aa1n03x7               g049(.a(new_n144), .b(new_n123), .c(new_n125), .out0(new_n145));
  aoai13aa1n06x5               g050(.a(new_n145), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n146));
  oaih12aa1n06x5               g051(.a(new_n141), .b(new_n140), .c(new_n135), .o1(new_n147));
  oai012aa1d24x5               g052(.a(new_n147), .b(new_n144), .c(new_n132), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  norp02aa1n24x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nand42aa1n03x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n146), .c(new_n149), .out0(\s[13] ));
  aobi12aa1n06x5               g058(.a(new_n152), .b(new_n146), .c(new_n149), .out0(new_n154));
  nor042aa1d18x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nand42aa1n04x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  obai22aa1n02x7               g061(.a(new_n156), .b(new_n155), .c(new_n154), .d(new_n150), .out0(new_n157));
  norb03aa1n02x5               g062(.a(new_n156), .b(new_n150), .c(new_n155), .out0(new_n158));
  oaib12aa1n02x5               g063(.a(new_n157), .b(new_n154), .c(new_n158), .out0(\s[14] ));
  tech160nm_fioai012aa1n03p5x5 g064(.a(new_n156), .b(new_n155), .c(new_n150), .o1(new_n160));
  nona23aa1n03x5               g065(.a(new_n156), .b(new_n151), .c(new_n150), .d(new_n155), .out0(new_n161));
  aoai13aa1n06x5               g066(.a(new_n160), .b(new_n161), .c(new_n146), .d(new_n149), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  xorc02aa1n02x5               g069(.a(\a[15] ), .b(\b[14] ), .out0(new_n165));
  tech160nm_fixnrc02aa1n03p5x5 g070(.a(\b[15] ), .b(\a[16] ), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n167));
  norp02aa1n02x5               g072(.a(new_n166), .b(new_n164), .o1(new_n168));
  aob012aa1n02x5               g073(.a(new_n168), .b(new_n162), .c(new_n165), .out0(new_n169));
  nanp02aa1n02x5               g074(.a(new_n167), .b(new_n169), .o1(\s[16] ));
  nano23aa1n06x5               g075(.a(new_n135), .b(new_n140), .c(new_n141), .d(new_n137), .out0(new_n171));
  nano23aa1n02x5               g076(.a(new_n150), .b(new_n155), .c(new_n156), .d(new_n151), .out0(new_n172));
  xorc02aa1n02x5               g077(.a(\a[16] ), .b(\b[15] ), .out0(new_n173));
  nanp03aa1n02x5               g078(.a(new_n172), .b(new_n165), .c(new_n173), .o1(new_n174));
  nano32aa1n03x7               g079(.a(new_n174), .b(new_n171), .c(new_n125), .d(new_n123), .out0(new_n175));
  aoai13aa1n12x5               g080(.a(new_n175), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n176));
  tech160nm_fixnrc02aa1n02p5x5 g081(.a(\b[14] ), .b(\a[15] ), .out0(new_n177));
  nor043aa1n03x5               g082(.a(new_n161), .b(new_n166), .c(new_n177), .o1(new_n178));
  orn002aa1n02x5               g083(.a(\a[15] ), .b(\b[14] ), .o(new_n179));
  oao003aa1n02x5               g084(.a(\a[16] ), .b(\b[15] ), .c(new_n179), .carry(new_n180));
  oai013aa1n03x5               g085(.a(new_n180), .b(new_n166), .c(new_n177), .d(new_n160), .o1(new_n181));
  aoi012aa1d18x5               g086(.a(new_n181), .b(new_n148), .c(new_n178), .o1(new_n182));
  xorc02aa1n02x5               g087(.a(\a[17] ), .b(\b[16] ), .out0(new_n183));
  xnbna2aa1n03x5               g088(.a(new_n183), .b(new_n176), .c(new_n182), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[17] ), .o1(new_n185));
  inv040aa1d32x5               g090(.a(\b[16] ), .o1(new_n186));
  nand42aa1d28x5               g091(.a(new_n186), .b(new_n185), .o1(new_n187));
  nand02aa1n02x5               g092(.a(new_n145), .b(new_n178), .o1(new_n188));
  aoai13aa1n09x5               g093(.a(new_n182), .b(new_n188), .c(new_n127), .d(new_n128), .o1(new_n189));
  nanp02aa1n03x5               g094(.a(new_n189), .b(new_n183), .o1(new_n190));
  norp02aa1n02x5               g095(.a(\b[17] ), .b(\a[18] ), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  xobna2aa1n03x5               g098(.a(new_n193), .b(new_n190), .c(new_n187), .out0(\s[18] ));
  inv000aa1d42x5               g099(.a(\a[18] ), .o1(new_n195));
  xroi22aa1d06x4               g100(.a(new_n185), .b(\b[16] ), .c(new_n195), .d(\b[17] ), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  oaoi03aa1n12x5               g102(.a(\a[18] ), .b(\b[17] ), .c(new_n187), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n197), .c(new_n176), .d(new_n182), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g106(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n09x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand42aa1n20x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nor042aa1n09x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand42aa1n20x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  aoai13aa1n02x5               g112(.a(new_n207), .b(new_n203), .c(new_n200), .d(new_n204), .o1(new_n208));
  nanp02aa1n03x5               g113(.a(new_n189), .b(new_n196), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n203), .b(new_n204), .out0(new_n210));
  norb03aa1n02x5               g115(.a(new_n206), .b(new_n203), .c(new_n205), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n210), .c(new_n209), .d(new_n199), .o1(new_n212));
  nanp02aa1n03x5               g117(.a(new_n208), .b(new_n212), .o1(\s[20] ));
  nano23aa1d15x5               g118(.a(new_n203), .b(new_n205), .c(new_n206), .d(new_n204), .out0(new_n214));
  nanb03aa1n06x5               g119(.a(new_n193), .b(new_n214), .c(new_n183), .out0(new_n215));
  nand22aa1n09x5               g120(.a(new_n214), .b(new_n198), .o1(new_n216));
  oaih12aa1n12x5               g121(.a(new_n206), .b(new_n205), .c(new_n203), .o1(new_n217));
  nand02aa1d04x5               g122(.a(new_n216), .b(new_n217), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n06x5               g124(.a(new_n219), .b(new_n215), .c(new_n176), .d(new_n182), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  nand02aa1d24x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  nor042aa1n06x5               g129(.a(\b[21] ), .b(\a[22] ), .o1(new_n225));
  nand02aa1d20x5               g130(.a(\b[21] ), .b(\a[22] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n228), .b(new_n222), .c(new_n220), .d(new_n224), .o1(new_n229));
  nand22aa1n03x5               g134(.a(new_n220), .b(new_n224), .o1(new_n230));
  norb03aa1n02x5               g135(.a(new_n226), .b(new_n222), .c(new_n225), .out0(new_n231));
  nand22aa1n03x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  nanp02aa1n03x5               g137(.a(new_n229), .b(new_n232), .o1(\s[22] ));
  nano23aa1d15x5               g138(.a(new_n222), .b(new_n225), .c(new_n226), .d(new_n223), .out0(new_n234));
  nanp03aa1n02x5               g139(.a(new_n196), .b(new_n214), .c(new_n234), .o1(new_n235));
  ao0012aa1n03x7               g140(.a(new_n225), .b(new_n222), .c(new_n226), .o(new_n236));
  tech160nm_fiaoi012aa1n04x5   g141(.a(new_n236), .b(new_n218), .c(new_n234), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n237), .b(new_n235), .c(new_n176), .d(new_n182), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  inv000aa1d42x5               g144(.a(new_n214), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n234), .o1(new_n241));
  nona32aa1n03x5               g146(.a(new_n189), .b(new_n241), .c(new_n240), .d(new_n197), .out0(new_n242));
  norp02aa1n24x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  nand02aa1d24x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  aoi012aa1n03x5               g151(.a(new_n246), .b(new_n242), .c(new_n237), .o1(new_n247));
  nor002aa1n10x5               g152(.a(\b[23] ), .b(\a[24] ), .o1(new_n248));
  nand02aa1d16x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  nanb02aa1n02x5               g154(.a(new_n248), .b(new_n249), .out0(new_n250));
  aoai13aa1n03x5               g155(.a(new_n250), .b(new_n243), .c(new_n238), .d(new_n245), .o1(new_n251));
  nona22aa1n03x5               g156(.a(new_n249), .b(new_n248), .c(new_n243), .out0(new_n252));
  tech160nm_fioai012aa1n02p5x5 g157(.a(new_n251), .b(new_n247), .c(new_n252), .o1(\s[24] ));
  nano23aa1n03x7               g158(.a(new_n243), .b(new_n248), .c(new_n249), .d(new_n244), .out0(new_n254));
  nona23aa1n02x4               g159(.a(new_n196), .b(new_n254), .c(new_n241), .d(new_n240), .out0(new_n255));
  nand22aa1n03x5               g160(.a(new_n254), .b(new_n234), .o1(new_n256));
  aoi022aa1n06x5               g161(.a(new_n254), .b(new_n236), .c(new_n249), .d(new_n252), .o1(new_n257));
  aoai13aa1n12x5               g162(.a(new_n257), .b(new_n256), .c(new_n216), .d(new_n217), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n255), .c(new_n176), .d(new_n182), .o1(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[24] ), .b(\a[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  xnrc02aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n262), .c(new_n260), .d(new_n264), .o1(new_n266));
  nona32aa1n03x5               g171(.a(new_n189), .b(new_n256), .c(new_n240), .d(new_n197), .out0(new_n267));
  norp02aa1n02x5               g172(.a(new_n265), .b(new_n262), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n263), .c(new_n267), .d(new_n259), .o1(new_n269));
  nanp02aa1n03x5               g174(.a(new_n266), .b(new_n269), .o1(\s[26] ));
  nor042aa1n02x5               g175(.a(new_n265), .b(new_n263), .o1(new_n271));
  nano32aa1n03x7               g176(.a(new_n215), .b(new_n271), .c(new_n234), .d(new_n254), .out0(new_n272));
  inv020aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\a[26] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(\b[25] ), .o1(new_n275));
  oaoi03aa1n02x5               g180(.a(new_n274), .b(new_n275), .c(new_n262), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  aoi012aa1n06x5               g182(.a(new_n277), .b(new_n258), .c(new_n271), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n273), .c(new_n176), .d(new_n182), .o1(new_n279));
  xorb03aa1n03x5               g184(.a(new_n279), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g185(.a(\b[26] ), .b(\a[27] ), .o1(new_n281));
  xorc02aa1n02x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n281), .c(new_n279), .d(new_n282), .o1(new_n284));
  nand22aa1n03x5               g189(.a(new_n258), .b(new_n271), .o1(new_n285));
  nand02aa1d04x5               g190(.a(new_n285), .b(new_n276), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n282), .b(new_n286), .c(new_n189), .d(new_n272), .o1(new_n287));
  nona22aa1n03x5               g192(.a(new_n287), .b(new_n283), .c(new_n281), .out0(new_n288));
  nanp02aa1n03x5               g193(.a(new_n284), .b(new_n288), .o1(\s[28] ));
  tech160nm_fixorc02aa1n03p5x5 g194(.a(\a[29] ), .b(\b[28] ), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  norb02aa1n02x5               g196(.a(new_n282), .b(new_n283), .out0(new_n292));
  inv000aa1d42x5               g197(.a(\a[28] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  oaoi03aa1n06x5               g199(.a(new_n293), .b(new_n294), .c(new_n281), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n291), .b(new_n296), .c(new_n279), .d(new_n292), .o1(new_n297));
  aoai13aa1n02x7               g202(.a(new_n292), .b(new_n286), .c(new_n189), .d(new_n272), .o1(new_n298));
  nona22aa1n03x5               g203(.a(new_n298), .b(new_n296), .c(new_n291), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g206(.a(new_n283), .b(new_n282), .c(new_n290), .out0(new_n302));
  oaoi03aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .o1(new_n303));
  tech160nm_fixorc02aa1n03p5x5 g208(.a(\a[30] ), .b(\b[29] ), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  aoai13aa1n02x7               g210(.a(new_n305), .b(new_n303), .c(new_n279), .d(new_n302), .o1(new_n306));
  aoai13aa1n02x7               g211(.a(new_n302), .b(new_n286), .c(new_n189), .d(new_n272), .o1(new_n307));
  nona22aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n305), .out0(new_n308));
  nanp02aa1n03x5               g213(.a(new_n306), .b(new_n308), .o1(\s[30] ));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  nano23aa1n02x4               g215(.a(new_n305), .b(new_n283), .c(new_n282), .d(new_n290), .out0(new_n311));
  and002aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .o(new_n312));
  oab012aa1n02x4               g217(.a(new_n312), .b(new_n303), .c(new_n305), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n310), .b(new_n313), .c(new_n279), .d(new_n311), .o1(new_n314));
  aoai13aa1n02x7               g219(.a(new_n311), .b(new_n286), .c(new_n189), .d(new_n272), .o1(new_n315));
  nona22aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n310), .out0(new_n316));
  nanp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[31] ));
  xnbna2aa1n03x5               g222(.a(new_n102), .b(new_n105), .c(new_n107), .out0(\s[3] ));
  orn002aa1n02x5               g223(.a(new_n102), .b(new_n106), .o(new_n319));
  xobna2aa1n03x5               g224(.a(new_n103), .b(new_n319), .c(new_n107), .out0(\s[4] ));
  xorb03aa1n02x5               g225(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g226(.a(new_n114), .b(new_n115), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n322), .b(new_n112), .c(new_n109), .d(new_n113), .o1(new_n323));
  aoi112aa1n02x5               g228(.a(new_n112), .b(new_n322), .c(new_n109), .d(new_n113), .o1(new_n324));
  nanb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(\s[6] ));
  oaib12aa1n02x5               g230(.a(new_n118), .b(new_n116), .c(new_n109), .out0(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g232(.a(new_n111), .b(new_n326), .out0(new_n328));
  xobna2aa1n03x5               g233(.a(new_n110), .b(new_n328), .c(new_n120), .out0(\s[8] ));
  xnbna2aa1n03x5               g234(.a(new_n123), .b(new_n127), .c(new_n128), .out0(\s[9] ));
endmodule


