// Benchmark "adder" written by ABC on Wed Jul 17 18:09:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n326, new_n327, new_n330, new_n331, new_n332, new_n334,
    new_n336, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n12x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nor002aa1n02x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand22aa1n03x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nanp02aa1n03x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai112aa1n06x5               g007(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n103));
  aoi113aa1n06x5               g008(.a(new_n100), .b(new_n99), .c(new_n103), .d(new_n102), .e(new_n101), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nanp02aa1n06x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nanp02aa1n09x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nano23aa1n09x5               g013(.a(new_n105), .b(new_n107), .c(new_n108), .d(new_n106), .out0(new_n109));
  inv000aa1d42x5               g014(.a(\a[6] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[5] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nand22aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand02aa1d06x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nor042aa1d18x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand02aa1n04x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanb02aa1n06x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  nano32aa1n03x7               g022(.a(new_n117), .b(new_n112), .c(new_n113), .d(new_n114), .out0(new_n118));
  nand22aa1n03x5               g023(.a(new_n118), .b(new_n109), .o1(new_n119));
  aob012aa1n03x5               g024(.a(new_n112), .b(new_n115), .c(new_n113), .out0(new_n120));
  inv000aa1d42x5               g025(.a(new_n107), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[8] ), .b(\b[7] ), .c(new_n121), .o1(new_n122));
  aoi012aa1n06x5               g027(.a(new_n122), .b(new_n109), .c(new_n120), .o1(new_n123));
  oai012aa1n18x5               g028(.a(new_n123), .b(new_n119), .c(new_n104), .o1(new_n124));
  xnrc02aa1n12x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(new_n124), .b(new_n126), .o1(new_n127));
  nor042aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand02aa1n04x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n03x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  aoai13aa1n06x5               g036(.a(new_n130), .b(new_n97), .c(new_n124), .d(new_n126), .o1(new_n132));
  tech160nm_fiaoi012aa1n05x5   g037(.a(new_n128), .b(new_n97), .c(new_n129), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanp02aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  inv000aa1d42x5               g041(.a(new_n136), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n132), .c(new_n133), .out0(\s[11] ));
  aob012aa1n03x5               g043(.a(new_n137), .b(new_n132), .c(new_n133), .out0(new_n139));
  nor042aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand02aa1n06x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  aoib12aa1n02x5               g048(.a(new_n134), .b(new_n141), .c(new_n140), .out0(new_n144));
  oai012aa1n02x5               g049(.a(new_n139), .b(\b[10] ), .c(\a[11] ), .o1(new_n145));
  aoi022aa1n02x5               g050(.a(new_n145), .b(new_n143), .c(new_n139), .d(new_n144), .o1(\s[12] ));
  inv040aa1n03x5               g051(.a(new_n130), .o1(new_n147));
  nona23aa1n02x4               g052(.a(new_n141), .b(new_n135), .c(new_n134), .d(new_n140), .out0(new_n148));
  nor003aa1n03x5               g053(.a(new_n148), .b(new_n147), .c(new_n125), .o1(new_n149));
  aoi012aa1n02x7               g054(.a(new_n140), .b(new_n134), .c(new_n141), .o1(new_n150));
  oai012aa1n02x5               g055(.a(new_n150), .b(new_n148), .c(new_n133), .o1(new_n151));
  inv040aa1n02x5               g056(.a(new_n151), .o1(new_n152));
  aob012aa1n06x5               g057(.a(new_n152), .b(new_n124), .c(new_n149), .out0(new_n153));
  nor002aa1d32x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand22aa1n06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n154), .b(new_n155), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoi112aa1n02x5               g062(.a(new_n157), .b(new_n151), .c(new_n124), .d(new_n149), .o1(new_n158));
  aoi012aa1n02x5               g063(.a(new_n158), .b(new_n153), .c(new_n157), .o1(\s[13] ));
  inv040aa1n08x5               g064(.a(new_n154), .o1(new_n160));
  aoai13aa1n02x5               g065(.a(new_n157), .b(new_n151), .c(new_n124), .d(new_n149), .o1(new_n161));
  nor042aa1n02x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand02aa1d04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  xobna2aa1n03x5               g069(.a(new_n164), .b(new_n161), .c(new_n160), .out0(\s[14] ));
  nano23aa1n06x5               g070(.a(new_n154), .b(new_n162), .c(new_n163), .d(new_n155), .out0(new_n166));
  oaoi03aa1n12x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .o1(new_n167));
  nor042aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n10x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n167), .c(new_n153), .d(new_n166), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n170), .b(new_n167), .c(new_n153), .d(new_n166), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[15] ));
  nor042aa1n09x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1d28x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  aoib12aa1n02x5               g081(.a(new_n168), .b(new_n175), .c(new_n174), .out0(new_n177));
  tech160nm_fioai012aa1n03p5x5 g082(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .o1(new_n178));
  aoi022aa1n02x7               g083(.a(new_n178), .b(new_n176), .c(new_n171), .d(new_n177), .o1(\s[16] ));
  nano23aa1n06x5               g084(.a(new_n134), .b(new_n140), .c(new_n141), .d(new_n135), .out0(new_n180));
  nano23aa1n09x5               g085(.a(new_n168), .b(new_n174), .c(new_n175), .d(new_n169), .out0(new_n181));
  nand02aa1d04x5               g086(.a(new_n181), .b(new_n166), .o1(new_n182));
  nano32aa1n03x7               g087(.a(new_n182), .b(new_n126), .c(new_n180), .d(new_n130), .out0(new_n183));
  nand02aa1n04x5               g088(.a(new_n124), .b(new_n183), .o1(new_n184));
  nanb02aa1n03x5               g089(.a(new_n133), .b(new_n180), .out0(new_n185));
  ao0012aa1n03x7               g090(.a(new_n174), .b(new_n168), .c(new_n175), .o(new_n186));
  aoi012aa1d24x5               g091(.a(new_n186), .b(new_n181), .c(new_n167), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n182), .c(new_n185), .d(new_n150), .o1(new_n188));
  nanb02aa1n12x5               g093(.a(new_n188), .b(new_n184), .out0(new_n189));
  tech160nm_fixorc02aa1n05x5   g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  nona23aa1n02x4               g095(.a(new_n163), .b(new_n155), .c(new_n154), .d(new_n162), .out0(new_n191));
  nano22aa1n02x4               g096(.a(new_n191), .b(new_n170), .c(new_n176), .out0(new_n192));
  inv000aa1d42x5               g097(.a(new_n187), .o1(new_n193));
  aoi112aa1n02x5               g098(.a(new_n193), .b(new_n190), .c(new_n151), .d(new_n192), .o1(new_n194));
  aoi022aa1n02x5               g099(.a(new_n189), .b(new_n190), .c(new_n184), .d(new_n194), .o1(\s[17] ));
  norp02aa1n02x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  aoai13aa1n02x5               g102(.a(new_n190), .b(new_n188), .c(new_n124), .d(new_n183), .o1(new_n198));
  xorc02aa1n12x5               g103(.a(\a[18] ), .b(\b[17] ), .out0(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n198), .c(new_n197), .out0(\s[18] ));
  and002aa1n02x5               g105(.a(new_n199), .b(new_n190), .o(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n188), .c(new_n124), .d(new_n183), .o1(new_n202));
  nor042aa1n02x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  aoi112aa1n09x5               g108(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n204));
  norp02aa1n02x5               g109(.a(new_n204), .b(new_n203), .o1(new_n205));
  nor002aa1d32x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand02aa1n08x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  norb02aa1n12x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n202), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g115(.a(new_n208), .b(new_n202), .c(new_n205), .out0(new_n211));
  nor042aa1n06x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand02aa1n08x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n06x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  aoib12aa1n02x5               g119(.a(new_n206), .b(new_n213), .c(new_n212), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n206), .o1(new_n216));
  nanp02aa1n03x5               g121(.a(new_n211), .b(new_n216), .o1(new_n217));
  aoi022aa1n02x5               g122(.a(new_n217), .b(new_n214), .c(new_n211), .d(new_n215), .o1(\s[20] ));
  nano23aa1n09x5               g123(.a(new_n206), .b(new_n212), .c(new_n213), .d(new_n207), .out0(new_n219));
  nand23aa1n06x5               g124(.a(new_n219), .b(new_n190), .c(new_n199), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n188), .c(new_n124), .d(new_n183), .o1(new_n222));
  oai112aa1n06x5               g127(.a(new_n208), .b(new_n214), .c(new_n204), .d(new_n203), .o1(new_n223));
  oaih12aa1n02x5               g128(.a(new_n213), .b(new_n212), .c(new_n206), .o1(new_n224));
  nanp02aa1n02x5               g129(.a(new_n223), .b(new_n224), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  xorc02aa1n12x5               g131(.a(\a[21] ), .b(\b[20] ), .out0(new_n227));
  xnbna2aa1n03x5               g132(.a(new_n227), .b(new_n222), .c(new_n226), .out0(\s[21] ));
  aob012aa1n03x5               g133(.a(new_n227), .b(new_n222), .c(new_n226), .out0(new_n229));
  xorc02aa1n02x5               g134(.a(\a[22] ), .b(\b[21] ), .out0(new_n230));
  norp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norp02aa1n02x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\a[21] ), .o1(new_n233));
  oaib12aa1n06x5               g138(.a(new_n229), .b(\b[20] ), .c(new_n233), .out0(new_n234));
  aoi022aa1n02x7               g139(.a(new_n234), .b(new_n230), .c(new_n229), .d(new_n232), .o1(\s[22] ));
  nand02aa1d04x5               g140(.a(new_n230), .b(new_n227), .o1(new_n236));
  nano32aa1n02x4               g141(.a(new_n236), .b(new_n219), .c(new_n199), .d(new_n190), .out0(new_n237));
  inv000aa1d42x5               g142(.a(\a[22] ), .o1(new_n238));
  oai022aa1n02x5               g143(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n239));
  oaib12aa1n02x5               g144(.a(new_n239), .b(new_n238), .c(\b[21] ), .out0(new_n240));
  aoai13aa1n12x5               g145(.a(new_n240), .b(new_n236), .c(new_n223), .d(new_n224), .o1(new_n241));
  xorc02aa1n02x5               g146(.a(\a[23] ), .b(\b[22] ), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n241), .c(new_n189), .d(new_n237), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(new_n242), .b(new_n241), .c(new_n189), .d(new_n237), .o1(new_n244));
  norb02aa1n03x4               g149(.a(new_n243), .b(new_n244), .out0(\s[23] ));
  xorc02aa1n02x5               g150(.a(\a[24] ), .b(\b[23] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(\a[23] ), .o1(new_n247));
  nanb02aa1n02x5               g152(.a(\b[22] ), .b(new_n247), .out0(new_n248));
  norb02aa1n02x5               g153(.a(new_n248), .b(new_n246), .out0(new_n249));
  nanp02aa1n03x5               g154(.a(new_n243), .b(new_n248), .o1(new_n250));
  aoi022aa1n02x7               g155(.a(new_n250), .b(new_n246), .c(new_n243), .d(new_n249), .o1(\s[24] ));
  xroi22aa1d04x5               g156(.a(new_n233), .b(\b[20] ), .c(new_n238), .d(\b[21] ), .out0(new_n252));
  inv000aa1d42x5               g157(.a(\a[24] ), .o1(new_n253));
  xroi22aa1d04x5               g158(.a(new_n247), .b(\b[22] ), .c(new_n253), .d(\b[23] ), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n220), .b(new_n252), .c(new_n254), .out0(new_n255));
  oaoi03aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n248), .o1(new_n256));
  tech160nm_fiao0012aa1n02p5x5 g161(.a(new_n256), .b(new_n241), .c(new_n254), .o(new_n257));
  tech160nm_fixorc02aa1n03p5x5 g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n257), .c(new_n189), .d(new_n255), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(new_n258), .b(new_n257), .c(new_n189), .d(new_n255), .o1(new_n260));
  norb02aa1n02x5               g165(.a(new_n259), .b(new_n260), .out0(\s[25] ));
  xorc02aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .out0(new_n262));
  orn002aa1n24x5               g167(.a(\a[25] ), .b(\b[24] ), .o(new_n263));
  norb02aa1n02x5               g168(.a(new_n263), .b(new_n262), .out0(new_n264));
  nanp02aa1n03x5               g169(.a(new_n259), .b(new_n263), .o1(new_n265));
  aoi022aa1n02x7               g170(.a(new_n265), .b(new_n262), .c(new_n259), .d(new_n264), .o1(\s[26] ));
  and002aa1n02x5               g171(.a(new_n262), .b(new_n258), .o(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n256), .c(new_n241), .d(new_n254), .o1(new_n268));
  nano32aa1n03x7               g173(.a(new_n220), .b(new_n267), .c(new_n252), .d(new_n254), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n188), .c(new_n124), .d(new_n183), .o1(new_n270));
  oaoi03aa1n02x5               g175(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .o1(new_n271));
  inv000aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  nand23aa1n06x5               g177(.a(new_n270), .b(new_n268), .c(new_n272), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  nona22aa1n02x4               g179(.a(new_n270), .b(new_n271), .c(new_n274), .out0(new_n275));
  aboi22aa1n03x5               g180(.a(new_n275), .b(new_n268), .c(new_n273), .d(new_n274), .out0(\s[27] ));
  nanp02aa1n06x5               g181(.a(new_n273), .b(new_n274), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[28] ), .b(\b[27] ), .out0(new_n278));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  norp02aa1n02x5               g184(.a(new_n278), .b(new_n279), .o1(new_n280));
  nor002aa1n02x5               g185(.a(new_n100), .b(new_n99), .o1(new_n281));
  inv000aa1d42x5               g186(.a(\a[3] ), .o1(new_n282));
  inv000aa1d42x5               g187(.a(\b[2] ), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n283), .b(new_n282), .o1(new_n284));
  nanp02aa1n02x5               g189(.a(new_n284), .b(new_n101), .o1(new_n285));
  norp02aa1n02x5               g190(.a(\b[1] ), .b(\a[2] ), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(\b[0] ), .b(\a[1] ), .o1(new_n287));
  oai012aa1n02x5               g192(.a(new_n102), .b(new_n286), .c(new_n287), .o1(new_n288));
  tech160nm_fioai012aa1n05x5   g193(.a(new_n281), .b(new_n288), .c(new_n285), .o1(new_n289));
  nanp03aa1n03x5               g194(.a(new_n289), .b(new_n109), .c(new_n118), .o1(new_n290));
  nanp02aa1n03x5               g195(.a(new_n149), .b(new_n192), .o1(new_n291));
  tech160nm_fiaoi012aa1n03p5x5 g196(.a(new_n291), .b(new_n290), .c(new_n123), .o1(new_n292));
  oaoi13aa1n06x5               g197(.a(new_n271), .b(new_n269), .c(new_n292), .d(new_n188), .o1(new_n293));
  inv000aa1n03x5               g198(.a(new_n279), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n274), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n294), .b(new_n295), .c(new_n293), .d(new_n268), .o1(new_n296));
  aoi022aa1n03x5               g201(.a(new_n296), .b(new_n278), .c(new_n277), .d(new_n280), .o1(\s[28] ));
  and002aa1n06x5               g202(.a(new_n278), .b(new_n274), .o(new_n298));
  tech160nm_finand02aa1n05x5   g203(.a(new_n273), .b(new_n298), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .out0(new_n300));
  oao003aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n294), .carry(new_n301));
  norb02aa1n02x5               g206(.a(new_n301), .b(new_n300), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n298), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n301), .b(new_n303), .c(new_n293), .d(new_n268), .o1(new_n304));
  aoi022aa1n03x5               g209(.a(new_n304), .b(new_n300), .c(new_n299), .d(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n287), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g211(.a(new_n295), .b(new_n278), .c(new_n300), .out0(new_n307));
  inv000aa1n02x5               g212(.a(new_n307), .o1(new_n308));
  aoi013aa1n03x5               g213(.a(new_n308), .b(new_n270), .c(new_n268), .d(new_n272), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .out0(new_n310));
  oab012aa1n02x4               g215(.a(new_n310), .b(\a[29] ), .c(\b[28] ), .out0(new_n311));
  aoai13aa1n02x5               g216(.a(new_n311), .b(new_n301), .c(\a[29] ), .d(\b[28] ), .o1(new_n312));
  tech160nm_fiaoi012aa1n05x5   g217(.a(new_n312), .b(new_n273), .c(new_n307), .o1(new_n313));
  oaoi03aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .o1(new_n314));
  oaoi13aa1n02x7               g219(.a(new_n313), .b(new_n310), .c(new_n314), .d(new_n309), .o1(\s[30] ));
  nanp03aa1n02x5               g220(.a(new_n298), .b(new_n300), .c(new_n310), .o1(new_n316));
  nanb02aa1n03x5               g221(.a(new_n316), .b(new_n273), .out0(new_n317));
  xorc02aa1n02x5               g222(.a(\a[31] ), .b(\b[30] ), .out0(new_n318));
  oabi12aa1n02x5               g223(.a(new_n314), .b(\a[30] ), .c(\b[29] ), .out0(new_n319));
  aob012aa1n02x5               g224(.a(new_n319), .b(\b[29] ), .c(\a[30] ), .out0(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n318), .out0(new_n321));
  aoai13aa1n02x5               g226(.a(new_n320), .b(new_n316), .c(new_n293), .d(new_n268), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n322), .b(new_n318), .c(new_n317), .d(new_n321), .o1(\s[31] ));
  xnbna2aa1n03x5               g228(.a(new_n285), .b(new_n103), .c(new_n102), .out0(\s[3] ));
  inv000aa1d42x5               g229(.a(new_n99), .o1(new_n325));
  norb02aa1n02x5               g230(.a(new_n114), .b(new_n99), .out0(new_n326));
  aoi113aa1n02x5               g231(.a(new_n100), .b(new_n326), .c(new_n103), .d(new_n102), .e(new_n101), .o1(new_n327));
  aoi013aa1n02x4               g232(.a(new_n327), .b(new_n289), .c(new_n114), .d(new_n325), .o1(\s[4] ));
  xnbna2aa1n03x5               g233(.a(new_n117), .b(new_n289), .c(new_n114), .out0(\s[5] ));
  xorc02aa1n02x5               g234(.a(\a[6] ), .b(\b[5] ), .out0(new_n330));
  aoi013aa1n02x4               g235(.a(new_n115), .b(new_n289), .c(new_n114), .d(new_n116), .o1(new_n331));
  aoi113aa1n02x5               g236(.a(new_n115), .b(new_n330), .c(new_n289), .d(new_n116), .e(new_n114), .o1(new_n332));
  aoib12aa1n02x5               g237(.a(new_n332), .b(new_n330), .c(new_n331), .out0(\s[6] ));
  aoi012aa1n02x5               g238(.a(new_n120), .b(new_n289), .c(new_n118), .o1(new_n334));
  xnbna2aa1n03x5               g239(.a(new_n334), .b(new_n121), .c(new_n108), .out0(\s[7] ));
  norb02aa1n02x5               g240(.a(new_n106), .b(new_n105), .out0(new_n336));
  nanb03aa1n02x5               g241(.a(new_n334), .b(new_n121), .c(new_n108), .out0(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n336), .b(new_n337), .c(new_n121), .out0(\s[8] ));
  xnbna2aa1n03x5               g243(.a(new_n126), .b(new_n290), .c(new_n123), .out0(\s[9] ));
endmodule


