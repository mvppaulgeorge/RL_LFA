// Benchmark "adder" written by ABC on Wed Jul 17 20:06:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n140, new_n141, new_n142, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n327, new_n328, new_n329, new_n331, new_n333,
    new_n334, new_n335, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nor022aa1n04x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nand42aa1n03x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nanb02aa1n12x5               g005(.a(new_n99), .b(new_n100), .out0(new_n101));
  orn002aa1n02x7               g006(.a(\a[2] ), .b(\b[1] ), .o(new_n102));
  nand42aa1n03x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  aob012aa1n03x5               g008(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(new_n104));
  nand42aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor002aa1n02x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb03aa1n03x4               g011(.a(new_n105), .b(new_n99), .c(new_n106), .out0(new_n107));
  aoai13aa1n06x5               g012(.a(new_n107), .b(new_n101), .c(new_n104), .d(new_n102), .o1(new_n108));
  nand02aa1d20x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[6] ), .o1(new_n110));
  nanb02aa1n02x5               g015(.a(\a[7] ), .b(new_n110), .out0(new_n111));
  nand42aa1n03x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor042aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanb02aa1n06x5               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  nano32aa1n09x5               g020(.a(new_n115), .b(new_n111), .c(new_n112), .d(new_n109), .out0(new_n116));
  nor042aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor022aa1n08x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nand42aa1n03x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n118), .b(new_n117), .c(new_n119), .d(new_n105), .out0(new_n120));
  nand23aa1n06x5               g025(.a(new_n108), .b(new_n116), .c(new_n120), .o1(new_n121));
  nor042aa1n02x5               g026(.a(new_n118), .b(new_n117), .o1(new_n122));
  inv040aa1n03x5               g027(.a(new_n122), .o1(new_n123));
  nor002aa1n02x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  tech160nm_fiaoi012aa1n05x5   g029(.a(new_n114), .b(new_n124), .c(new_n113), .o1(new_n125));
  inv030aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  aoi012aa1n12x5               g031(.a(new_n126), .b(new_n116), .c(new_n123), .o1(new_n127));
  nand02aa1n08x5               g032(.a(new_n121), .b(new_n127), .o1(new_n128));
  oaoi03aa1n02x5               g033(.a(new_n97), .b(new_n98), .c(new_n128), .o1(new_n129));
  nor002aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  inv020aa1n02x5               g035(.a(new_n130), .o1(new_n131));
  nand02aa1n10x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(new_n98), .b(new_n97), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[8] ), .b(\a[9] ), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(new_n133), .b(new_n134), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n132), .o1(new_n136));
  aoi112aa1n09x5               g041(.a(new_n136), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n137));
  aoai13aa1n06x5               g042(.a(new_n137), .b(new_n135), .c(new_n121), .d(new_n127), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n129), .c(new_n132), .d(new_n131), .o1(\s[10] ));
  nand02aa1d06x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nor042aa1n06x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n132), .out0(\s[11] ));
  aoi013aa1n02x4               g048(.a(new_n141), .b(new_n138), .c(new_n140), .d(new_n132), .o1(new_n144));
  xnrb03aa1n02x5               g049(.a(new_n144), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n04x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand22aa1n12x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nano23aa1n06x5               g052(.a(new_n146), .b(new_n141), .c(new_n147), .d(new_n140), .out0(new_n148));
  oai112aa1n03x5               g053(.a(new_n133), .b(new_n134), .c(\b[9] ), .d(\a[10] ), .o1(new_n149));
  nona22aa1n02x4               g054(.a(new_n148), .b(new_n149), .c(new_n136), .out0(new_n150));
  nona23aa1d18x5               g055(.a(new_n140), .b(new_n147), .c(new_n146), .d(new_n141), .out0(new_n151));
  aoi012aa1d24x5               g056(.a(new_n146), .b(new_n141), .c(new_n147), .o1(new_n152));
  oai013aa1d12x5               g057(.a(new_n152), .b(new_n151), .c(new_n137), .d(new_n136), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n150), .c(new_n121), .d(new_n127), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d24x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nanp02aa1n06x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  aoi012aa1n03x5               g063(.a(new_n157), .b(new_n155), .c(new_n158), .o1(new_n159));
  xnrb03aa1n03x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n10x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanp02aa1n06x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nano23aa1n06x5               g067(.a(new_n157), .b(new_n161), .c(new_n162), .d(new_n158), .out0(new_n163));
  tech160nm_fioai012aa1n04x5   g068(.a(new_n162), .b(new_n161), .c(new_n157), .o1(new_n164));
  inv030aa1n03x5               g069(.a(new_n164), .o1(new_n165));
  xorc02aa1n12x5               g070(.a(\a[15] ), .b(\b[14] ), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n165), .c(new_n155), .d(new_n163), .o1(new_n167));
  aoi112aa1n02x5               g072(.a(new_n166), .b(new_n165), .c(new_n155), .d(new_n163), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n167), .b(new_n168), .out0(\s[15] ));
  norp02aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  tech160nm_fixorc02aa1n05x5   g075(.a(\a[16] ), .b(\b[15] ), .out0(new_n171));
  nona22aa1n03x5               g076(.a(new_n167), .b(new_n171), .c(new_n170), .out0(new_n172));
  xnrc02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .out0(new_n173));
  oaoi13aa1n04x5               g078(.a(new_n173), .b(new_n167), .c(\a[15] ), .d(\b[14] ), .o1(new_n174));
  norb02aa1n03x4               g079(.a(new_n172), .b(new_n174), .out0(\s[16] ));
  norb02aa1n02x7               g080(.a(new_n112), .b(new_n124), .out0(new_n176));
  norb02aa1n02x5               g081(.a(new_n113), .b(new_n114), .out0(new_n177));
  nona23aa1n02x4               g082(.a(new_n105), .b(new_n119), .c(new_n118), .d(new_n117), .out0(new_n178));
  nano32aa1n03x5               g083(.a(new_n178), .b(new_n177), .c(new_n176), .d(new_n109), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n109), .o1(new_n180));
  nona23aa1n03x5               g085(.a(new_n177), .b(new_n176), .c(new_n122), .d(new_n180), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n181), .b(new_n125), .o1(new_n182));
  aoi012aa1n03x5               g087(.a(new_n182), .b(new_n179), .c(new_n108), .o1(new_n183));
  nona23aa1n03x5               g088(.a(new_n162), .b(new_n158), .c(new_n157), .d(new_n161), .out0(new_n184));
  xnrc02aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .out0(new_n185));
  norp03aa1n02x5               g090(.a(new_n184), .b(new_n185), .c(new_n173), .o1(new_n186));
  nona32aa1n03x5               g091(.a(new_n186), .b(new_n151), .c(new_n149), .d(new_n136), .out0(new_n187));
  inv000aa1d42x5               g092(.a(\a[16] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[15] ), .o1(new_n189));
  oaoi03aa1n02x5               g094(.a(new_n188), .b(new_n189), .c(new_n170), .o1(new_n190));
  oai013aa1n02x4               g095(.a(new_n190), .b(new_n185), .c(new_n173), .d(new_n164), .o1(new_n191));
  tech160nm_fiaoi012aa1n05x5   g096(.a(new_n191), .b(new_n153), .c(new_n186), .o1(new_n192));
  oai012aa1n06x5               g097(.a(new_n192), .b(new_n183), .c(new_n187), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g099(.a(\a[18] ), .o1(new_n195));
  aoi012aa1n06x5               g100(.a(new_n187), .b(new_n121), .c(new_n127), .o1(new_n196));
  oai112aa1n02x5               g101(.a(new_n131), .b(new_n132), .c(\b[8] ), .d(\a[9] ), .o1(new_n197));
  nanp03aa1n06x5               g102(.a(new_n148), .b(new_n132), .c(new_n197), .o1(new_n198));
  nand03aa1n03x5               g103(.a(new_n163), .b(new_n166), .c(new_n171), .o1(new_n199));
  inv000aa1n02x5               g104(.a(new_n190), .o1(new_n200));
  aoi013aa1n06x4               g105(.a(new_n200), .b(new_n165), .c(new_n166), .d(new_n171), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n201), .b(new_n199), .c(new_n198), .d(new_n152), .o1(new_n202));
  norp02aa1n02x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  xorc02aa1n02x5               g108(.a(\a[17] ), .b(\b[16] ), .out0(new_n204));
  oaoi13aa1n06x5               g109(.a(new_n203), .b(new_n204), .c(new_n196), .d(new_n202), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[17] ), .c(new_n195), .out0(\s[18] ));
  nor042aa1n04x5               g111(.a(new_n150), .b(new_n199), .o1(new_n207));
  inv000aa1d42x5               g112(.a(\a[17] ), .o1(new_n208));
  xroi22aa1d06x4               g113(.a(new_n208), .b(\b[16] ), .c(new_n195), .d(\b[17] ), .out0(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n202), .c(new_n128), .d(new_n207), .o1(new_n210));
  oai022aa1d24x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  oaib12aa1n18x5               g116(.a(new_n211), .b(new_n195), .c(\b[17] ), .out0(new_n212));
  nor002aa1d32x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand42aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n210), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g122(.a(new_n213), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n215), .o1(new_n219));
  aoi012aa1n02x5               g124(.a(new_n219), .b(new_n210), .c(new_n212), .o1(new_n220));
  nor022aa1n06x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand42aa1n04x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanb02aa1n02x5               g127(.a(new_n221), .b(new_n222), .out0(new_n223));
  nano22aa1n02x4               g128(.a(new_n220), .b(new_n218), .c(new_n223), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n212), .o1(new_n225));
  oaoi13aa1n03x5               g130(.a(new_n225), .b(new_n209), .c(new_n196), .d(new_n202), .o1(new_n226));
  oaoi13aa1n03x5               g131(.a(new_n223), .b(new_n218), .c(new_n226), .d(new_n219), .o1(new_n227));
  norp02aa1n03x5               g132(.a(new_n227), .b(new_n224), .o1(\s[20] ));
  nona23aa1n09x5               g133(.a(new_n222), .b(new_n214), .c(new_n213), .d(new_n221), .out0(new_n229));
  norb02aa1n02x5               g134(.a(new_n209), .b(new_n229), .out0(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n202), .c(new_n128), .d(new_n207), .o1(new_n231));
  oaoi03aa1n02x5               g136(.a(\a[20] ), .b(\b[19] ), .c(new_n218), .o1(new_n232));
  oabi12aa1n18x5               g137(.a(new_n232), .b(new_n229), .c(new_n212), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .out0(new_n235));
  xobna2aa1n03x5               g140(.a(new_n235), .b(new_n231), .c(new_n234), .out0(\s[21] ));
  orn002aa1n03x5               g141(.a(\a[21] ), .b(\b[20] ), .o(new_n237));
  aoi012aa1n03x5               g142(.a(new_n235), .b(new_n231), .c(new_n234), .o1(new_n238));
  tech160nm_fixnrc02aa1n04x5   g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  nano22aa1n02x4               g144(.a(new_n238), .b(new_n237), .c(new_n239), .out0(new_n240));
  oaoi13aa1n03x5               g145(.a(new_n233), .b(new_n230), .c(new_n196), .d(new_n202), .o1(new_n241));
  oaoi13aa1n03x5               g146(.a(new_n239), .b(new_n237), .c(new_n241), .d(new_n235), .o1(new_n242));
  norp02aa1n03x5               g147(.a(new_n242), .b(new_n240), .o1(\s[22] ));
  nano23aa1n06x5               g148(.a(new_n213), .b(new_n221), .c(new_n222), .d(new_n214), .out0(new_n244));
  norp02aa1n12x5               g149(.a(new_n239), .b(new_n235), .o1(new_n245));
  nand23aa1n09x5               g150(.a(new_n209), .b(new_n245), .c(new_n244), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n202), .c(new_n128), .d(new_n207), .o1(new_n248));
  tech160nm_fioaoi03aa1n02p5x5 g153(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .o1(new_n249));
  tech160nm_fiaoi012aa1n02p5x5 g154(.a(new_n249), .b(new_n233), .c(new_n245), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  xnbna2aa1n03x5               g156(.a(new_n251), .b(new_n248), .c(new_n250), .out0(\s[23] ));
  inv000aa1d42x5               g157(.a(\a[23] ), .o1(new_n253));
  nanb02aa1n02x5               g158(.a(\b[22] ), .b(new_n253), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n251), .o1(new_n255));
  tech160nm_fiaoi012aa1n05x5   g160(.a(new_n255), .b(new_n248), .c(new_n250), .o1(new_n256));
  xorc02aa1n12x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  nano22aa1n03x7               g163(.a(new_n256), .b(new_n254), .c(new_n258), .out0(new_n259));
  inv000aa1n03x5               g164(.a(new_n250), .o1(new_n260));
  oaoi13aa1n03x5               g165(.a(new_n260), .b(new_n247), .c(new_n196), .d(new_n202), .o1(new_n261));
  oaoi13aa1n03x5               g166(.a(new_n258), .b(new_n254), .c(new_n261), .d(new_n255), .o1(new_n262));
  norp02aa1n03x5               g167(.a(new_n262), .b(new_n259), .o1(\s[24] ));
  and002aa1n12x5               g168(.a(new_n257), .b(new_n251), .o(new_n264));
  inv000aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  nano32aa1n02x4               g170(.a(new_n265), .b(new_n209), .c(new_n245), .d(new_n244), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n202), .c(new_n128), .d(new_n207), .o1(new_n267));
  nand23aa1d12x5               g172(.a(new_n233), .b(new_n245), .c(new_n264), .o1(new_n268));
  norp02aa1n02x5               g173(.a(\b[23] ), .b(\a[24] ), .o1(new_n269));
  aoi112aa1n02x5               g174(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n270));
  aoi113aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n249), .d(new_n257), .e(new_n251), .o1(new_n271));
  nand02aa1d10x5               g176(.a(new_n268), .b(new_n271), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  tech160nm_fixnrc02aa1n04x5   g178(.a(\b[24] ), .b(\a[25] ), .out0(new_n274));
  xobna2aa1n03x5               g179(.a(new_n274), .b(new_n267), .c(new_n273), .out0(\s[25] ));
  nor042aa1n03x5               g180(.a(\b[24] ), .b(\a[25] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoi012aa1n03x5               g182(.a(new_n274), .b(new_n267), .c(new_n273), .o1(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  nano22aa1n02x4               g184(.a(new_n278), .b(new_n277), .c(new_n279), .out0(new_n280));
  oaoi13aa1n03x5               g185(.a(new_n272), .b(new_n266), .c(new_n196), .d(new_n202), .o1(new_n281));
  oaoi13aa1n03x5               g186(.a(new_n279), .b(new_n277), .c(new_n281), .d(new_n274), .o1(new_n282));
  norp02aa1n03x5               g187(.a(new_n282), .b(new_n280), .o1(\s[26] ));
  nor042aa1n06x5               g188(.a(new_n279), .b(new_n274), .o1(new_n284));
  nano22aa1d15x5               g189(.a(new_n246), .b(new_n264), .c(new_n284), .out0(new_n285));
  aoai13aa1n12x5               g190(.a(new_n285), .b(new_n202), .c(new_n128), .d(new_n207), .o1(new_n286));
  oao003aa1n02x5               g191(.a(\a[26] ), .b(\b[25] ), .c(new_n277), .carry(new_n287));
  aobi12aa1n18x5               g192(.a(new_n287), .b(new_n272), .c(new_n284), .out0(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  xnbna2aa1n03x5               g194(.a(new_n289), .b(new_n288), .c(new_n286), .out0(\s[27] ));
  norp02aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o1(new_n291));
  inv040aa1n03x5               g196(.a(new_n291), .o1(new_n292));
  aobi12aa1n06x5               g197(.a(new_n289), .b(new_n288), .c(new_n286), .out0(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[27] ), .b(\a[28] ), .out0(new_n294));
  nano22aa1n03x7               g199(.a(new_n293), .b(new_n292), .c(new_n294), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n284), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n287), .b(new_n296), .c(new_n268), .d(new_n271), .o1(new_n297));
  aoai13aa1n02x5               g202(.a(new_n289), .b(new_n297), .c(new_n193), .d(new_n285), .o1(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n294), .b(new_n298), .c(new_n292), .o1(new_n299));
  norp02aa1n03x5               g204(.a(new_n299), .b(new_n295), .o1(\s[28] ));
  norb02aa1n02x5               g205(.a(new_n289), .b(new_n294), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n297), .c(new_n193), .d(new_n285), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  aoi012aa1n02x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  aobi12aa1n06x5               g210(.a(new_n301), .b(new_n288), .c(new_n286), .out0(new_n306));
  nano22aa1n03x7               g211(.a(new_n306), .b(new_n303), .c(new_n304), .out0(new_n307));
  norp02aa1n03x5               g212(.a(new_n305), .b(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g214(.a(new_n289), .b(new_n304), .c(new_n294), .out0(new_n310));
  aoai13aa1n02x5               g215(.a(new_n310), .b(new_n297), .c(new_n193), .d(new_n285), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[29] ), .b(\a[30] ), .out0(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n313), .b(new_n311), .c(new_n312), .o1(new_n314));
  aobi12aa1n06x5               g219(.a(new_n310), .b(new_n288), .c(new_n286), .out0(new_n315));
  nano22aa1n03x7               g220(.a(new_n315), .b(new_n312), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[30] ));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n310), .b(new_n313), .out0(new_n319));
  aobi12aa1n06x5               g224(.a(new_n319), .b(new_n288), .c(new_n286), .out0(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n321));
  nano22aa1n03x7               g226(.a(new_n320), .b(new_n318), .c(new_n321), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n319), .b(new_n297), .c(new_n193), .d(new_n285), .o1(new_n323));
  aoi012aa1n02x5               g228(.a(new_n318), .b(new_n323), .c(new_n321), .o1(new_n324));
  norp02aa1n03x5               g229(.a(new_n324), .b(new_n322), .o1(\s[31] ));
  xobna2aa1n03x5               g230(.a(new_n101), .b(new_n104), .c(new_n102), .out0(\s[3] ));
  norb02aa1n02x5               g231(.a(new_n105), .b(new_n106), .out0(new_n327));
  nanp02aa1n02x5               g232(.a(new_n104), .b(new_n102), .o1(new_n328));
  aoi012aa1n02x5               g233(.a(new_n99), .b(new_n328), .c(new_n100), .o1(new_n329));
  oai012aa1n02x5               g234(.a(new_n108), .b(new_n329), .c(new_n327), .o1(\s[4] ));
  nanb02aa1n02x5               g235(.a(new_n118), .b(new_n119), .out0(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n331), .b(new_n108), .c(new_n105), .out0(\s[5] ));
  nanb03aa1n02x5               g237(.a(new_n331), .b(new_n108), .c(new_n105), .out0(new_n333));
  obai22aa1n02x7               g238(.a(new_n333), .b(new_n118), .c(new_n180), .d(new_n117), .out0(new_n334));
  nona32aa1n02x4               g239(.a(new_n333), .b(new_n118), .c(new_n117), .d(new_n180), .out0(new_n335));
  nanp02aa1n02x5               g240(.a(new_n334), .b(new_n335), .o1(\s[6] ));
  xobna2aa1n03x5               g241(.a(new_n176), .b(new_n335), .c(new_n109), .out0(\s[7] ));
  nanp03aa1n02x5               g242(.a(new_n335), .b(new_n109), .c(new_n176), .o1(new_n338));
  xnbna2aa1n03x5               g243(.a(new_n177), .b(new_n338), .c(new_n111), .out0(\s[8] ));
  xobna2aa1n03x5               g244(.a(new_n135), .b(new_n121), .c(new_n127), .out0(\s[9] ));
endmodule


