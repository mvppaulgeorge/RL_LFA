// Benchmark "adder" written by ABC on Thu Jul 18 06:29:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n322, new_n323,
    new_n324, new_n325, new_n327, new_n329, new_n330, new_n331, new_n333,
    new_n335, new_n336, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1n08x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n12x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor002aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n06x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  oai012aa1n02x7               g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oai012aa1n12x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nand02aa1n06x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nor022aa1n06x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor022aa1n08x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n110), .b(new_n113), .c(new_n112), .d(new_n111), .out0(new_n114));
  tech160nm_fixnrc02aa1n05x5   g019(.a(\b[7] ), .b(\a[8] ), .out0(new_n115));
  nor022aa1n08x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nanb02aa1n02x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  nor043aa1n03x5               g023(.a(new_n114), .b(new_n115), .c(new_n118), .o1(new_n119));
  nanb03aa1n09x5               g024(.a(new_n116), .b(new_n117), .c(new_n110), .out0(new_n120));
  norp02aa1n04x5               g025(.a(new_n112), .b(new_n111), .o1(new_n121));
  aoi112aa1n02x5               g026(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n122));
  oab012aa1n02x4               g027(.a(new_n122), .b(\a[8] ), .c(\b[7] ), .out0(new_n123));
  oai013aa1d12x5               g028(.a(new_n123), .b(new_n120), .c(new_n115), .d(new_n121), .o1(new_n124));
  nand42aa1n03x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n97), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n127));
  norp02aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  nona23aa1n02x4               g035(.a(new_n127), .b(new_n129), .c(new_n128), .d(new_n97), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n130), .c(new_n98), .d(new_n127), .o1(\s[10] ));
  nano23aa1n06x5               g037(.a(new_n97), .b(new_n128), .c(new_n129), .d(new_n125), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n134));
  oaoi03aa1n12x5               g039(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nor002aa1n02x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand42aa1n10x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n134), .c(new_n136), .out0(\s[11] ));
  aobi12aa1n02x5               g045(.a(new_n139), .b(new_n134), .c(new_n136), .out0(new_n141));
  nand42aa1n20x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  inv030aa1n03x5               g047(.a(new_n142), .o1(new_n143));
  norp02aa1n02x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n144), .b(new_n142), .out0(new_n145));
  oai012aa1n02x5               g050(.a(new_n145), .b(new_n141), .c(new_n137), .o1(new_n146));
  oai022aa1n02x5               g051(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n147));
  oai013aa1n02x4               g052(.a(new_n146), .b(new_n143), .c(new_n141), .d(new_n147), .o1(\s[12] ));
  nano32aa1n03x7               g053(.a(new_n145), .b(new_n139), .c(new_n130), .d(new_n126), .out0(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n150));
  oai012aa1n02x5               g055(.a(new_n138), .b(\b[11] ), .c(\a[12] ), .o1(new_n151));
  nona32aa1n06x5               g056(.a(new_n135), .b(new_n151), .c(new_n143), .d(new_n137), .out0(new_n152));
  oaib12aa1n18x5               g057(.a(new_n152), .b(new_n143), .c(new_n147), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  nor022aa1n12x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n150), .c(new_n154), .out0(\s[13] ));
  inv000aa1d42x5               g063(.a(new_n155), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(new_n109), .b(new_n119), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n124), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(new_n160), .b(new_n161), .o1(new_n162));
  aoai13aa1n02x5               g067(.a(new_n157), .b(new_n153), .c(new_n162), .d(new_n149), .o1(new_n163));
  norp02aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  oai022aa1n02x5               g071(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n167));
  nanb03aa1n02x5               g072(.a(new_n167), .b(new_n163), .c(new_n165), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n166), .c(new_n159), .d(new_n163), .o1(\s[14] ));
  nano23aa1n06x5               g074(.a(new_n155), .b(new_n164), .c(new_n165), .d(new_n156), .out0(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n153), .c(new_n162), .d(new_n149), .o1(new_n171));
  oai012aa1n02x5               g076(.a(new_n165), .b(new_n164), .c(new_n155), .o1(new_n172));
  nor022aa1n08x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  xobna2aa1n03x5               g080(.a(new_n175), .b(new_n171), .c(new_n172), .out0(\s[15] ));
  nona23aa1n02x4               g081(.a(new_n165), .b(new_n156), .c(new_n155), .d(new_n164), .out0(new_n177));
  aoai13aa1n02x7               g082(.a(new_n172), .b(new_n177), .c(new_n150), .d(new_n154), .o1(new_n178));
  nor022aa1n06x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanp02aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n173), .c(new_n178), .d(new_n174), .o1(new_n182));
  nor042aa1n04x5               g087(.a(new_n179), .b(new_n173), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n180), .b(new_n175), .c(new_n171), .d(new_n172), .o1(new_n185));
  oai012aa1n02x5               g090(.a(new_n182), .b(new_n185), .c(new_n184), .o1(\s[16] ));
  nano23aa1n02x5               g091(.a(new_n137), .b(new_n144), .c(new_n142), .d(new_n138), .out0(new_n187));
  nano23aa1n06x5               g092(.a(new_n173), .b(new_n179), .c(new_n180), .d(new_n174), .out0(new_n188));
  nand02aa1n02x5               g093(.a(new_n188), .b(new_n170), .o1(new_n189));
  nano22aa1n02x5               g094(.a(new_n189), .b(new_n133), .c(new_n187), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n191));
  nor043aa1n02x5               g096(.a(new_n177), .b(new_n175), .c(new_n181), .o1(new_n192));
  nanb03aa1n02x5               g097(.a(new_n179), .b(new_n180), .c(new_n174), .out0(new_n193));
  oai112aa1n02x5               g098(.a(new_n167), .b(new_n165), .c(\b[14] ), .d(\a[15] ), .o1(new_n194));
  obai22aa1n09x5               g099(.a(new_n180), .b(new_n183), .c(new_n194), .d(new_n193), .out0(new_n195));
  aoi012aa1d18x5               g100(.a(new_n195), .b(new_n153), .c(new_n192), .o1(new_n196));
  tech160nm_finor002aa1n05x5   g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nand42aa1d28x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n191), .c(new_n196), .out0(\s[17] ));
  nanp02aa1n09x5               g105(.a(new_n191), .b(new_n196), .o1(new_n201));
  aoi012aa1n02x5               g106(.a(new_n197), .b(new_n201), .c(new_n198), .o1(new_n202));
  norp02aa1n04x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand42aa1d28x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  oaih22aa1n06x5               g110(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n206));
  aoi122aa1n06x5               g111(.a(new_n206), .b(\b[17] ), .c(\a[18] ), .d(new_n201), .e(new_n199), .o1(new_n207));
  oabi12aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n205), .out0(\s[18] ));
  nano23aa1d15x5               g113(.a(new_n197), .b(new_n203), .c(new_n204), .d(new_n198), .out0(new_n209));
  nand22aa1n03x5               g114(.a(new_n201), .b(new_n209), .o1(new_n210));
  oai012aa1n02x5               g115(.a(new_n204), .b(new_n203), .c(new_n197), .o1(new_n211));
  norp02aa1n02x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nand42aa1n03x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  norb02aa1n09x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  xnbna2aa1n03x5               g119(.a(new_n214), .b(new_n210), .c(new_n211), .out0(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g121(.a(new_n209), .o1(new_n217));
  aoai13aa1n02x7               g122(.a(new_n211), .b(new_n217), .c(new_n191), .d(new_n196), .o1(new_n218));
  orn002aa1n02x7               g123(.a(\a[20] ), .b(\b[19] ), .o(new_n219));
  nand22aa1n03x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(new_n219), .b(new_n220), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n212), .c(new_n218), .d(new_n213), .o1(new_n222));
  oai022aa1n02x5               g127(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n214), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n220), .b(new_n224), .c(new_n210), .d(new_n211), .o1(new_n225));
  oai012aa1n03x5               g130(.a(new_n222), .b(new_n225), .c(new_n223), .o1(\s[20] ));
  nanb03aa1d24x5               g131(.a(new_n221), .b(new_n209), .c(new_n214), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  nanp03aa1n02x5               g133(.a(new_n219), .b(new_n213), .c(new_n220), .o1(new_n229));
  oai112aa1n02x5               g134(.a(new_n206), .b(new_n204), .c(\b[18] ), .d(\a[19] ), .o1(new_n230));
  nanp02aa1n02x5               g135(.a(new_n223), .b(new_n220), .o1(new_n231));
  tech160nm_fioai012aa1n04x5   g136(.a(new_n231), .b(new_n230), .c(new_n229), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[21] ), .b(\b[20] ), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n232), .c(new_n201), .d(new_n228), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n233), .b(new_n232), .c(new_n201), .d(new_n228), .o1(new_n235));
  norb02aa1n03x4               g140(.a(new_n234), .b(new_n235), .out0(\s[21] ));
  inv000aa1d42x5               g141(.a(\a[21] ), .o1(new_n237));
  nanb02aa1n02x5               g142(.a(\b[20] ), .b(new_n237), .out0(new_n238));
  xorc02aa1n02x5               g143(.a(\a[22] ), .b(\b[21] ), .out0(new_n239));
  and002aa1n02x5               g144(.a(\b[21] ), .b(\a[22] ), .o(new_n240));
  oai022aa1n02x5               g145(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n241));
  nona22aa1n02x5               g146(.a(new_n234), .b(new_n240), .c(new_n241), .out0(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n239), .c(new_n238), .d(new_n234), .o1(\s[22] ));
  inv000aa1d42x5               g148(.a(\a[22] ), .o1(new_n244));
  xroi22aa1d04x5               g149(.a(new_n237), .b(\b[20] ), .c(new_n244), .d(\b[21] ), .out0(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n227), .out0(new_n246));
  oaoi03aa1n02x5               g151(.a(\a[22] ), .b(\b[21] ), .c(new_n238), .o1(new_n247));
  tech160nm_fiao0012aa1n02p5x5 g152(.a(new_n247), .b(new_n232), .c(new_n245), .o(new_n248));
  xorc02aa1n12x5               g153(.a(\a[23] ), .b(\b[22] ), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n248), .c(new_n201), .d(new_n246), .o1(new_n250));
  aoi112aa1n02x5               g155(.a(new_n249), .b(new_n248), .c(new_n201), .d(new_n246), .o1(new_n251));
  norb02aa1n03x4               g156(.a(new_n250), .b(new_n251), .out0(\s[23] ));
  norp02aa1n02x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[24] ), .b(\b[23] ), .out0(new_n255));
  and002aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o(new_n256));
  oai022aa1n02x5               g161(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n257));
  nona22aa1n02x5               g162(.a(new_n250), .b(new_n256), .c(new_n257), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n255), .c(new_n254), .d(new_n250), .o1(\s[24] ));
  nano32aa1n02x5               g164(.a(new_n227), .b(new_n255), .c(new_n245), .d(new_n249), .out0(new_n260));
  aob012aa1n02x5               g165(.a(new_n257), .b(\b[23] ), .c(\a[24] ), .out0(new_n261));
  and002aa1n02x5               g166(.a(new_n255), .b(new_n249), .o(new_n262));
  aoai13aa1n06x5               g167(.a(new_n262), .b(new_n247), .c(new_n232), .d(new_n245), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(new_n263), .b(new_n261), .o1(new_n264));
  xnrc02aa1n12x5               g169(.a(\b[24] ), .b(\a[25] ), .out0(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n264), .c(new_n201), .d(new_n260), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n266), .b(new_n264), .c(new_n201), .d(new_n260), .o1(new_n268));
  norb02aa1n02x5               g173(.a(new_n267), .b(new_n268), .out0(\s[25] ));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  tech160nm_fixorc02aa1n04x5   g176(.a(\a[26] ), .b(\b[25] ), .out0(new_n272));
  and002aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .o(new_n273));
  oai022aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n274));
  nona22aa1n02x5               g179(.a(new_n267), .b(new_n273), .c(new_n274), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n272), .c(new_n271), .d(new_n267), .o1(\s[26] ));
  nanb02aa1n09x5               g181(.a(new_n265), .b(new_n272), .out0(new_n277));
  nona23aa1n09x5               g182(.a(new_n245), .b(new_n262), .c(new_n227), .d(new_n277), .out0(new_n278));
  nanb02aa1n06x5               g183(.a(new_n278), .b(new_n201), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n277), .o1(new_n280));
  aob012aa1n02x5               g185(.a(new_n274), .b(\b[25] ), .c(\a[26] ), .out0(new_n281));
  aobi12aa1n02x5               g186(.a(new_n281), .b(new_n264), .c(new_n280), .out0(new_n282));
  xorc02aa1n02x5               g187(.a(\a[27] ), .b(\b[26] ), .out0(new_n283));
  xnbna2aa1n03x5               g188(.a(new_n283), .b(new_n282), .c(new_n279), .out0(\s[27] ));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  aoi012aa1n06x5               g191(.a(new_n278), .b(new_n191), .c(new_n196), .o1(new_n287));
  aoai13aa1n06x5               g192(.a(new_n281), .b(new_n277), .c(new_n263), .d(new_n261), .o1(new_n288));
  oaih12aa1n02x5               g193(.a(new_n283), .b(new_n288), .c(new_n287), .o1(new_n289));
  xorc02aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .out0(new_n290));
  oai022aa1n02x5               g195(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n291));
  aoi012aa1n02x5               g196(.a(new_n291), .b(\a[28] ), .c(\b[27] ), .o1(new_n292));
  tech160nm_finand02aa1n03p5x5 g197(.a(new_n289), .b(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n289), .d(new_n286), .o1(\s[28] ));
  xorc02aa1n02x5               g199(.a(\a[29] ), .b(\b[28] ), .out0(new_n295));
  and002aa1n02x5               g200(.a(new_n290), .b(new_n283), .o(new_n296));
  inv000aa1d42x5               g201(.a(\b[27] ), .o1(new_n297));
  oaib12aa1n09x5               g202(.a(new_n291), .b(new_n297), .c(\a[28] ), .out0(new_n298));
  inv000aa1d42x5               g203(.a(new_n298), .o1(new_n299));
  oaoi13aa1n03x5               g204(.a(new_n299), .b(new_n296), .c(new_n288), .d(new_n287), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n295), .o1(new_n301));
  oaih12aa1n02x5               g206(.a(new_n296), .b(new_n288), .c(new_n287), .o1(new_n302));
  nona22aa1n02x5               g207(.a(new_n302), .b(new_n299), .c(new_n301), .out0(new_n303));
  oai012aa1n03x5               g208(.a(new_n303), .b(new_n300), .c(new_n295), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g210(.a(new_n301), .b(new_n283), .c(new_n290), .out0(new_n306));
  oaoi03aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .o1(new_n307));
  oaoi13aa1n03x5               g212(.a(new_n307), .b(new_n306), .c(new_n288), .d(new_n287), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .out0(new_n309));
  oaih12aa1n02x5               g214(.a(new_n306), .b(new_n288), .c(new_n287), .o1(new_n310));
  norb02aa1n02x5               g215(.a(new_n309), .b(new_n307), .out0(new_n311));
  tech160nm_finand02aa1n03p5x5 g216(.a(new_n310), .b(new_n311), .o1(new_n312));
  oai012aa1n03x5               g217(.a(new_n312), .b(new_n308), .c(new_n309), .o1(\s[30] ));
  nano32aa1n02x4               g218(.a(new_n301), .b(new_n309), .c(new_n283), .d(new_n290), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n314), .b(new_n288), .c(new_n287), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n316));
  xorc02aa1n02x5               g221(.a(\a[31] ), .b(\b[30] ), .out0(new_n317));
  oai012aa1n02x5               g222(.a(new_n317), .b(\b[29] ), .c(\a[30] ), .o1(new_n318));
  aoi012aa1n02x5               g223(.a(new_n318), .b(new_n307), .c(new_n309), .o1(new_n319));
  nand42aa1n02x5               g224(.a(new_n315), .b(new_n319), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n317), .c(new_n315), .d(new_n316), .o1(\s[31] ));
  aoi022aa1n02x5               g226(.a(new_n100), .b(new_n99), .c(\a[1] ), .d(\b[0] ), .o1(new_n322));
  oaib12aa1n02x5               g227(.a(new_n322), .b(new_n100), .c(\a[2] ), .out0(new_n323));
  norb02aa1n02x5               g228(.a(new_n106), .b(new_n105), .out0(new_n324));
  aboi22aa1n03x5               g229(.a(new_n105), .b(new_n106), .c(new_n99), .d(new_n100), .out0(new_n325));
  aboi22aa1n03x5               g230(.a(new_n102), .b(new_n324), .c(new_n325), .d(new_n323), .out0(\s[3] ));
  oaoi03aa1n02x5               g231(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  inv000aa1d42x5               g233(.a(new_n102), .o1(new_n329));
  nanb02aa1n02x5               g234(.a(new_n107), .b(new_n329), .out0(new_n330));
  nanb02aa1n02x5               g235(.a(new_n112), .b(new_n113), .out0(new_n331));
  xobna2aa1n03x5               g236(.a(new_n331), .b(new_n330), .c(new_n108), .out0(\s[5] ));
  aoi012aa1n02x5               g237(.a(new_n112), .b(new_n109), .c(new_n113), .o1(new_n333));
  xnrb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g239(.a(new_n114), .b(new_n109), .out0(new_n335));
  oaib12aa1n02x5               g240(.a(new_n335), .b(new_n121), .c(new_n110), .out0(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g242(.a(new_n116), .b(new_n336), .c(new_n117), .o1(new_n338));
  xnrb03aa1n02x5               g243(.a(new_n338), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g244(.a(new_n126), .b(new_n160), .c(new_n161), .out0(\s[9] ));
endmodule


