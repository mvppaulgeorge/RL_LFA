// Benchmark "adder" written by ABC on Thu Jul 18 03:12:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n341, new_n342, new_n344, new_n347,
    new_n348, new_n349, new_n352, new_n354, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  and002aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n09x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  nand42aa1n03x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norb02aa1n03x4               g007(.a(new_n101), .b(new_n102), .out0(new_n103));
  xorc02aa1n12x5               g008(.a(\a[3] ), .b(\b[2] ), .out0(new_n104));
  nanp03aa1n04x5               g009(.a(new_n100), .b(new_n104), .c(new_n103), .o1(new_n105));
  norp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  aoi012aa1n02x7               g011(.a(new_n102), .b(new_n106), .c(new_n101), .o1(new_n107));
  nand42aa1n02x5               g012(.a(new_n105), .b(new_n107), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nand42aa1n04x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  norb02aa1n02x7               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  nor002aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  norb02aa1n06x4               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  tech160nm_fixorc02aa1n05x5   g019(.a(\a[8] ), .b(\b[7] ), .out0(new_n115));
  nand42aa1n03x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor022aa1n06x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  norb02aa1n09x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  inv000aa1d42x5               g023(.a(new_n118), .o1(new_n119));
  nano32aa1n03x7               g024(.a(new_n119), .b(new_n115), .c(new_n114), .d(new_n111), .out0(new_n120));
  nano22aa1n03x5               g025(.a(new_n117), .b(new_n110), .c(new_n116), .out0(new_n121));
  oai022aa1n02x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  nanp03aa1n02x5               g027(.a(new_n121), .b(new_n115), .c(new_n122), .o1(new_n123));
  inv000aa1n02x5               g028(.a(new_n117), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  nanb02aa1n02x5               g030(.a(new_n125), .b(new_n123), .out0(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n126), .c(new_n108), .d(new_n120), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  oai022aa1d24x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nand42aa1n03x5               g037(.a(new_n128), .b(new_n132), .o1(new_n133));
  nand42aa1n02x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nand42aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor042aa1n09x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb03aa1n02x5               g041(.a(new_n136), .b(new_n134), .c(new_n135), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n136), .o1(new_n138));
  aoi022aa1n02x5               g043(.a(new_n133), .b(new_n134), .c(new_n138), .d(new_n135), .o1(new_n139));
  aoib12aa1n02x5               g044(.a(new_n139), .b(new_n133), .c(new_n137), .out0(\s[11] ));
  nor042aa1n06x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1n03x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  aoi113aa1n02x5               g048(.a(new_n143), .b(new_n136), .c(new_n133), .d(new_n135), .e(new_n134), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n138), .b(new_n137), .c(new_n128), .d(new_n132), .o1(new_n145));
  aoi012aa1n02x5               g050(.a(new_n144), .b(new_n143), .c(new_n145), .o1(\s[12] ));
  nano23aa1n09x5               g051(.a(new_n141), .b(new_n136), .c(new_n142), .d(new_n135), .out0(new_n147));
  nanp03aa1d12x5               g052(.a(new_n147), .b(new_n127), .c(new_n129), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n126), .c(new_n108), .d(new_n120), .o1(new_n150));
  aoi022aa1n06x5               g055(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n151));
  aoai13aa1n12x5               g056(.a(new_n151), .b(new_n136), .c(new_n131), .d(new_n134), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  nona22aa1n02x4               g058(.a(new_n150), .b(new_n153), .c(new_n141), .out0(new_n154));
  xnrc02aa1n12x5               g059(.a(\b[12] ), .b(\a[13] ), .out0(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n141), .o1(new_n157));
  nano22aa1n02x4               g062(.a(new_n153), .b(new_n157), .c(new_n155), .out0(new_n158));
  aoi022aa1n02x5               g063(.a(new_n154), .b(new_n156), .c(new_n150), .d(new_n158), .o1(\s[13] ));
  orn002aa1n02x5               g064(.a(\a[13] ), .b(\b[12] ), .o(new_n160));
  nano23aa1n02x5               g065(.a(new_n109), .b(new_n112), .c(new_n113), .d(new_n110), .out0(new_n161));
  nanp03aa1n03x5               g066(.a(new_n161), .b(new_n115), .c(new_n118), .o1(new_n162));
  aoi013aa1n03x5               g067(.a(new_n125), .b(new_n121), .c(new_n115), .d(new_n122), .o1(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n162), .c(new_n105), .d(new_n107), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(new_n152), .b(new_n157), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n156), .b(new_n165), .c(new_n164), .d(new_n149), .o1(new_n166));
  xnrc02aa1n03x5               g071(.a(\b[13] ), .b(\a[14] ), .out0(new_n167));
  xobna2aa1n03x5               g072(.a(new_n167), .b(new_n166), .c(new_n160), .out0(\s[14] ));
  norp02aa1n04x5               g073(.a(new_n167), .b(new_n155), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n165), .c(new_n164), .d(new_n149), .o1(new_n170));
  oaoi03aa1n02x5               g075(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  xnrc02aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n172), .out0(\s[15] ));
  aob012aa1n02x5               g080(.a(new_n174), .b(new_n170), .c(new_n172), .out0(new_n176));
  tech160nm_fixnrc02aa1n02p5x5 g081(.a(\b[15] ), .b(\a[16] ), .out0(new_n177));
  orn002aa1n02x5               g082(.a(\a[15] ), .b(\b[14] ), .o(new_n178));
  and002aa1n02x5               g083(.a(new_n177), .b(new_n178), .o(new_n179));
  aoai13aa1n02x5               g084(.a(new_n178), .b(new_n173), .c(new_n170), .d(new_n172), .o1(new_n180));
  aboi22aa1n03x5               g085(.a(new_n177), .b(new_n180), .c(new_n176), .d(new_n179), .out0(\s[16] ));
  nor042aa1n02x5               g086(.a(new_n177), .b(new_n173), .o1(new_n182));
  nano22aa1n12x5               g087(.a(new_n148), .b(new_n169), .c(new_n182), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n126), .c(new_n108), .d(new_n120), .o1(new_n184));
  nand02aa1n02x5               g089(.a(new_n182), .b(new_n169), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[14] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[13] ), .o1(new_n187));
  nor042aa1n02x5               g092(.a(\b[12] ), .b(\a[13] ), .o1(new_n188));
  aoi022aa1d24x5               g093(.a(\b[14] ), .b(\a[15] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n188), .c(new_n186), .d(new_n187), .o1(new_n190));
  oa0022aa1n06x5               g095(.a(\a[16] ), .b(\b[15] ), .c(\a[15] ), .d(\b[14] ), .o(new_n191));
  aoi022aa1n06x5               g096(.a(new_n190), .b(new_n191), .c(\b[15] ), .d(\a[16] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  aoai13aa1n12x5               g098(.a(new_n193), .b(new_n185), .c(new_n157), .d(new_n152), .o1(new_n194));
  nanb02aa1n12x5               g099(.a(new_n194), .b(new_n184), .out0(new_n195));
  xorc02aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  aoi113aa1n02x5               g101(.a(new_n192), .b(new_n196), .c(new_n165), .d(new_n169), .e(new_n182), .o1(new_n197));
  aoi022aa1n02x5               g102(.a(new_n195), .b(new_n196), .c(new_n184), .d(new_n197), .o1(\s[17] ));
  nor042aa1n09x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n199), .o1(new_n200));
  aoai13aa1n03x5               g105(.a(new_n196), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n201));
  nor002aa1n03x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand02aa1n03x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norb02aa1n06x4               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n201), .c(new_n200), .out0(\s[18] ));
  and002aa1n02x5               g110(.a(new_n196), .b(new_n204), .o(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n207));
  oaoi03aa1n02x5               g112(.a(\a[18] ), .b(\b[17] ), .c(new_n200), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  nor042aa1n09x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nand02aa1d04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  norb02aa1n12x5               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n207), .c(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g119(.a(new_n212), .b(new_n207), .c(new_n209), .out0(new_n215));
  nor042aa1n06x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand22aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1n06x4               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  inv000aa1d42x5               g123(.a(\a[19] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(\b[18] ), .o1(new_n220));
  aboi22aa1n03x5               g125(.a(new_n216), .b(new_n217), .c(new_n219), .d(new_n220), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n210), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n212), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n222), .b(new_n223), .c(new_n207), .d(new_n209), .o1(new_n224));
  aoi022aa1n02x5               g129(.a(new_n224), .b(new_n218), .c(new_n215), .d(new_n221), .o1(\s[20] ));
  nano32aa1n03x7               g130(.a(new_n223), .b(new_n196), .c(new_n218), .d(new_n204), .out0(new_n226));
  aoai13aa1n02x5               g131(.a(new_n226), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n227));
  nanb03aa1n12x5               g132(.a(new_n216), .b(new_n217), .c(new_n211), .out0(new_n228));
  oai112aa1n06x5               g133(.a(new_n222), .b(new_n203), .c(new_n202), .d(new_n199), .o1(new_n229));
  aoi012aa1n12x5               g134(.a(new_n216), .b(new_n210), .c(new_n217), .o1(new_n230));
  oai012aa1d24x5               g135(.a(new_n230), .b(new_n229), .c(new_n228), .o1(new_n231));
  nor042aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nand42aa1n02x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1d21x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n231), .c(new_n195), .d(new_n226), .o1(new_n235));
  nano22aa1n12x5               g140(.a(new_n216), .b(new_n211), .c(new_n217), .out0(new_n236));
  oai012aa1n02x5               g141(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .o1(new_n237));
  oab012aa1n02x5               g142(.a(new_n237), .b(new_n199), .c(new_n202), .out0(new_n238));
  inv030aa1n02x5               g143(.a(new_n230), .o1(new_n239));
  aoi112aa1n02x5               g144(.a(new_n239), .b(new_n234), .c(new_n238), .d(new_n236), .o1(new_n240));
  aobi12aa1n03x7               g145(.a(new_n235), .b(new_n240), .c(new_n227), .out0(\s[21] ));
  nor042aa1n02x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  nand22aa1n04x5               g147(.a(\b[21] ), .b(\a[22] ), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n243), .b(new_n242), .out0(new_n244));
  aoib12aa1n02x5               g149(.a(new_n232), .b(new_n243), .c(new_n242), .out0(new_n245));
  inv000aa1d42x5               g150(.a(new_n231), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n232), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n234), .o1(new_n248));
  aoai13aa1n02x7               g153(.a(new_n247), .b(new_n248), .c(new_n227), .d(new_n246), .o1(new_n249));
  aoi022aa1n02x7               g154(.a(new_n249), .b(new_n244), .c(new_n235), .d(new_n245), .o1(\s[22] ));
  inv020aa1n02x5               g155(.a(new_n226), .o1(new_n251));
  nano22aa1n02x5               g156(.a(new_n251), .b(new_n234), .c(new_n244), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n253));
  nano23aa1n06x5               g158(.a(new_n232), .b(new_n242), .c(new_n243), .d(new_n233), .out0(new_n254));
  aoi012aa1d18x5               g159(.a(new_n242), .b(new_n232), .c(new_n243), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoi012aa1n02x5               g161(.a(new_n256), .b(new_n231), .c(new_n254), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[23] ), .b(\b[22] ), .out0(new_n258));
  aob012aa1n03x5               g163(.a(new_n258), .b(new_n253), .c(new_n257), .out0(new_n259));
  aoi112aa1n02x5               g164(.a(new_n258), .b(new_n256), .c(new_n231), .d(new_n254), .o1(new_n260));
  aobi12aa1n02x7               g165(.a(new_n259), .b(new_n260), .c(new_n253), .out0(\s[23] ));
  tech160nm_fixorc02aa1n02p5x5 g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  nor042aa1n06x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  norp02aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n263), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n258), .o1(new_n266));
  aoai13aa1n02x5               g171(.a(new_n265), .b(new_n266), .c(new_n253), .d(new_n257), .o1(new_n267));
  aoi022aa1n02x7               g172(.a(new_n267), .b(new_n262), .c(new_n259), .d(new_n264), .o1(\s[24] ));
  and002aa1n18x5               g173(.a(new_n262), .b(new_n258), .o(new_n269));
  nano22aa1n02x5               g174(.a(new_n251), .b(new_n269), .c(new_n254), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n254), .b(new_n239), .c(new_n238), .d(new_n236), .o1(new_n272));
  inv030aa1n02x5               g177(.a(new_n269), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[24] ), .b(\b[23] ), .c(new_n265), .carry(new_n274));
  aoai13aa1n12x5               g179(.a(new_n274), .b(new_n273), .c(new_n272), .d(new_n255), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  aob012aa1n03x5               g182(.a(new_n277), .b(new_n271), .c(new_n276), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n269), .b(new_n256), .c(new_n231), .d(new_n254), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n277), .o1(new_n280));
  and003aa1n02x5               g185(.a(new_n279), .b(new_n280), .c(new_n274), .o(new_n281));
  aobi12aa1n02x7               g186(.a(new_n278), .b(new_n281), .c(new_n271), .out0(\s[25] ));
  xorc02aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .out0(new_n283));
  nor042aa1n03x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  norp02aa1n02x5               g189(.a(new_n283), .b(new_n284), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n284), .o1(new_n286));
  aoai13aa1n02x5               g191(.a(new_n286), .b(new_n280), .c(new_n271), .d(new_n276), .o1(new_n287));
  aoi022aa1n02x7               g192(.a(new_n287), .b(new_n283), .c(new_n278), .d(new_n285), .o1(\s[26] ));
  and002aa1n12x5               g193(.a(new_n283), .b(new_n277), .o(new_n289));
  nano32aa1d12x5               g194(.a(new_n251), .b(new_n289), .c(new_n254), .d(new_n269), .out0(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n194), .c(new_n164), .d(new_n183), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n289), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .c(new_n286), .carry(new_n293));
  aoai13aa1n04x5               g198(.a(new_n293), .b(new_n292), .c(new_n279), .d(new_n274), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n294), .c(new_n195), .d(new_n290), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n293), .o1(new_n297));
  aoi112aa1n02x5               g202(.a(new_n295), .b(new_n297), .c(new_n275), .d(new_n289), .o1(new_n298));
  aobi12aa1n03x7               g203(.a(new_n296), .b(new_n298), .c(new_n291), .out0(\s[27] ));
  xorc02aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .out0(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  norp02aa1n02x5               g206(.a(new_n300), .b(new_n301), .o1(new_n302));
  aoi012aa1n09x5               g207(.a(new_n297), .b(new_n275), .c(new_n289), .o1(new_n303));
  inv000aa1n03x5               g208(.a(new_n301), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n295), .o1(new_n305));
  aoai13aa1n02x7               g210(.a(new_n304), .b(new_n305), .c(new_n303), .d(new_n291), .o1(new_n306));
  aoi022aa1n02x7               g211(.a(new_n306), .b(new_n300), .c(new_n296), .d(new_n302), .o1(\s[28] ));
  and002aa1n02x5               g212(.a(new_n300), .b(new_n295), .o(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n294), .c(new_n195), .d(new_n290), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n308), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n311));
  aoai13aa1n02x7               g216(.a(new_n311), .b(new_n310), .c(new_n303), .d(new_n291), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n311), .b(new_n313), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[29] ));
  xnrb03aa1n02x5               g220(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g221(.a(new_n305), .b(new_n300), .c(new_n313), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n294), .c(new_n195), .d(new_n290), .o1(new_n318));
  inv000aa1n02x5               g223(.a(new_n317), .o1(new_n319));
  inv000aa1d42x5               g224(.a(\b[28] ), .o1(new_n320));
  inv000aa1d42x5               g225(.a(\a[29] ), .o1(new_n321));
  oaib12aa1n02x5               g226(.a(new_n311), .b(\b[28] ), .c(new_n321), .out0(new_n322));
  oaib12aa1n02x5               g227(.a(new_n322), .b(new_n320), .c(\a[29] ), .out0(new_n323));
  aoai13aa1n03x5               g228(.a(new_n323), .b(new_n319), .c(new_n303), .d(new_n291), .o1(new_n324));
  xorc02aa1n02x5               g229(.a(\a[30] ), .b(\b[29] ), .out0(new_n325));
  oaoi13aa1n02x5               g230(.a(new_n325), .b(new_n322), .c(new_n321), .d(new_n320), .o1(new_n326));
  aoi022aa1n03x5               g231(.a(new_n324), .b(new_n325), .c(new_n318), .d(new_n326), .o1(\s[30] ));
  nano32aa1n06x5               g232(.a(new_n305), .b(new_n325), .c(new_n300), .d(new_n313), .out0(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n294), .c(new_n195), .d(new_n290), .o1(new_n329));
  aoi022aa1n02x5               g234(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n330));
  norb02aa1n02x5               g235(.a(\b[30] ), .b(\a[31] ), .out0(new_n331));
  obai22aa1n02x7               g236(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n332));
  aoi112aa1n02x5               g237(.a(new_n332), .b(new_n331), .c(new_n322), .d(new_n330), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  inv000aa1d42x5               g239(.a(new_n328), .o1(new_n335));
  norp02aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .o1(new_n336));
  aoi012aa1n02x5               g241(.a(new_n336), .b(new_n322), .c(new_n330), .o1(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n335), .c(new_n303), .d(new_n291), .o1(new_n338));
  aoi022aa1n03x5               g243(.a(new_n338), .b(new_n334), .c(new_n329), .d(new_n333), .o1(\s[31] ));
  orn002aa1n02x5               g244(.a(\a[2] ), .b(\b[1] ), .o(new_n340));
  nanp02aa1n02x5               g245(.a(\b[1] ), .b(\a[2] ), .o1(new_n341));
  nanb03aa1n02x5               g246(.a(new_n99), .b(new_n340), .c(new_n341), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n104), .b(new_n342), .c(new_n340), .out0(\s[3] ));
  aoi112aa1n02x5               g248(.a(new_n106), .b(new_n103), .c(new_n100), .d(new_n104), .o1(new_n344));
  oaoi13aa1n02x5               g249(.a(new_n344), .b(new_n108), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g250(.a(new_n114), .b(new_n105), .c(new_n107), .out0(\s[5] ));
  aoi012aa1n02x5               g251(.a(new_n112), .b(new_n108), .c(new_n113), .o1(new_n347));
  norb03aa1n02x5               g252(.a(new_n110), .b(new_n109), .c(new_n112), .out0(new_n348));
  aob012aa1n02x5               g253(.a(new_n348), .b(new_n108), .c(new_n114), .out0(new_n349));
  oai012aa1n02x5               g254(.a(new_n349), .b(new_n347), .c(new_n111), .o1(\s[6] ));
  xnbna2aa1n03x5               g255(.a(new_n119), .b(new_n349), .c(new_n110), .out0(\s[7] ));
  nanp02aa1n02x5               g256(.a(new_n349), .b(new_n121), .o1(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n115), .b(new_n352), .c(new_n124), .out0(\s[8] ));
  nanp02aa1n02x5               g258(.a(new_n108), .b(new_n120), .o1(new_n354));
  aoi113aa1n02x5               g259(.a(new_n127), .b(new_n125), .c(new_n121), .d(new_n115), .e(new_n122), .o1(new_n355));
  aoi022aa1n02x5               g260(.a(new_n164), .b(new_n127), .c(new_n354), .d(new_n355), .o1(\s[9] ));
endmodule


