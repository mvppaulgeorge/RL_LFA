// Benchmark "adder" written by ABC on Wed Jul 17 15:32:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n375, new_n377, new_n379, new_n380, new_n382,
    new_n383, new_n385, new_n386, new_n387, new_n388, new_n389, new_n391,
    new_n392, new_n394, new_n395;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n04x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  inv000aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nand22aa1n03x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1d06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n02x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .out0(new_n101));
  nor042aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand22aa1n12x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n02x7               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor042aa1n09x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n16x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n02x7               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nand23aa1n04x5               g012(.a(new_n101), .b(new_n104), .c(new_n107), .o1(new_n108));
  aoi012aa1n06x5               g013(.a(new_n102), .b(new_n105), .c(new_n103), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  norb02aa1n03x5               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  nor002aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand42aa1n06x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  norb02aa1n06x4               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  nor002aa1d32x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand02aa1d28x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor042aa1n09x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand02aa1n08x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nand23aa1n02x5               g025(.a(new_n120), .b(new_n112), .c(new_n115), .o1(new_n121));
  inv040aa1n08x5               g026(.a(new_n110), .o1(new_n122));
  oaoi03aa1n12x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  tech160nm_fiao0012aa1n02p5x5 g028(.a(new_n116), .b(new_n118), .c(new_n117), .o(new_n124));
  aoi012aa1d24x5               g029(.a(new_n124), .b(new_n120), .c(new_n123), .o1(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n121), .c(new_n108), .d(new_n109), .o1(new_n126));
  nor042aa1n06x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nand42aa1n03x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nor042aa1n06x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand02aa1n06x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n127), .c(new_n126), .d(new_n128), .o1(new_n133));
  nona22aa1n02x4               g038(.a(new_n131), .b(new_n130), .c(new_n127), .out0(new_n134));
  aoai13aa1n02x5               g039(.a(new_n133), .b(new_n134), .c(new_n129), .d(new_n126), .o1(\s[10] ));
  nano23aa1d15x5               g040(.a(new_n127), .b(new_n130), .c(new_n131), .d(new_n128), .out0(new_n136));
  aoi012aa1n06x5               g041(.a(new_n130), .b(new_n127), .c(new_n131), .o1(new_n137));
  inv030aa1n06x5               g042(.a(new_n137), .o1(new_n138));
  nor002aa1n20x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nanp02aa1n04x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  aoai13aa1n06x5               g046(.a(new_n141), .b(new_n138), .c(new_n126), .d(new_n136), .o1(new_n142));
  aoi112aa1n02x5               g047(.a(new_n141), .b(new_n130), .c(new_n131), .d(new_n127), .o1(new_n143));
  aobi12aa1n02x5               g048(.a(new_n143), .b(new_n126), .c(new_n136), .out0(new_n144));
  norb02aa1n02x5               g049(.a(new_n142), .b(new_n144), .out0(\s[11] ));
  inv000aa1d42x5               g050(.a(new_n139), .o1(new_n146));
  norp02aa1n09x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  nona23aa1n03x5               g054(.a(new_n142), .b(new_n148), .c(new_n147), .d(new_n139), .out0(new_n150));
  aoai13aa1n03x5               g055(.a(new_n150), .b(new_n149), .c(new_n146), .d(new_n142), .o1(\s[12] ));
  nano23aa1n03x7               g056(.a(new_n139), .b(new_n147), .c(new_n148), .d(new_n140), .out0(new_n152));
  nand02aa1n04x5               g057(.a(new_n152), .b(new_n136), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(new_n126), .b(new_n154), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n97), .b(new_n99), .c(new_n100), .o1(new_n156));
  nanb02aa1n02x5               g061(.a(new_n102), .b(new_n103), .out0(new_n157));
  inv000aa1d42x5               g062(.a(\a[3] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(\b[2] ), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(new_n159), .b(new_n158), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(new_n160), .b(new_n106), .o1(new_n161));
  nor003aa1n02x5               g066(.a(new_n156), .b(new_n157), .c(new_n161), .o1(new_n162));
  inv000aa1n02x5               g067(.a(new_n109), .o1(new_n163));
  nona23aa1n03x5               g068(.a(new_n119), .b(new_n117), .c(new_n116), .d(new_n118), .out0(new_n164));
  nano22aa1n03x7               g069(.a(new_n164), .b(new_n112), .c(new_n115), .out0(new_n165));
  tech160nm_fioai012aa1n05x5   g070(.a(new_n165), .b(new_n162), .c(new_n163), .o1(new_n166));
  tech160nm_fiaoi012aa1n03p5x5 g071(.a(new_n147), .b(new_n139), .c(new_n148), .o1(new_n167));
  aobi12aa1n06x5               g072(.a(new_n167), .b(new_n152), .c(new_n138), .out0(new_n168));
  aoai13aa1n04x5               g073(.a(new_n168), .b(new_n153), .c(new_n166), .d(new_n125), .o1(new_n169));
  xnrc02aa1n12x5               g074(.a(\b[12] ), .b(\a[13] ), .out0(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  nanb03aa1n02x5               g076(.a(new_n147), .b(new_n148), .c(new_n139), .out0(new_n172));
  oai112aa1n02x5               g077(.a(new_n172), .b(new_n170), .c(\b[11] ), .d(\a[12] ), .o1(new_n173));
  aoi012aa1n02x5               g078(.a(new_n173), .b(new_n138), .c(new_n152), .o1(new_n174));
  aoi022aa1n02x5               g079(.a(new_n169), .b(new_n171), .c(new_n155), .d(new_n174), .o1(\s[13] ));
  nor042aa1d18x5               g080(.a(\b[12] ), .b(\a[13] ), .o1(new_n176));
  inv040aa1d32x5               g081(.a(\a[14] ), .o1(new_n177));
  inv040aa1d32x5               g082(.a(\b[13] ), .o1(new_n178));
  nand22aa1n12x5               g083(.a(new_n178), .b(new_n177), .o1(new_n179));
  nand02aa1n02x5               g084(.a(\b[13] ), .b(\a[14] ), .o1(new_n180));
  nanp02aa1n03x5               g085(.a(new_n179), .b(new_n180), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n176), .c(new_n169), .d(new_n171), .o1(new_n182));
  oai112aa1n02x5               g087(.a(new_n179), .b(new_n180), .c(\b[12] ), .d(\a[13] ), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n171), .d(new_n169), .o1(\s[14] ));
  nona23aa1n09x5               g089(.a(new_n148), .b(new_n140), .c(new_n139), .d(new_n147), .out0(new_n185));
  oai012aa1n02x7               g090(.a(new_n167), .b(new_n185), .c(new_n137), .o1(new_n186));
  nor042aa1n06x5               g091(.a(new_n170), .b(new_n181), .o1(new_n187));
  aoai13aa1n06x5               g092(.a(new_n187), .b(new_n186), .c(new_n126), .d(new_n154), .o1(new_n188));
  oaoi03aa1n12x5               g093(.a(new_n177), .b(new_n178), .c(new_n176), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  norp02aa1n24x5               g095(.a(\b[14] ), .b(\a[15] ), .o1(new_n191));
  nand22aa1n04x5               g096(.a(\b[14] ), .b(\a[15] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  aoai13aa1n03x5               g099(.a(new_n194), .b(new_n190), .c(new_n169), .d(new_n187), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n179), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n191), .o1(new_n197));
  aoi122aa1n02x5               g102(.a(new_n196), .b(new_n176), .c(new_n180), .d(new_n197), .e(new_n192), .o1(new_n198));
  aobi12aa1n02x5               g103(.a(new_n195), .b(new_n198), .c(new_n188), .out0(\s[15] ));
  nor022aa1n06x5               g104(.a(\b[15] ), .b(\a[16] ), .o1(new_n200));
  nand22aa1n04x5               g105(.a(\b[15] ), .b(\a[16] ), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  norb03aa1n02x5               g107(.a(new_n201), .b(new_n191), .c(new_n200), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n193), .c(new_n188), .d(new_n189), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n204), .b(new_n202), .c(new_n195), .d(new_n197), .o1(\s[16] ));
  nona23aa1d18x5               g110(.a(new_n201), .b(new_n192), .c(new_n191), .d(new_n200), .out0(new_n206));
  nona23aa1d18x5               g111(.a(new_n187), .b(new_n136), .c(new_n206), .d(new_n185), .out0(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(new_n126), .b(new_n208), .o1(new_n209));
  nor003aa1n02x5               g114(.a(new_n206), .b(new_n181), .c(new_n170), .o1(new_n210));
  aoi012aa1n02x5               g115(.a(new_n200), .b(new_n191), .c(new_n201), .o1(new_n211));
  oaih12aa1n02x5               g116(.a(new_n211), .b(new_n206), .c(new_n189), .o1(new_n212));
  aoi012aa1n06x5               g117(.a(new_n212), .b(new_n186), .c(new_n210), .o1(new_n213));
  aoai13aa1n12x5               g118(.a(new_n213), .b(new_n207), .c(new_n166), .d(new_n125), .o1(new_n214));
  tech160nm_fixorc02aa1n03p5x5 g119(.a(\a[17] ), .b(\b[16] ), .out0(new_n215));
  aoi112aa1n02x5               g120(.a(new_n215), .b(new_n200), .c(new_n201), .d(new_n191), .o1(new_n216));
  oai012aa1n02x5               g121(.a(new_n216), .b(new_n206), .c(new_n189), .o1(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(new_n186), .c(new_n210), .o1(new_n218));
  aoi022aa1n02x5               g123(.a(new_n214), .b(new_n215), .c(new_n209), .d(new_n218), .o1(\s[17] ));
  nor042aa1n12x5               g124(.a(\b[16] ), .b(\a[17] ), .o1(new_n220));
  aoi012aa1n02x5               g125(.a(new_n220), .b(new_n214), .c(new_n215), .o1(new_n221));
  nor002aa1n10x5               g126(.a(\b[17] ), .b(\a[18] ), .o1(new_n222));
  nand02aa1d24x5               g127(.a(\b[17] ), .b(\a[18] ), .o1(new_n223));
  norb02aa1n02x7               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  norb03aa1n02x5               g129(.a(new_n223), .b(new_n220), .c(new_n222), .out0(new_n225));
  aob012aa1n02x5               g130(.a(new_n225), .b(new_n214), .c(new_n215), .out0(new_n226));
  oai012aa1n02x5               g131(.a(new_n226), .b(new_n221), .c(new_n224), .o1(\s[18] ));
  nanb02aa1n09x5               g132(.a(new_n206), .b(new_n187), .out0(new_n228));
  oabi12aa1n18x5               g133(.a(new_n212), .b(new_n168), .c(new_n228), .out0(new_n229));
  and002aa1n06x5               g134(.a(new_n215), .b(new_n224), .o(new_n230));
  aoai13aa1n03x5               g135(.a(new_n230), .b(new_n229), .c(new_n126), .d(new_n208), .o1(new_n231));
  aoi012aa1d24x5               g136(.a(new_n222), .b(new_n220), .c(new_n223), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  xorc02aa1n12x5               g138(.a(\a[19] ), .b(\b[18] ), .out0(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n233), .c(new_n214), .d(new_n230), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n234), .b(new_n222), .c(new_n223), .d(new_n220), .o1(new_n236));
  aobi12aa1n02x7               g141(.a(new_n235), .b(new_n236), .c(new_n231), .out0(\s[19] ));
  xnrc02aa1n02x5               g142(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g143(.a(\b[18] ), .b(\a[19] ), .o1(new_n239));
  inv000aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  nor042aa1n04x5               g145(.a(\b[19] ), .b(\a[20] ), .o1(new_n241));
  and002aa1n06x5               g146(.a(\b[19] ), .b(\a[20] ), .o(new_n242));
  nor042aa1n02x5               g147(.a(new_n242), .b(new_n241), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[18] ), .b(\a[19] ), .out0(new_n244));
  norp03aa1n02x5               g149(.a(new_n242), .b(new_n241), .c(new_n239), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n245), .b(new_n244), .c(new_n231), .d(new_n232), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n243), .c(new_n235), .d(new_n240), .o1(\s[20] ));
  nano32aa1n02x4               g152(.a(new_n244), .b(new_n215), .c(new_n243), .d(new_n224), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n229), .c(new_n126), .d(new_n208), .o1(new_n249));
  xnrc02aa1n12x5               g154(.a(\b[19] ), .b(\a[20] ), .out0(new_n250));
  oab012aa1d15x5               g155(.a(new_n241), .b(new_n240), .c(new_n242), .out0(new_n251));
  oai013aa1d12x5               g156(.a(new_n251), .b(new_n244), .c(new_n250), .d(new_n232), .o1(new_n252));
  nor042aa1d18x5               g157(.a(\b[20] ), .b(\a[21] ), .o1(new_n253));
  nanp02aa1n24x5               g158(.a(\b[20] ), .b(\a[21] ), .o1(new_n254));
  nanb02aa1n02x5               g159(.a(new_n253), .b(new_n254), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n03x5               g161(.a(new_n256), .b(new_n252), .c(new_n214), .d(new_n248), .o1(new_n257));
  nanb03aa1n06x5               g162(.a(new_n232), .b(new_n234), .c(new_n243), .out0(new_n258));
  nona22aa1n02x4               g163(.a(new_n239), .b(new_n242), .c(new_n241), .out0(new_n259));
  nano32aa1n02x4               g164(.a(new_n241), .b(new_n255), .c(new_n258), .d(new_n259), .out0(new_n260));
  aobi12aa1n02x7               g165(.a(new_n257), .b(new_n260), .c(new_n249), .out0(\s[21] ));
  inv000aa1d42x5               g166(.a(new_n253), .o1(new_n262));
  nor042aa1n06x5               g167(.a(\b[21] ), .b(\a[22] ), .o1(new_n263));
  nand42aa1d28x5               g168(.a(\b[21] ), .b(\a[22] ), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n264), .b(new_n263), .out0(new_n265));
  inv000aa1d42x5               g170(.a(new_n252), .o1(new_n266));
  norb03aa1n02x5               g171(.a(new_n264), .b(new_n253), .c(new_n263), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n255), .c(new_n249), .d(new_n266), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n265), .c(new_n257), .d(new_n262), .o1(\s[22] ));
  norp02aa1n02x5               g174(.a(new_n250), .b(new_n244), .o1(new_n270));
  nona23aa1n02x4               g175(.a(new_n264), .b(new_n254), .c(new_n253), .d(new_n263), .out0(new_n271));
  nano32aa1n02x4               g176(.a(new_n271), .b(new_n270), .c(new_n224), .d(new_n215), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n229), .c(new_n126), .d(new_n208), .o1(new_n273));
  nano23aa1n06x5               g178(.a(new_n253), .b(new_n263), .c(new_n264), .d(new_n254), .out0(new_n274));
  tech160nm_fiaoi012aa1n05x5   g179(.a(new_n263), .b(new_n253), .c(new_n264), .o1(new_n275));
  inv020aa1n03x5               g180(.a(new_n275), .o1(new_n276));
  aoi012aa1n12x5               g181(.a(new_n276), .b(new_n252), .c(new_n274), .o1(new_n277));
  inv000aa1n02x5               g182(.a(new_n277), .o1(new_n278));
  xorc02aa1n12x5               g183(.a(\a[23] ), .b(\b[22] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n278), .c(new_n214), .d(new_n272), .o1(new_n280));
  aoi112aa1n02x5               g185(.a(new_n279), .b(new_n263), .c(new_n264), .d(new_n253), .o1(new_n281));
  aobi12aa1n02x5               g186(.a(new_n281), .b(new_n252), .c(new_n274), .out0(new_n282));
  aobi12aa1n02x7               g187(.a(new_n280), .b(new_n282), .c(new_n273), .out0(\s[23] ));
  nor002aa1n06x5               g188(.a(\b[22] ), .b(\a[23] ), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[24] ), .b(\b[23] ), .out0(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[22] ), .b(\a[23] ), .out0(new_n287));
  orn002aa1n02x7               g192(.a(\a[24] ), .b(\b[23] ), .o(new_n288));
  nanp02aa1n02x5               g193(.a(\b[23] ), .b(\a[24] ), .o1(new_n289));
  nano22aa1n02x4               g194(.a(new_n284), .b(new_n288), .c(new_n289), .out0(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n287), .c(new_n273), .d(new_n277), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n286), .c(new_n280), .d(new_n285), .o1(\s[24] ));
  nand23aa1n02x5               g197(.a(new_n274), .b(new_n279), .c(new_n286), .o1(new_n293));
  nano32aa1n02x4               g198(.a(new_n293), .b(new_n270), .c(new_n224), .d(new_n215), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n229), .c(new_n126), .d(new_n208), .o1(new_n295));
  aob012aa1n06x5               g200(.a(new_n288), .b(new_n284), .c(new_n289), .out0(new_n296));
  aoi013aa1n06x4               g201(.a(new_n296), .b(new_n276), .c(new_n279), .d(new_n286), .o1(new_n297));
  aoai13aa1n12x5               g202(.a(new_n297), .b(new_n293), .c(new_n258), .d(new_n251), .o1(new_n298));
  xorc02aa1n12x5               g203(.a(\a[25] ), .b(\b[24] ), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n298), .c(new_n214), .d(new_n294), .o1(new_n300));
  norb03aa1n02x5               g205(.a(new_n286), .b(new_n271), .c(new_n287), .out0(new_n301));
  norb03aa1n02x5               g206(.a(new_n286), .b(new_n275), .c(new_n287), .out0(new_n302));
  nanp03aa1n02x5               g207(.a(new_n288), .b(new_n284), .c(new_n289), .o1(new_n303));
  nanb03aa1n02x5               g208(.a(new_n299), .b(new_n288), .c(new_n303), .out0(new_n304));
  aoi112aa1n02x5               g209(.a(new_n304), .b(new_n302), .c(new_n252), .d(new_n301), .o1(new_n305));
  aobi12aa1n02x7               g210(.a(new_n300), .b(new_n305), .c(new_n295), .out0(\s[25] ));
  nor042aa1n03x5               g211(.a(\b[24] ), .b(\a[25] ), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  norp02aa1n12x5               g213(.a(\b[25] ), .b(\a[26] ), .o1(new_n309));
  and002aa1n12x5               g214(.a(\b[25] ), .b(\a[26] ), .o(new_n310));
  norp02aa1n06x5               g215(.a(new_n310), .b(new_n309), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n298), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n299), .o1(new_n313));
  norp03aa1n02x5               g218(.a(new_n310), .b(new_n309), .c(new_n307), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n313), .c(new_n295), .d(new_n312), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n300), .d(new_n308), .o1(\s[26] ));
  and002aa1n12x5               g221(.a(new_n299), .b(new_n311), .o(new_n317));
  nano32aa1n03x7               g222(.a(new_n293), .b(new_n317), .c(new_n230), .d(new_n270), .out0(new_n318));
  aoai13aa1n09x5               g223(.a(new_n318), .b(new_n229), .c(new_n126), .d(new_n208), .o1(new_n319));
  nanp02aa1n03x5               g224(.a(new_n252), .b(new_n301), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n317), .o1(new_n321));
  oab012aa1n02x4               g226(.a(new_n309), .b(new_n308), .c(new_n310), .out0(new_n322));
  aoai13aa1n04x5               g227(.a(new_n322), .b(new_n321), .c(new_n320), .d(new_n297), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[27] ), .b(\b[26] ), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n323), .c(new_n214), .d(new_n318), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n309), .o1(new_n326));
  inv000aa1n02x5               g231(.a(new_n324), .o1(new_n327));
  oai112aa1n02x5               g232(.a(new_n327), .b(new_n326), .c(new_n310), .d(new_n308), .o1(new_n328));
  aoi012aa1n02x5               g233(.a(new_n328), .b(new_n298), .c(new_n317), .o1(new_n329));
  aobi12aa1n02x7               g234(.a(new_n325), .b(new_n329), .c(new_n319), .out0(\s[27] ));
  nor042aa1n03x5               g235(.a(\b[26] ), .b(\a[27] ), .o1(new_n331));
  inv020aa1n02x5               g236(.a(new_n331), .o1(new_n332));
  nor042aa1n03x5               g237(.a(\b[27] ), .b(\a[28] ), .o1(new_n333));
  and002aa1n12x5               g238(.a(\b[27] ), .b(\a[28] ), .o(new_n334));
  norp02aa1n02x5               g239(.a(new_n334), .b(new_n333), .o1(new_n335));
  aobi12aa1n06x5               g240(.a(new_n322), .b(new_n298), .c(new_n317), .out0(new_n336));
  norp03aa1n02x5               g241(.a(new_n334), .b(new_n333), .c(new_n331), .o1(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n327), .c(new_n319), .d(new_n336), .o1(new_n338));
  aoai13aa1n03x5               g243(.a(new_n338), .b(new_n335), .c(new_n325), .d(new_n332), .o1(\s[28] ));
  inv000aa1d42x5               g244(.a(\a[28] ), .o1(new_n340));
  inv000aa1d42x5               g245(.a(\b[26] ), .o1(new_n341));
  xroi22aa1d04x5               g246(.a(\a[27] ), .b(new_n341), .c(new_n340), .d(\b[27] ), .out0(new_n342));
  aoai13aa1n02x5               g247(.a(new_n342), .b(new_n323), .c(new_n214), .d(new_n318), .o1(new_n343));
  oab012aa1n06x5               g248(.a(new_n333), .b(new_n332), .c(new_n334), .out0(new_n344));
  norp02aa1n02x5               g249(.a(\b[28] ), .b(\a[29] ), .o1(new_n345));
  nand42aa1n03x5               g250(.a(\b[28] ), .b(\a[29] ), .o1(new_n346));
  norb02aa1n02x5               g251(.a(new_n346), .b(new_n345), .out0(new_n347));
  inv000aa1d42x5               g252(.a(new_n342), .o1(new_n348));
  nona22aa1n02x4               g253(.a(new_n331), .b(new_n334), .c(new_n333), .out0(new_n349));
  nano23aa1n02x4               g254(.a(new_n333), .b(new_n345), .c(new_n349), .d(new_n346), .out0(new_n350));
  aoai13aa1n03x5               g255(.a(new_n350), .b(new_n348), .c(new_n319), .d(new_n336), .o1(new_n351));
  aoai13aa1n03x5               g256(.a(new_n351), .b(new_n347), .c(new_n343), .d(new_n344), .o1(\s[29] ));
  xorb03aa1n02x5               g257(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g258(.a(new_n327), .b(new_n335), .c(new_n347), .out0(new_n354));
  aoai13aa1n03x5               g259(.a(new_n354), .b(new_n323), .c(new_n214), .d(new_n318), .o1(new_n355));
  tech160nm_fioaoi03aa1n03p5x5 g260(.a(\a[29] ), .b(\b[28] ), .c(new_n344), .o1(new_n356));
  inv000aa1d42x5               g261(.a(new_n356), .o1(new_n357));
  norp02aa1n02x5               g262(.a(\b[29] ), .b(\a[30] ), .o1(new_n358));
  nanp02aa1n02x5               g263(.a(\b[29] ), .b(\a[30] ), .o1(new_n359));
  norb02aa1n02x5               g264(.a(new_n359), .b(new_n358), .out0(new_n360));
  inv000aa1d42x5               g265(.a(new_n354), .o1(new_n361));
  nanb02aa1n02x5               g266(.a(new_n344), .b(new_n347), .out0(new_n362));
  nano23aa1n02x4               g267(.a(new_n345), .b(new_n358), .c(new_n362), .d(new_n359), .out0(new_n363));
  aoai13aa1n03x5               g268(.a(new_n363), .b(new_n361), .c(new_n319), .d(new_n336), .o1(new_n364));
  aoai13aa1n03x5               g269(.a(new_n364), .b(new_n360), .c(new_n355), .d(new_n357), .o1(\s[30] ));
  nano32aa1n03x7               g270(.a(new_n327), .b(new_n360), .c(new_n335), .d(new_n347), .out0(new_n366));
  aoai13aa1n03x5               g271(.a(new_n366), .b(new_n323), .c(new_n214), .d(new_n318), .o1(new_n367));
  aoi012aa1n02x5               g272(.a(new_n358), .b(new_n356), .c(new_n359), .o1(new_n368));
  xnrc02aa1n02x5               g273(.a(\b[30] ), .b(\a[31] ), .out0(new_n369));
  inv000aa1d42x5               g274(.a(new_n369), .o1(new_n370));
  inv000aa1d42x5               g275(.a(new_n366), .o1(new_n371));
  aoi112aa1n02x5               g276(.a(new_n358), .b(new_n369), .c(new_n356), .d(new_n360), .o1(new_n372));
  aoai13aa1n03x5               g277(.a(new_n372), .b(new_n371), .c(new_n319), .d(new_n336), .o1(new_n373));
  aoai13aa1n03x5               g278(.a(new_n373), .b(new_n370), .c(new_n367), .d(new_n368), .o1(\s[31] ));
  aoi112aa1n02x5               g279(.a(new_n107), .b(new_n97), .c(new_n99), .d(new_n100), .o1(new_n375));
  aoi012aa1n02x5               g280(.a(new_n375), .b(new_n101), .c(new_n107), .o1(\s[3] ));
  aoai13aa1n02x5               g281(.a(new_n107), .b(new_n97), .c(new_n100), .d(new_n99), .o1(new_n377));
  xnbna2aa1n03x5               g282(.a(new_n104), .b(new_n377), .c(new_n160), .out0(\s[4] ));
  oai013aa1n02x4               g283(.a(new_n109), .b(new_n156), .c(new_n157), .d(new_n161), .o1(new_n379));
  aoi112aa1n02x5               g284(.a(new_n112), .b(new_n102), .c(new_n103), .d(new_n105), .o1(new_n380));
  aoi022aa1n02x5               g285(.a(new_n379), .b(new_n112), .c(new_n108), .d(new_n380), .o1(\s[5] ));
  oai012aa1n02x5               g286(.a(new_n112), .b(new_n162), .c(new_n163), .o1(new_n382));
  nona23aa1n02x4               g287(.a(new_n382), .b(new_n114), .c(new_n110), .d(new_n113), .out0(new_n383));
  aoai13aa1n02x5               g288(.a(new_n383), .b(new_n115), .c(new_n122), .d(new_n382), .o1(\s[6] ));
  nanp03aa1n02x5               g289(.a(new_n379), .b(new_n112), .c(new_n115), .o1(new_n385));
  norb02aa1n02x5               g290(.a(new_n119), .b(new_n118), .out0(new_n386));
  inv000aa1d42x5               g291(.a(new_n123), .o1(new_n387));
  aobi12aa1n02x5               g292(.a(new_n386), .b(new_n385), .c(new_n387), .out0(new_n388));
  aoi112aa1n02x5               g293(.a(new_n386), .b(new_n113), .c(new_n114), .d(new_n110), .o1(new_n389));
  aoi012aa1n02x5               g294(.a(new_n388), .b(new_n385), .c(new_n389), .o1(\s[7] ));
  obai22aa1n02x7               g295(.a(new_n117), .b(new_n116), .c(new_n388), .d(new_n118), .out0(new_n391));
  norb03aa1n02x5               g296(.a(new_n117), .b(new_n116), .c(new_n118), .out0(new_n392));
  oaib12aa1n02x5               g297(.a(new_n391), .b(new_n388), .c(new_n392), .out0(\s[8] ));
  aoi112aa1n02x5               g298(.a(new_n129), .b(new_n116), .c(new_n117), .d(new_n118), .o1(new_n394));
  aobi12aa1n02x5               g299(.a(new_n394), .b(new_n123), .c(new_n120), .out0(new_n395));
  aoi022aa1n02x5               g300(.a(new_n126), .b(new_n129), .c(new_n166), .d(new_n395), .o1(\s[9] ));
endmodule


