// Benchmark "adder" written by ABC on Wed Jul 17 19:05:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n336, new_n339, new_n340,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n348;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  oai022aa1n02x7               g003(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n99));
  tech160nm_fixorc02aa1n04x5   g004(.a(\a[7] ), .b(\b[6] ), .out0(new_n100));
  aoi022aa1d24x5               g005(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n101));
  orn002aa1n24x5               g006(.a(\a[7] ), .b(\b[6] ), .o(new_n102));
  oaoi03aa1n12x5               g007(.a(\a[8] ), .b(\b[7] ), .c(new_n102), .o1(new_n103));
  aoi013aa1n06x4               g008(.a(new_n103), .b(new_n100), .c(new_n101), .d(new_n99), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  and002aa1n02x5               g010(.a(\b[4] ), .b(\a[5] ), .o(new_n106));
  nano32aa1n03x7               g011(.a(new_n106), .b(new_n101), .c(new_n102), .d(new_n105), .out0(new_n107));
  and002aa1n03x5               g012(.a(\b[0] ), .b(\a[1] ), .o(new_n108));
  oaoi03aa1n03x5               g013(.a(\a[2] ), .b(\b[1] ), .c(new_n108), .o1(new_n109));
  nor022aa1n16x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nand02aa1n08x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nor002aa1n03x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nand02aa1n03x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nano23aa1n06x5               g018(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n114));
  inv000aa1d42x5               g019(.a(\a[3] ), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\b[2] ), .o1(new_n116));
  aoai13aa1n06x5               g021(.a(new_n111), .b(new_n110), .c(new_n115), .d(new_n116), .o1(new_n117));
  inv040aa1n03x5               g022(.a(new_n117), .o1(new_n118));
  aoai13aa1n06x5               g023(.a(new_n107), .b(new_n118), .c(new_n114), .d(new_n109), .o1(new_n119));
  nanp02aa1n09x5               g024(.a(new_n119), .b(new_n104), .o1(new_n120));
  oaoi03aa1n09x5               g025(.a(new_n97), .b(new_n98), .c(new_n120), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\a[10] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[9] ), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n123), .b(new_n122), .o1(new_n124));
  nand42aa1n16x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n121), .b(new_n125), .c(new_n124), .out0(\s[10] ));
  nanp02aa1n09x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nor002aa1d32x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  norb02aa1n12x5               g033(.a(new_n127), .b(new_n128), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  nanp02aa1n03x5               g035(.a(new_n121), .b(new_n124), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n130), .b(new_n131), .c(new_n125), .out0(\s[11] ));
  inv000aa1d42x5               g037(.a(new_n128), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n125), .o1(new_n134));
  nona22aa1n02x4               g039(.a(new_n131), .b(new_n130), .c(new_n134), .out0(new_n135));
  nor002aa1n02x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand22aa1n12x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aobi12aa1n06x5               g043(.a(new_n138), .b(new_n135), .c(new_n133), .out0(new_n139));
  aoi112aa1n03x5               g044(.a(new_n130), .b(new_n134), .c(new_n121), .d(new_n124), .o1(new_n140));
  norp03aa1n02x5               g045(.a(new_n140), .b(new_n138), .c(new_n128), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n139), .b(new_n141), .o1(\s[12] ));
  inv040aa1n02x5               g047(.a(new_n137), .o1(new_n143));
  oai022aa1d18x5               g048(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n144));
  inv000aa1n04x5               g049(.a(new_n144), .o1(new_n145));
  nanb03aa1d24x5               g050(.a(new_n128), .b(new_n125), .c(new_n127), .out0(new_n146));
  tech160nm_fioai012aa1n04x5   g051(.a(new_n137), .b(new_n136), .c(new_n128), .o1(new_n147));
  oai013aa1d12x5               g052(.a(new_n147), .b(new_n146), .c(new_n143), .d(new_n145), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nanp03aa1n02x5               g054(.a(new_n101), .b(new_n102), .c(new_n105), .o1(new_n150));
  inv000aa1n02x5               g055(.a(new_n103), .o1(new_n151));
  oaib12aa1n02x5               g056(.a(new_n151), .b(new_n150), .c(new_n99), .out0(new_n152));
  inv000aa1d42x5               g057(.a(\a[1] ), .o1(new_n153));
  inv000aa1d42x5               g058(.a(\b[0] ), .o1(new_n154));
  norp02aa1n02x5               g059(.a(\b[1] ), .b(\a[2] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(\b[1] ), .b(\a[2] ), .o1(new_n156));
  oaoi13aa1n09x5               g061(.a(new_n155), .b(new_n156), .c(new_n153), .d(new_n154), .o1(new_n157));
  nona23aa1n09x5               g062(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n158));
  oai012aa1n18x5               g063(.a(new_n117), .b(new_n158), .c(new_n157), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(\b[8] ), .b(\a[9] ), .o1(new_n160));
  nano22aa1n03x7               g065(.a(new_n146), .b(new_n160), .c(new_n137), .out0(new_n161));
  aoai13aa1n06x5               g066(.a(new_n161), .b(new_n152), .c(new_n159), .d(new_n107), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(new_n162), .b(new_n149), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n03x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  tech160nm_finand02aa1n03p5x5 g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n165), .b(new_n163), .c(new_n166), .o1(new_n167));
  xnrb03aa1n02x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nona23aa1n09x5               g075(.a(new_n170), .b(new_n166), .c(new_n165), .d(new_n169), .out0(new_n171));
  aoi012aa1n02x5               g076(.a(new_n169), .b(new_n165), .c(new_n170), .o1(new_n172));
  aoai13aa1n04x5               g077(.a(new_n172), .b(new_n171), .c(new_n162), .d(new_n149), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv000aa1d42x5               g079(.a(\a[15] ), .o1(new_n175));
  nanb02aa1d36x5               g080(.a(\b[14] ), .b(new_n175), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  xnrc02aa1n12x5               g083(.a(\b[15] ), .b(\a[16] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n177), .b(new_n180), .c(new_n173), .d(new_n178), .o1(new_n181));
  aoai13aa1n03x5               g086(.a(new_n180), .b(new_n177), .c(new_n173), .d(new_n178), .o1(new_n182));
  norb02aa1n02x7               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  aoi012aa1n03x5               g088(.a(new_n152), .b(new_n159), .c(new_n107), .o1(new_n184));
  nona22aa1n03x5               g089(.a(new_n129), .b(new_n143), .c(new_n134), .out0(new_n185));
  nano32aa1n03x7               g090(.a(new_n185), .b(new_n147), .c(new_n145), .d(new_n160), .out0(new_n186));
  nand02aa1n03x5               g091(.a(new_n176), .b(new_n178), .o1(new_n187));
  nor043aa1n03x5               g092(.a(new_n171), .b(new_n187), .c(new_n179), .o1(new_n188));
  nand22aa1n03x5               g093(.a(new_n186), .b(new_n188), .o1(new_n189));
  norp02aa1n02x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  aoai13aa1n02x5               g095(.a(new_n178), .b(new_n169), .c(new_n165), .d(new_n170), .o1(new_n191));
  aoi022aa1n03x5               g096(.a(new_n191), .b(new_n176), .c(\a[16] ), .d(\b[15] ), .o1(new_n192));
  aoi112aa1n02x7               g097(.a(new_n190), .b(new_n192), .c(new_n148), .d(new_n188), .o1(new_n193));
  oai012aa1n06x5               g098(.a(new_n193), .b(new_n184), .c(new_n189), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  aoi012aa1n12x5               g100(.a(new_n189), .b(new_n119), .c(new_n104), .o1(new_n196));
  nano22aa1n03x7               g101(.a(new_n146), .b(new_n137), .c(new_n144), .out0(new_n197));
  oaib12aa1n06x5               g102(.a(new_n188), .b(new_n197), .c(new_n147), .out0(new_n198));
  nona22aa1n12x5               g103(.a(new_n198), .b(new_n192), .c(new_n190), .out0(new_n199));
  nor042aa1d18x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  nand42aa1n16x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  oaoi13aa1n03x5               g106(.a(new_n200), .b(new_n201), .c(new_n196), .d(new_n199), .o1(new_n202));
  xnrb03aa1n03x5               g107(.a(new_n202), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nano23aa1n02x5               g108(.a(new_n165), .b(new_n169), .c(new_n170), .d(new_n166), .out0(new_n204));
  norp02aa1n02x5               g109(.a(new_n179), .b(new_n187), .o1(new_n205));
  nano32aa1n03x7               g110(.a(new_n148), .b(new_n205), .c(new_n161), .d(new_n204), .out0(new_n206));
  nor042aa1n12x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nand02aa1d28x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nano23aa1n06x5               g113(.a(new_n200), .b(new_n207), .c(new_n208), .d(new_n201), .out0(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n199), .c(new_n120), .d(new_n206), .o1(new_n210));
  tech160nm_fiao0012aa1n02p5x5 g115(.a(new_n207), .b(new_n200), .c(new_n208), .o(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  orn002aa1n24x5               g117(.a(\a[19] ), .b(\b[18] ), .o(new_n213));
  nand42aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand02aa1d04x5               g119(.a(new_n213), .b(new_n214), .o1(new_n215));
  xobna2aa1n03x5               g120(.a(new_n215), .b(new_n210), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoi012aa1n06x5               g122(.a(new_n215), .b(new_n210), .c(new_n212), .o1(new_n218));
  xnrc02aa1n03x5               g123(.a(\b[19] ), .b(\a[20] ), .out0(new_n219));
  nano22aa1n03x7               g124(.a(new_n218), .b(new_n213), .c(new_n219), .out0(new_n220));
  oaoi13aa1n02x5               g125(.a(new_n211), .b(new_n209), .c(new_n196), .d(new_n199), .o1(new_n221));
  oaoi13aa1n02x5               g126(.a(new_n219), .b(new_n213), .c(new_n221), .d(new_n215), .o1(new_n222));
  norp02aa1n03x5               g127(.a(new_n222), .b(new_n220), .o1(\s[20] ));
  inv000aa1d42x5               g128(.a(\a[21] ), .o1(new_n224));
  nona22aa1d18x5               g129(.a(new_n209), .b(new_n219), .c(new_n215), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  orn002aa1n02x5               g131(.a(\a[20] ), .b(\b[19] ), .o(new_n227));
  and002aa1n02x5               g132(.a(\b[19] ), .b(\a[20] ), .o(new_n228));
  aoai13aa1n12x5               g133(.a(new_n214), .b(new_n207), .c(new_n200), .d(new_n208), .o1(new_n229));
  aoai13aa1n12x5               g134(.a(new_n227), .b(new_n228), .c(new_n229), .d(new_n213), .o1(new_n230));
  oaoi13aa1n06x5               g135(.a(new_n230), .b(new_n226), .c(new_n196), .d(new_n199), .o1(new_n231));
  xorb03aa1n03x5               g136(.a(new_n231), .b(\b[20] ), .c(new_n224), .out0(\s[21] ));
  nor042aa1d18x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoi012aa1n02x5               g139(.a(new_n199), .b(new_n120), .c(new_n206), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n230), .o1(new_n236));
  xorc02aa1n12x5               g141(.a(\a[21] ), .b(\b[20] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  oaoi13aa1n02x5               g143(.a(new_n238), .b(new_n236), .c(new_n235), .d(new_n225), .o1(new_n239));
  nor002aa1n12x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nand42aa1d28x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  norb02aa1d27x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  inv000aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  nano22aa1n02x4               g148(.a(new_n239), .b(new_n234), .c(new_n243), .out0(new_n244));
  oaoi13aa1n03x5               g149(.a(new_n243), .b(new_n234), .c(new_n231), .d(new_n238), .o1(new_n245));
  norp02aa1n02x5               g150(.a(new_n245), .b(new_n244), .o1(\s[22] ));
  nand22aa1n12x5               g151(.a(new_n237), .b(new_n242), .o1(new_n247));
  nor042aa1n02x5               g152(.a(new_n225), .b(new_n247), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n247), .o1(new_n249));
  aoi012aa1n02x5               g154(.a(new_n240), .b(new_n233), .c(new_n241), .o1(new_n250));
  aob012aa1n06x5               g155(.a(new_n250), .b(new_n230), .c(new_n249), .out0(new_n251));
  oaoi13aa1n09x5               g156(.a(new_n251), .b(new_n248), .c(new_n196), .d(new_n199), .o1(new_n252));
  orn002aa1n24x5               g157(.a(\a[23] ), .b(\b[22] ), .o(new_n253));
  nand02aa1n06x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n252), .b(new_n254), .c(new_n253), .out0(\s[23] ));
  aoai13aa1n02x5               g160(.a(new_n248), .b(new_n199), .c(new_n120), .d(new_n206), .o1(new_n256));
  nanp02aa1n02x5               g161(.a(new_n253), .b(new_n254), .o1(new_n257));
  aoib12aa1n02x7               g162(.a(new_n257), .b(new_n256), .c(new_n251), .out0(new_n258));
  xorc02aa1n12x5               g163(.a(\a[24] ), .b(\b[23] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  nano22aa1n03x5               g165(.a(new_n258), .b(new_n253), .c(new_n260), .out0(new_n261));
  oaoi13aa1n03x5               g166(.a(new_n260), .b(new_n253), .c(new_n252), .d(new_n257), .o1(new_n262));
  norp02aa1n03x5               g167(.a(new_n262), .b(new_n261), .o1(\s[24] ));
  nona23aa1n06x5               g168(.a(new_n259), .b(new_n237), .c(new_n243), .d(new_n257), .out0(new_n264));
  nor042aa1n02x5               g169(.a(new_n264), .b(new_n225), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n199), .c(new_n120), .d(new_n206), .o1(new_n266));
  nano32aa1d12x5               g171(.a(new_n247), .b(new_n259), .c(new_n253), .d(new_n254), .out0(new_n267));
  nanp02aa1n12x5               g172(.a(new_n267), .b(new_n230), .o1(new_n268));
  inv000aa1d42x5               g173(.a(\a[24] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(\b[23] ), .o1(new_n270));
  nanp02aa1n02x5               g175(.a(new_n270), .b(new_n269), .o1(new_n271));
  and002aa1n02x5               g176(.a(\b[23] ), .b(\a[24] ), .o(new_n272));
  aoai13aa1n02x5               g177(.a(new_n254), .b(new_n240), .c(new_n233), .d(new_n241), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n271), .b(new_n272), .c(new_n273), .d(new_n253), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nand22aa1n12x5               g180(.a(new_n268), .b(new_n275), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  xnrc02aa1n12x5               g182(.a(\b[24] ), .b(\a[25] ), .out0(new_n278));
  xobna2aa1n03x5               g183(.a(new_n278), .b(new_n266), .c(new_n277), .out0(\s[25] ));
  inv000aa1d42x5               g184(.a(\a[25] ), .o1(new_n280));
  nanb02aa1n02x5               g185(.a(\b[24] ), .b(new_n280), .out0(new_n281));
  tech160nm_fiaoi012aa1n02p5x5 g186(.a(new_n278), .b(new_n266), .c(new_n277), .o1(new_n282));
  xnrc02aa1n06x5               g187(.a(\b[25] ), .b(\a[26] ), .out0(new_n283));
  nano22aa1n03x7               g188(.a(new_n282), .b(new_n281), .c(new_n283), .out0(new_n284));
  oaoi13aa1n04x5               g189(.a(new_n276), .b(new_n265), .c(new_n196), .d(new_n199), .o1(new_n285));
  oaoi13aa1n03x5               g190(.a(new_n283), .b(new_n281), .c(new_n285), .d(new_n278), .o1(new_n286));
  norp02aa1n03x5               g191(.a(new_n286), .b(new_n284), .o1(\s[26] ));
  nor042aa1n02x5               g192(.a(new_n283), .b(new_n278), .o1(new_n288));
  norb03aa1n06x5               g193(.a(new_n288), .b(new_n264), .c(new_n225), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n199), .c(new_n120), .d(new_n206), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n281), .carry(new_n291));
  aobi12aa1n18x5               g196(.a(new_n291), .b(new_n276), .c(new_n288), .out0(new_n292));
  xorc02aa1n12x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  xnbna2aa1n03x5               g198(.a(new_n293), .b(new_n292), .c(new_n290), .out0(\s[27] ));
  norp02aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  inv040aa1n03x5               g200(.a(new_n295), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n293), .o1(new_n297));
  tech160nm_fiaoi012aa1n05x5   g202(.a(new_n297), .b(new_n292), .c(new_n290), .o1(new_n298));
  tech160nm_fixnrc02aa1n04x5   g203(.a(\b[27] ), .b(\a[28] ), .out0(new_n299));
  nano22aa1n03x7               g204(.a(new_n298), .b(new_n296), .c(new_n299), .out0(new_n300));
  aoai13aa1n06x5               g205(.a(new_n288), .b(new_n274), .c(new_n267), .d(new_n230), .o1(new_n301));
  nand22aa1n03x5               g206(.a(new_n301), .b(new_n291), .o1(new_n302));
  aoai13aa1n02x5               g207(.a(new_n293), .b(new_n302), .c(new_n194), .d(new_n289), .o1(new_n303));
  aoi012aa1n02x5               g208(.a(new_n299), .b(new_n303), .c(new_n296), .o1(new_n304));
  norp02aa1n03x5               g209(.a(new_n304), .b(new_n300), .o1(\s[28] ));
  norb02aa1n06x5               g210(.a(new_n293), .b(new_n299), .out0(new_n306));
  aoai13aa1n02x5               g211(.a(new_n306), .b(new_n302), .c(new_n194), .d(new_n289), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n296), .carry(new_n308));
  xnrc02aa1n12x5               g213(.a(\b[28] ), .b(\a[29] ), .out0(new_n309));
  aoi012aa1n03x5               g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n306), .o1(new_n311));
  tech160nm_fiaoi012aa1n05x5   g216(.a(new_n311), .b(new_n292), .c(new_n290), .o1(new_n312));
  nano22aa1n03x7               g217(.a(new_n312), .b(new_n308), .c(new_n309), .out0(new_n313));
  nor002aa1n02x5               g218(.a(new_n310), .b(new_n313), .o1(\s[29] ));
  xnrb03aa1n02x5               g219(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1d15x5               g220(.a(new_n293), .b(new_n309), .c(new_n299), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n302), .c(new_n194), .d(new_n289), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .carry(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .out0(new_n319));
  aoi012aa1n02x5               g224(.a(new_n319), .b(new_n317), .c(new_n318), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n316), .o1(new_n321));
  tech160nm_fiaoi012aa1n05x5   g226(.a(new_n321), .b(new_n292), .c(new_n290), .o1(new_n322));
  nano22aa1n03x7               g227(.a(new_n322), .b(new_n318), .c(new_n319), .out0(new_n323));
  norp02aa1n03x5               g228(.a(new_n320), .b(new_n323), .o1(\s[30] ));
  norb02aa1n06x5               g229(.a(new_n316), .b(new_n319), .out0(new_n325));
  aoai13aa1n02x5               g230(.a(new_n325), .b(new_n302), .c(new_n194), .d(new_n289), .o1(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n318), .carry(new_n327));
  xnrc02aa1n02x5               g232(.a(\b[30] ), .b(\a[31] ), .out0(new_n328));
  aoi012aa1n03x5               g233(.a(new_n328), .b(new_n326), .c(new_n327), .o1(new_n329));
  inv000aa1d42x5               g234(.a(new_n325), .o1(new_n330));
  tech160nm_fiaoi012aa1n05x5   g235(.a(new_n330), .b(new_n292), .c(new_n290), .o1(new_n331));
  nano22aa1n03x7               g236(.a(new_n331), .b(new_n327), .c(new_n328), .out0(new_n332));
  nor002aa1n02x5               g237(.a(new_n329), .b(new_n332), .o1(\s[31] ));
  xorb03aa1n02x5               g238(.a(new_n157), .b(\b[2] ), .c(new_n115), .out0(\s[3] ));
  nanb03aa1n02x5               g239(.a(new_n112), .b(new_n109), .c(new_n113), .out0(new_n335));
  aboi22aa1n03x5               g240(.a(new_n110), .b(new_n111), .c(new_n115), .d(new_n116), .out0(new_n336));
  aboi22aa1n03x5               g241(.a(new_n110), .b(new_n159), .c(new_n335), .d(new_n336), .out0(\s[4] ));
  xorb03aa1n02x5               g242(.a(new_n159), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1n06x5               g243(.a(new_n159), .o1(new_n339));
  oaoi03aa1n09x5               g244(.a(\a[5] ), .b(\b[4] ), .c(new_n339), .o1(new_n340));
  xorb03aa1n02x5               g245(.a(new_n340), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  orn002aa1n02x5               g246(.a(\a[6] ), .b(\b[5] ), .o(new_n342));
  inv000aa1d42x5               g247(.a(new_n342), .o1(new_n343));
  nanp02aa1n02x5               g248(.a(\b[5] ), .b(\a[6] ), .o1(new_n344));
  aoi112aa1n02x5               g249(.a(new_n343), .b(new_n100), .c(new_n340), .d(new_n344), .o1(new_n345));
  aoai13aa1n06x5               g250(.a(new_n100), .b(new_n343), .c(new_n340), .d(new_n344), .o1(new_n346));
  norb02aa1n02x5               g251(.a(new_n346), .b(new_n345), .out0(\s[7] ));
  xorc02aa1n02x5               g252(.a(\a[8] ), .b(\b[7] ), .out0(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n348), .b(new_n346), .c(new_n102), .out0(\s[8] ));
  xorb03aa1n02x5               g254(.a(new_n120), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


