// Benchmark "adder" written by ABC on Wed Jul 17 15:21:24 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n341, new_n342, new_n343, new_n345,
    new_n346, new_n349, new_n350, new_n351, new_n352, new_n354, new_n355,
    new_n357;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  and002aa1n03x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n09x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano23aa1n06x5               g009(.a(new_n103), .b(new_n102), .c(new_n104), .d(new_n101), .out0(new_n105));
  nanp02aa1n03x5               g010(.a(new_n105), .b(new_n100), .o1(new_n106));
  aoi012aa1n02x5               g011(.a(new_n102), .b(new_n103), .c(new_n101), .o1(new_n107));
  nand02aa1d04x5               g012(.a(new_n106), .b(new_n107), .o1(new_n108));
  nand02aa1n08x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor002aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  norp02aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nano23aa1n06x5               g017(.a(new_n111), .b(new_n110), .c(new_n112), .d(new_n109), .out0(new_n113));
  xorc02aa1n12x5               g018(.a(\a[5] ), .b(\b[4] ), .out0(new_n114));
  nor042aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand02aa1d24x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  norb02aa1n03x4               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nand23aa1n04x5               g022(.a(new_n113), .b(new_n114), .c(new_n117), .o1(new_n118));
  inv000aa1n06x5               g023(.a(new_n118), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n109), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n110), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n111), .o1(new_n122));
  nor042aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  aoai13aa1n06x5               g028(.a(new_n112), .b(new_n115), .c(new_n123), .d(new_n116), .o1(new_n124));
  aoai13aa1n02x7               g029(.a(new_n121), .b(new_n120), .c(new_n124), .d(new_n122), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n125), .c(new_n119), .d(new_n108), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[10] ), .b(\b[9] ), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  aobi12aa1n06x5               g034(.a(new_n107), .b(new_n105), .c(new_n100), .out0(new_n130));
  nand02aa1n02x5               g035(.a(new_n124), .b(new_n122), .o1(new_n131));
  aoi012aa1n02x7               g036(.a(new_n110), .b(new_n131), .c(new_n109), .o1(new_n132));
  oai012aa1n12x5               g037(.a(new_n132), .b(new_n130), .c(new_n118), .o1(new_n133));
  aoai13aa1n06x5               g038(.a(new_n128), .b(new_n97), .c(new_n133), .d(new_n126), .o1(new_n134));
  norp02aa1n04x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  oai012aa1n12x5               g041(.a(new_n136), .b(new_n135), .c(new_n97), .o1(new_n137));
  nor002aa1d24x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nanp02aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n06x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n134), .c(new_n137), .out0(\s[11] ));
  nand02aa1n03x5               g046(.a(new_n127), .b(new_n98), .o1(new_n142));
  inv040aa1n02x5               g047(.a(new_n137), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n140), .b(new_n143), .c(new_n142), .d(new_n128), .o1(new_n144));
  nor022aa1n08x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand02aa1n06x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nanb02aa1n03x5               g051(.a(new_n145), .b(new_n146), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  aoib12aa1n02x5               g053(.a(new_n138), .b(new_n146), .c(new_n145), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n138), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n140), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n150), .b(new_n151), .c(new_n134), .d(new_n137), .o1(new_n152));
  aoi022aa1n03x5               g057(.a(new_n152), .b(new_n148), .c(new_n144), .d(new_n149), .o1(\s[12] ));
  nano23aa1n06x5               g058(.a(new_n138), .b(new_n145), .c(new_n146), .d(new_n139), .out0(new_n154));
  nand23aa1d12x5               g059(.a(new_n154), .b(new_n126), .c(new_n128), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  aoai13aa1n04x5               g061(.a(new_n156), .b(new_n125), .c(new_n119), .d(new_n108), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n145), .b(new_n138), .c(new_n146), .o1(new_n158));
  aobi12aa1n06x5               g063(.a(new_n158), .b(new_n154), .c(new_n143), .out0(new_n159));
  xnrc02aa1n12x5               g064(.a(\b[12] ), .b(\a[13] ), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n157), .c(new_n159), .out0(\s[13] ));
  nor042aa1n06x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  inv000aa1n02x5               g068(.a(new_n163), .o1(new_n164));
  oai013aa1n09x5               g069(.a(new_n158), .b(new_n151), .c(new_n137), .d(new_n147), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n161), .b(new_n165), .c(new_n133), .d(new_n156), .o1(new_n166));
  xnrc02aa1n12x5               g071(.a(\b[13] ), .b(\a[14] ), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n166), .c(new_n164), .out0(\s[14] ));
  nor042aa1n06x5               g074(.a(new_n167), .b(new_n160), .o1(new_n170));
  aoai13aa1n03x5               g075(.a(new_n170), .b(new_n165), .c(new_n133), .d(new_n156), .o1(new_n171));
  oaoi03aa1n02x5               g076(.a(\a[14] ), .b(\b[13] ), .c(new_n164), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  xorc02aa1n02x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n171), .c(new_n173), .out0(\s[15] ));
  nanp02aa1n02x5               g080(.a(new_n157), .b(new_n159), .o1(new_n176));
  aoai13aa1n03x5               g081(.a(new_n174), .b(new_n172), .c(new_n176), .d(new_n170), .o1(new_n177));
  xorc02aa1n02x5               g082(.a(\a[16] ), .b(\b[15] ), .out0(new_n178));
  inv000aa1d42x5               g083(.a(\a[15] ), .o1(new_n179));
  inv000aa1d42x5               g084(.a(\b[14] ), .o1(new_n180));
  orn002aa1n02x5               g085(.a(\a[16] ), .b(\b[15] ), .o(new_n181));
  and002aa1n02x5               g086(.a(\b[15] ), .b(\a[16] ), .o(new_n182));
  aboi22aa1n03x5               g087(.a(new_n182), .b(new_n181), .c(new_n180), .d(new_n179), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n180), .b(new_n179), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n174), .o1(new_n185));
  aoai13aa1n02x5               g090(.a(new_n184), .b(new_n185), .c(new_n171), .d(new_n173), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(new_n186), .b(new_n178), .c(new_n177), .d(new_n183), .o1(\s[16] ));
  nanp02aa1n02x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  nano32aa1n03x7               g093(.a(new_n182), .b(new_n181), .c(new_n184), .d(new_n188), .out0(new_n189));
  nano22aa1d15x5               g094(.a(new_n155), .b(new_n170), .c(new_n189), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n125), .c(new_n119), .d(new_n108), .o1(new_n191));
  nand42aa1n02x5               g096(.a(new_n170), .b(new_n189), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(\b[13] ), .b(\a[14] ), .o1(new_n193));
  oai022aa1n02x7               g098(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n194));
  nanp03aa1n02x5               g099(.a(new_n194), .b(new_n193), .c(new_n188), .o1(new_n195));
  aoai13aa1n03x5               g100(.a(new_n181), .b(new_n182), .c(new_n195), .d(new_n184), .o1(new_n196));
  oab012aa1n06x5               g101(.a(new_n196), .b(new_n159), .c(new_n192), .out0(new_n197));
  nand02aa1d06x5               g102(.a(new_n191), .b(new_n197), .o1(new_n198));
  xorc02aa1n12x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  aoi113aa1n02x5               g104(.a(new_n196), .b(new_n199), .c(new_n165), .d(new_n170), .e(new_n189), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n198), .b(new_n199), .c(new_n191), .d(new_n200), .o1(\s[17] ));
  inv000aa1d42x5               g106(.a(\a[17] ), .o1(new_n202));
  nanb02aa1n02x5               g107(.a(\b[16] ), .b(new_n202), .out0(new_n203));
  oabi12aa1n09x5               g108(.a(new_n196), .b(new_n159), .c(new_n192), .out0(new_n204));
  aoai13aa1n02x5               g109(.a(new_n199), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n205));
  nor042aa1n06x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand02aa1n08x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  norb02aa1n06x4               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n205), .c(new_n203), .out0(\s[18] ));
  and002aa1n02x5               g114(.a(new_n199), .b(new_n208), .o(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n211));
  oaoi03aa1n02x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n203), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  nor002aa1d32x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand02aa1n06x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norb02aa1d21x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n211), .c(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g123(.a(new_n216), .b(new_n212), .c(new_n198), .d(new_n210), .o1(new_n219));
  nor042aa1n06x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nand22aa1n12x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  inv000aa1d42x5               g127(.a(\a[19] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[18] ), .o1(new_n224));
  aboi22aa1n03x5               g129(.a(new_n220), .b(new_n221), .c(new_n223), .d(new_n224), .out0(new_n225));
  inv030aa1n03x5               g130(.a(new_n214), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n216), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n226), .b(new_n227), .c(new_n211), .d(new_n213), .o1(new_n228));
  aoi022aa1n03x5               g133(.a(new_n228), .b(new_n222), .c(new_n219), .d(new_n225), .o1(\s[20] ));
  nano32aa1n03x7               g134(.a(new_n227), .b(new_n199), .c(new_n222), .d(new_n208), .out0(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n231));
  nanb03aa1n12x5               g136(.a(new_n220), .b(new_n221), .c(new_n215), .out0(new_n232));
  nor042aa1n04x5               g137(.a(\b[16] ), .b(\a[17] ), .o1(new_n233));
  oai112aa1n06x5               g138(.a(new_n226), .b(new_n207), .c(new_n206), .d(new_n233), .o1(new_n234));
  aoi012aa1n12x5               g139(.a(new_n220), .b(new_n214), .c(new_n221), .o1(new_n235));
  oai012aa1d24x5               g140(.a(new_n235), .b(new_n234), .c(new_n232), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nor002aa1d32x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  nanp02aa1n04x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  norb02aa1n03x5               g144(.a(new_n239), .b(new_n238), .out0(new_n240));
  xnbna2aa1n03x5               g145(.a(new_n240), .b(new_n231), .c(new_n237), .out0(\s[21] ));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n236), .c(new_n198), .d(new_n230), .o1(new_n242));
  nor042aa1n03x5               g147(.a(\b[21] ), .b(\a[22] ), .o1(new_n243));
  nanp02aa1n04x5               g148(.a(\b[21] ), .b(\a[22] ), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  aoib12aa1n02x5               g150(.a(new_n238), .b(new_n244), .c(new_n243), .out0(new_n246));
  inv000aa1n06x5               g151(.a(new_n238), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n240), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n247), .b(new_n248), .c(new_n231), .d(new_n237), .o1(new_n249));
  aoi022aa1n02x5               g154(.a(new_n249), .b(new_n245), .c(new_n242), .d(new_n246), .o1(\s[22] ));
  inv000aa1n02x5               g155(.a(new_n230), .o1(new_n251));
  nano22aa1n02x5               g156(.a(new_n251), .b(new_n240), .c(new_n245), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n253));
  nano23aa1d15x5               g158(.a(new_n238), .b(new_n243), .c(new_n244), .d(new_n239), .out0(new_n254));
  oaoi03aa1n09x5               g159(.a(\a[22] ), .b(\b[21] ), .c(new_n247), .o1(new_n255));
  aoi012aa1d18x5               g160(.a(new_n255), .b(new_n236), .c(new_n254), .o1(new_n256));
  xorc02aa1n12x5               g161(.a(\a[23] ), .b(\b[22] ), .out0(new_n257));
  xnbna2aa1n03x5               g162(.a(new_n257), .b(new_n253), .c(new_n256), .out0(\s[23] ));
  inv000aa1d42x5               g163(.a(new_n256), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n257), .b(new_n259), .c(new_n198), .d(new_n252), .o1(new_n260));
  xorc02aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .out0(new_n261));
  nor042aa1n06x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  norp02aa1n02x5               g167(.a(new_n261), .b(new_n262), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n262), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n257), .o1(new_n265));
  aoai13aa1n02x5               g170(.a(new_n264), .b(new_n265), .c(new_n253), .d(new_n256), .o1(new_n266));
  aoi022aa1n02x5               g171(.a(new_n266), .b(new_n261), .c(new_n260), .d(new_n263), .o1(\s[24] ));
  and002aa1n12x5               g172(.a(new_n261), .b(new_n257), .o(new_n268));
  nano22aa1n02x5               g173(.a(new_n251), .b(new_n268), .c(new_n254), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n268), .b(new_n255), .c(new_n236), .d(new_n254), .o1(new_n271));
  nano22aa1n02x4               g176(.a(new_n220), .b(new_n215), .c(new_n221), .out0(new_n272));
  oai012aa1n02x5               g177(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .o1(new_n273));
  oab012aa1n02x4               g178(.a(new_n273), .b(new_n233), .c(new_n206), .out0(new_n274));
  inv000aa1n02x5               g179(.a(new_n235), .o1(new_n275));
  aoai13aa1n06x5               g180(.a(new_n254), .b(new_n275), .c(new_n274), .d(new_n272), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n255), .o1(new_n277));
  inv000aa1n06x5               g182(.a(new_n268), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[24] ), .b(\b[23] ), .c(new_n264), .carry(new_n279));
  aoai13aa1n12x5               g184(.a(new_n279), .b(new_n278), .c(new_n276), .d(new_n277), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  aoi012aa1n02x5               g188(.a(new_n283), .b(new_n270), .c(new_n281), .o1(new_n284));
  norb02aa1n02x5               g189(.a(new_n279), .b(new_n282), .out0(new_n285));
  aoi013aa1n02x4               g190(.a(new_n284), .b(new_n271), .c(new_n270), .d(new_n285), .o1(\s[25] ));
  aoai13aa1n02x5               g191(.a(new_n282), .b(new_n280), .c(new_n198), .d(new_n269), .o1(new_n287));
  tech160nm_fixorc02aa1n02p5x5 g192(.a(\a[26] ), .b(\b[25] ), .out0(new_n288));
  nor042aa1n03x5               g193(.a(\b[24] ), .b(\a[25] ), .o1(new_n289));
  norp02aa1n02x5               g194(.a(new_n288), .b(new_n289), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n289), .o1(new_n291));
  aoai13aa1n04x5               g196(.a(new_n291), .b(new_n283), .c(new_n270), .d(new_n281), .o1(new_n292));
  aoi022aa1n02x5               g197(.a(new_n292), .b(new_n288), .c(new_n287), .d(new_n290), .o1(\s[26] ));
  and002aa1n12x5               g198(.a(new_n288), .b(new_n282), .o(new_n294));
  nano32aa1n03x7               g199(.a(new_n251), .b(new_n294), .c(new_n254), .d(new_n268), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n204), .c(new_n133), .d(new_n190), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n294), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[26] ), .b(\b[25] ), .c(new_n291), .carry(new_n298));
  aoai13aa1n04x5               g203(.a(new_n298), .b(new_n297), .c(new_n271), .d(new_n279), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n299), .c(new_n198), .d(new_n295), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n298), .o1(new_n302));
  aoi112aa1n02x5               g207(.a(new_n300), .b(new_n302), .c(new_n280), .d(new_n294), .o1(new_n303));
  aobi12aa1n03x7               g208(.a(new_n301), .b(new_n303), .c(new_n296), .out0(\s[27] ));
  xorc02aa1n02x5               g209(.a(\a[28] ), .b(\b[27] ), .out0(new_n305));
  norp02aa1n02x5               g210(.a(\b[26] ), .b(\a[27] ), .o1(new_n306));
  norp02aa1n02x5               g211(.a(new_n305), .b(new_n306), .o1(new_n307));
  tech160nm_fiaoi012aa1n05x5   g212(.a(new_n302), .b(new_n280), .c(new_n294), .o1(new_n308));
  inv000aa1n03x5               g213(.a(new_n306), .o1(new_n309));
  inv000aa1n02x5               g214(.a(new_n300), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n309), .b(new_n310), .c(new_n308), .d(new_n296), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n311), .b(new_n305), .c(new_n301), .d(new_n307), .o1(\s[28] ));
  and002aa1n02x5               g217(.a(new_n305), .b(new_n300), .o(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n299), .c(new_n198), .d(new_n295), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .c(new_n309), .carry(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n308), .d(new_n296), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n316), .b(new_n318), .out0(new_n319));
  aoi022aa1n03x5               g224(.a(new_n317), .b(new_n318), .c(new_n314), .d(new_n319), .o1(\s[29] ));
  xnrb03aa1n02x5               g225(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g226(.a(new_n310), .b(new_n305), .c(new_n318), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n299), .c(new_n198), .d(new_n295), .o1(new_n323));
  inv000aa1d42x5               g228(.a(new_n322), .o1(new_n324));
  oao003aa1n02x5               g229(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .carry(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n324), .c(new_n308), .d(new_n296), .o1(new_n326));
  xorc02aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .out0(new_n327));
  norb02aa1n02x5               g232(.a(new_n325), .b(new_n327), .out0(new_n328));
  aoi022aa1n03x5               g233(.a(new_n326), .b(new_n327), .c(new_n323), .d(new_n328), .o1(\s[30] ));
  nano32aa1n06x5               g234(.a(new_n310), .b(new_n327), .c(new_n305), .d(new_n318), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n299), .c(new_n198), .d(new_n295), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[31] ), .b(\b[30] ), .out0(new_n332));
  and002aa1n02x5               g237(.a(\b[29] ), .b(\a[30] ), .o(new_n333));
  oabi12aa1n02x5               g238(.a(new_n332), .b(\a[30] ), .c(\b[29] ), .out0(new_n334));
  oab012aa1n02x4               g239(.a(new_n334), .b(new_n325), .c(new_n333), .out0(new_n335));
  inv000aa1d42x5               g240(.a(new_n330), .o1(new_n336));
  oao003aa1n02x5               g241(.a(\a[30] ), .b(\b[29] ), .c(new_n325), .carry(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n336), .c(new_n308), .d(new_n296), .o1(new_n338));
  aoi022aa1n03x5               g243(.a(new_n338), .b(new_n332), .c(new_n331), .d(new_n335), .o1(\s[31] ));
  orn002aa1n02x5               g244(.a(\a[2] ), .b(\b[1] ), .o(new_n340));
  nanp02aa1n02x5               g245(.a(\b[1] ), .b(\a[2] ), .o1(new_n341));
  nanb03aa1n02x5               g246(.a(new_n99), .b(new_n340), .c(new_n341), .out0(new_n342));
  norb02aa1n02x5               g247(.a(new_n104), .b(new_n103), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n342), .c(new_n340), .out0(\s[3] ));
  obai22aa1n02x7               g249(.a(new_n101), .b(new_n102), .c(\a[3] ), .d(\b[2] ), .out0(new_n345));
  aoi012aa1n02x5               g250(.a(new_n345), .b(new_n100), .c(new_n343), .o1(new_n346));
  oaoi13aa1n02x5               g251(.a(new_n346), .b(new_n108), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g252(.a(new_n114), .b(new_n106), .c(new_n107), .out0(\s[5] ));
  aoi012aa1n02x5               g253(.a(new_n123), .b(new_n108), .c(new_n114), .o1(new_n349));
  inv000aa1d42x5               g254(.a(new_n116), .o1(new_n350));
  nanp02aa1n02x5               g255(.a(new_n108), .b(new_n114), .o1(new_n351));
  nona32aa1n03x5               g256(.a(new_n351), .b(new_n350), .c(new_n115), .d(new_n123), .out0(new_n352));
  oai012aa1n02x5               g257(.a(new_n352), .b(new_n349), .c(new_n117), .o1(\s[6] ));
  aoi022aa1n02x5               g258(.a(new_n352), .b(new_n116), .c(new_n122), .d(new_n112), .o1(new_n354));
  nona23aa1n06x5               g259(.a(new_n352), .b(new_n112), .c(new_n111), .d(new_n350), .out0(new_n355));
  norb02aa1n02x5               g260(.a(new_n355), .b(new_n354), .out0(\s[7] ));
  norb02aa1n02x5               g261(.a(new_n109), .b(new_n110), .out0(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n357), .b(new_n355), .c(new_n122), .out0(\s[8] ));
  xorb03aa1n02x5               g263(.a(new_n133), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


