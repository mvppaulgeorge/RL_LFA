// Benchmark "adder" written by ABC on Thu Jul 18 12:16:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n330,
    new_n331, new_n333, new_n334, new_n336, new_n338, new_n339, new_n340,
    new_n342, new_n344, new_n345, new_n346, new_n348, new_n349, new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  and002aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n12x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  nor042aa1n03x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nand02aa1n03x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norb02aa1n06x5               g007(.a(new_n102), .b(new_n101), .out0(new_n103));
  nor042aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  norb02aa1n09x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nanp03aa1d12x5               g011(.a(new_n100), .b(new_n103), .c(new_n106), .o1(new_n107));
  aoi012aa1n06x5               g012(.a(new_n101), .b(new_n104), .c(new_n102), .o1(new_n108));
  oai022aa1n02x5               g013(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n109));
  nand42aa1n02x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nano22aa1n03x5               g016(.a(new_n109), .b(new_n110), .c(new_n111), .out0(new_n112));
  nand22aa1n09x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor042aa1n04x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nor042aa1n04x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nanp02aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n09x5               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  nand02aa1n02x5               g022(.a(new_n117), .b(new_n112), .o1(new_n118));
  orn002aa1n03x5               g023(.a(\a[5] ), .b(\b[4] ), .o(new_n119));
  oaoi03aa1n03x5               g024(.a(\a[6] ), .b(\b[5] ), .c(new_n119), .o1(new_n120));
  tech160nm_fiaoi012aa1n02p5x5 g025(.a(new_n115), .b(new_n114), .c(new_n113), .o1(new_n121));
  aobi12aa1n06x5               g026(.a(new_n121), .b(new_n117), .c(new_n120), .out0(new_n122));
  aoai13aa1n12x5               g027(.a(new_n122), .b(new_n118), .c(new_n107), .d(new_n108), .o1(new_n123));
  xorc02aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  nanp02aa1n03x5               g029(.a(new_n123), .b(new_n124), .o1(new_n125));
  xorc02aa1n02x5               g030(.a(\a[10] ), .b(\b[9] ), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n126), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  oa0022aa1n03x5               g032(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n128));
  nanp02aa1n02x5               g033(.a(new_n125), .b(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n03x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor002aa1n10x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nanb03aa1n02x5               g037(.a(new_n132), .b(new_n130), .c(new_n131), .out0(new_n133));
  nanb02aa1n03x5               g038(.a(new_n133), .b(new_n129), .out0(new_n134));
  inv000aa1d42x5               g039(.a(new_n132), .o1(new_n135));
  aoi022aa1n02x5               g040(.a(new_n129), .b(new_n130), .c(new_n135), .d(new_n131), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n134), .b(new_n136), .out0(\s[11] ));
  nor002aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoib12aa1n02x5               g045(.a(new_n132), .b(new_n139), .c(new_n138), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n135), .b(new_n133), .c(new_n125), .d(new_n128), .o1(new_n142));
  aoi022aa1n02x5               g047(.a(new_n134), .b(new_n141), .c(new_n142), .d(new_n140), .o1(\s[12] ));
  nano23aa1n02x5               g048(.a(new_n138), .b(new_n132), .c(new_n139), .d(new_n131), .out0(new_n144));
  and003aa1n02x5               g049(.a(new_n144), .b(new_n126), .c(new_n124), .o(new_n145));
  nano22aa1n03x5               g050(.a(new_n138), .b(new_n131), .c(new_n139), .out0(new_n146));
  nona23aa1n06x5               g051(.a(new_n146), .b(new_n130), .c(new_n128), .d(new_n132), .out0(new_n147));
  aoi012aa1n02x7               g052(.a(new_n138), .b(new_n132), .c(new_n139), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  xnrc02aa1n12x5               g054(.a(\b[12] ), .b(\a[13] ), .out0(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n149), .c(new_n123), .d(new_n145), .o1(new_n152));
  and003aa1n02x5               g057(.a(new_n147), .b(new_n150), .c(new_n148), .o(new_n153));
  aobi12aa1n02x5               g058(.a(new_n153), .b(new_n145), .c(new_n123), .out0(new_n154));
  norb02aa1n02x5               g059(.a(new_n152), .b(new_n154), .out0(\s[13] ));
  orn002aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .o(new_n156));
  xorc02aa1n12x5               g061(.a(\a[14] ), .b(\b[13] ), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n152), .c(new_n156), .out0(\s[14] ));
  xnrc02aa1n02x5               g063(.a(\b[13] ), .b(\a[14] ), .out0(new_n159));
  norp02aa1n02x5               g064(.a(new_n159), .b(new_n150), .o1(new_n160));
  aoai13aa1n06x5               g065(.a(new_n160), .b(new_n149), .c(new_n123), .d(new_n145), .o1(new_n161));
  oaoi03aa1n02x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nor002aa1n20x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand42aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n161), .c(new_n163), .out0(\s[15] ));
  aob012aa1n02x5               g072(.a(new_n166), .b(new_n161), .c(new_n163), .out0(new_n168));
  tech160nm_fixorc02aa1n03p5x5 g073(.a(\a[16] ), .b(\b[15] ), .out0(new_n169));
  inv000aa1d42x5               g074(.a(\a[16] ), .o1(new_n170));
  inv000aa1d42x5               g075(.a(\b[15] ), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n170), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  aoi012aa1n02x5               g078(.a(new_n164), .b(new_n172), .c(new_n173), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n164), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n164), .b(new_n165), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n175), .b(new_n176), .c(new_n161), .d(new_n163), .o1(new_n177));
  aoi022aa1n02x5               g082(.a(new_n177), .b(new_n169), .c(new_n168), .d(new_n174), .o1(\s[16] ));
  nona23aa1d18x5               g083(.a(new_n169), .b(new_n157), .c(new_n150), .d(new_n176), .out0(new_n179));
  nano32aa1d12x5               g084(.a(new_n179), .b(new_n144), .c(new_n126), .d(new_n124), .out0(new_n180));
  nanp02aa1n06x5               g085(.a(new_n123), .b(new_n180), .o1(new_n181));
  nanp03aa1n02x5               g086(.a(new_n172), .b(new_n165), .c(new_n173), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(\b[13] ), .b(\a[14] ), .o1(new_n183));
  oai022aa1n02x5               g088(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n184));
  oai112aa1n02x5               g089(.a(new_n184), .b(new_n183), .c(\b[14] ), .d(\a[15] ), .o1(new_n185));
  oaoi03aa1n02x5               g090(.a(new_n170), .b(new_n171), .c(new_n164), .o1(new_n186));
  oa0012aa1n02x5               g091(.a(new_n186), .b(new_n185), .c(new_n182), .o(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n179), .c(new_n147), .d(new_n148), .o1(new_n188));
  nanb02aa1n06x5               g093(.a(new_n188), .b(new_n181), .out0(new_n189));
  xorc02aa1n02x5               g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  xnrc02aa1n02x5               g095(.a(\b[16] ), .b(\a[17] ), .out0(new_n191));
  oai112aa1n02x5               g096(.a(new_n186), .b(new_n191), .c(new_n185), .d(new_n182), .o1(new_n192));
  aoib12aa1n02x5               g097(.a(new_n192), .b(new_n149), .c(new_n179), .out0(new_n193));
  aoi022aa1n02x5               g098(.a(new_n189), .b(new_n190), .c(new_n181), .d(new_n193), .o1(\s[17] ));
  nor042aa1d18x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  aoai13aa1n02x5               g101(.a(new_n190), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n197));
  nor042aa1n04x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nanp02aa1n04x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  norb02aa1n06x4               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n200), .b(new_n197), .c(new_n196), .out0(\s[18] ));
  norb02aa1n02x5               g106(.a(new_n200), .b(new_n191), .out0(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n203));
  oaoi03aa1n02x5               g108(.a(\a[18] ), .b(\b[17] ), .c(new_n196), .o1(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  nor022aa1n16x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand42aa1n20x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  norb02aa1n12x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n203), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g115(.a(new_n208), .b(new_n203), .c(new_n205), .out0(new_n211));
  norp02aa1n09x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand42aa1n10x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  inv000aa1d42x5               g119(.a(\a[19] ), .o1(new_n215));
  inv000aa1d42x5               g120(.a(\b[18] ), .o1(new_n216));
  aboi22aa1n03x5               g121(.a(new_n212), .b(new_n213), .c(new_n215), .d(new_n216), .out0(new_n217));
  inv030aa1n02x5               g122(.a(new_n206), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n208), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n218), .b(new_n219), .c(new_n203), .d(new_n205), .o1(new_n220));
  aoi022aa1n02x5               g125(.a(new_n220), .b(new_n214), .c(new_n211), .d(new_n217), .o1(\s[20] ));
  nano32aa1n03x7               g126(.a(new_n191), .b(new_n214), .c(new_n200), .d(new_n208), .out0(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n223));
  nanb03aa1n06x5               g128(.a(new_n212), .b(new_n213), .c(new_n207), .out0(new_n224));
  oai112aa1n06x5               g129(.a(new_n218), .b(new_n199), .c(new_n198), .d(new_n195), .o1(new_n225));
  aoi012aa1n09x5               g130(.a(new_n212), .b(new_n206), .c(new_n213), .o1(new_n226));
  oai012aa1n18x5               g131(.a(new_n226), .b(new_n225), .c(new_n224), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  nor002aa1n10x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  nand42aa1n02x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  norb02aa1n03x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  aob012aa1n03x5               g136(.a(new_n231), .b(new_n223), .c(new_n228), .out0(new_n232));
  nano22aa1n02x4               g137(.a(new_n212), .b(new_n207), .c(new_n213), .out0(new_n233));
  oai012aa1n02x5               g138(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .o1(new_n234));
  oab012aa1n04x5               g139(.a(new_n234), .b(new_n195), .c(new_n198), .out0(new_n235));
  inv020aa1n02x5               g140(.a(new_n226), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(new_n236), .b(new_n231), .c(new_n235), .d(new_n233), .o1(new_n237));
  aobi12aa1n02x7               g142(.a(new_n232), .b(new_n237), .c(new_n223), .out0(\s[21] ));
  nor002aa1n04x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nand42aa1n04x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  aoib12aa1n02x5               g146(.a(new_n229), .b(new_n240), .c(new_n239), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n229), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n231), .o1(new_n244));
  aoai13aa1n02x5               g149(.a(new_n243), .b(new_n244), .c(new_n223), .d(new_n228), .o1(new_n245));
  aoi022aa1n03x5               g150(.a(new_n245), .b(new_n241), .c(new_n232), .d(new_n242), .o1(\s[22] ));
  inv000aa1n02x5               g151(.a(new_n222), .o1(new_n247));
  nano22aa1n02x4               g152(.a(new_n247), .b(new_n231), .c(new_n241), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n249));
  nano23aa1n06x5               g154(.a(new_n229), .b(new_n239), .c(new_n240), .d(new_n230), .out0(new_n250));
  aoi012aa1n02x5               g155(.a(new_n239), .b(new_n229), .c(new_n240), .o1(new_n251));
  inv020aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  aoi012aa1n02x5               g157(.a(new_n252), .b(new_n227), .c(new_n250), .o1(new_n253));
  xorc02aa1n12x5               g158(.a(\a[23] ), .b(\b[22] ), .out0(new_n254));
  aob012aa1n03x5               g159(.a(new_n254), .b(new_n249), .c(new_n253), .out0(new_n255));
  aoi112aa1n02x5               g160(.a(new_n254), .b(new_n252), .c(new_n227), .d(new_n250), .o1(new_n256));
  aobi12aa1n02x7               g161(.a(new_n255), .b(new_n256), .c(new_n249), .out0(\s[23] ));
  xorc02aa1n02x5               g162(.a(\a[24] ), .b(\b[23] ), .out0(new_n258));
  nor042aa1n06x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  norp02aa1n02x5               g164(.a(new_n258), .b(new_n259), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n259), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n254), .o1(new_n262));
  aoai13aa1n02x5               g167(.a(new_n261), .b(new_n262), .c(new_n249), .d(new_n253), .o1(new_n263));
  aoi022aa1n03x5               g168(.a(new_n263), .b(new_n258), .c(new_n255), .d(new_n260), .o1(\s[24] ));
  and002aa1n12x5               g169(.a(new_n258), .b(new_n254), .o(new_n265));
  nano22aa1n03x5               g170(.a(new_n247), .b(new_n265), .c(new_n250), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n250), .b(new_n236), .c(new_n235), .d(new_n233), .o1(new_n268));
  inv040aa1n02x5               g173(.a(new_n265), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[24] ), .b(\b[23] ), .c(new_n261), .carry(new_n270));
  aoai13aa1n12x5               g175(.a(new_n270), .b(new_n269), .c(new_n268), .d(new_n251), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  xorc02aa1n12x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  aob012aa1n03x5               g178(.a(new_n273), .b(new_n267), .c(new_n272), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n265), .b(new_n252), .c(new_n227), .d(new_n250), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n273), .o1(new_n276));
  and003aa1n02x5               g181(.a(new_n275), .b(new_n276), .c(new_n270), .o(new_n277));
  aobi12aa1n02x7               g182(.a(new_n274), .b(new_n277), .c(new_n267), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  nor042aa1n06x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n280), .o1(new_n282));
  aoai13aa1n02x5               g187(.a(new_n282), .b(new_n276), .c(new_n267), .d(new_n272), .o1(new_n283));
  aoi022aa1n02x5               g188(.a(new_n283), .b(new_n279), .c(new_n274), .d(new_n281), .o1(\s[26] ));
  and002aa1n12x5               g189(.a(new_n279), .b(new_n273), .o(new_n285));
  nano32aa1n03x7               g190(.a(new_n247), .b(new_n285), .c(new_n250), .d(new_n265), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n188), .c(new_n123), .d(new_n180), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[26] ), .b(\b[25] ), .c(new_n282), .carry(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n288), .c(new_n275), .d(new_n270), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n290), .c(new_n189), .d(new_n286), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n289), .o1(new_n293));
  aoi112aa1n02x5               g198(.a(new_n291), .b(new_n293), .c(new_n271), .d(new_n285), .o1(new_n294));
  aobi12aa1n03x7               g199(.a(new_n292), .b(new_n294), .c(new_n287), .out0(\s[27] ));
  xorc02aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .out0(new_n296));
  norp02aa1n02x5               g201(.a(\b[26] ), .b(\a[27] ), .o1(new_n297));
  norp02aa1n02x5               g202(.a(new_n296), .b(new_n297), .o1(new_n298));
  aoi012aa1n06x5               g203(.a(new_n293), .b(new_n271), .c(new_n285), .o1(new_n299));
  inv000aa1n03x5               g204(.a(new_n297), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n291), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n300), .b(new_n301), .c(new_n299), .d(new_n287), .o1(new_n302));
  aoi022aa1n03x5               g207(.a(new_n302), .b(new_n296), .c(new_n292), .d(new_n298), .o1(\s[28] ));
  and002aa1n02x5               g208(.a(new_n296), .b(new_n291), .o(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n290), .c(new_n189), .d(new_n286), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[28] ), .b(\b[27] ), .c(new_n300), .carry(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n306), .c(new_n299), .d(new_n287), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n307), .b(new_n309), .out0(new_n310));
  aoi022aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n305), .d(new_n310), .o1(\s[29] ));
  xnrb03aa1n02x5               g216(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g217(.a(new_n301), .b(new_n296), .c(new_n309), .out0(new_n313));
  aoai13aa1n06x5               g218(.a(new_n313), .b(new_n290), .c(new_n189), .d(new_n286), .o1(new_n314));
  inv000aa1n02x5               g219(.a(new_n313), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[29] ), .b(\b[28] ), .c(new_n307), .carry(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n299), .d(new_n287), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n316), .b(new_n318), .out0(new_n319));
  aoi022aa1n03x5               g224(.a(new_n317), .b(new_n318), .c(new_n314), .d(new_n319), .o1(\s[30] ));
  nano32aa1n06x5               g225(.a(new_n301), .b(new_n318), .c(new_n296), .d(new_n309), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n290), .c(new_n189), .d(new_n286), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[31] ), .b(\b[30] ), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n316), .carry(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(new_n325));
  inv000aa1d42x5               g230(.a(new_n321), .o1(new_n326));
  aoai13aa1n03x5               g231(.a(new_n324), .b(new_n326), .c(new_n299), .d(new_n287), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n323), .c(new_n322), .d(new_n325), .o1(\s[31] ));
  orn002aa1n02x5               g233(.a(\a[2] ), .b(\b[1] ), .o(new_n329));
  nanp02aa1n02x5               g234(.a(\b[1] ), .b(\a[2] ), .o1(new_n330));
  nanb03aa1n02x5               g235(.a(new_n99), .b(new_n330), .c(new_n329), .out0(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n106), .b(new_n331), .c(new_n329), .out0(\s[3] ));
  aoai13aa1n02x5               g237(.a(new_n103), .b(new_n104), .c(new_n100), .d(new_n105), .o1(new_n333));
  aoi112aa1n02x5               g238(.a(new_n104), .b(new_n103), .c(new_n100), .d(new_n106), .o1(new_n334));
  norb02aa1n02x5               g239(.a(new_n333), .b(new_n334), .out0(\s[4] ));
  xorc02aa1n02x5               g240(.a(\a[5] ), .b(\b[4] ), .out0(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n336), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  aob012aa1n02x5               g242(.a(new_n336), .b(new_n107), .c(new_n108), .out0(new_n338));
  xorc02aa1n02x5               g243(.a(\a[6] ), .b(\b[5] ), .out0(new_n339));
  nanb03aa1n02x5               g244(.a(new_n109), .b(new_n338), .c(new_n110), .out0(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n339), .c(new_n119), .d(new_n338), .o1(\s[6] ));
  norb02aa1n02x5               g246(.a(new_n116), .b(new_n114), .out0(new_n342));
  xobna2aa1n03x5               g247(.a(new_n342), .b(new_n340), .c(new_n110), .out0(\s[7] ));
  aoi013aa1n02x4               g248(.a(new_n114), .b(new_n340), .c(new_n110), .d(new_n342), .o1(new_n344));
  norb02aa1n02x5               g249(.a(new_n113), .b(new_n115), .out0(new_n345));
  aoi113aa1n02x5               g250(.a(new_n345), .b(new_n114), .c(new_n340), .d(new_n342), .e(new_n110), .o1(new_n346));
  aoib12aa1n02x5               g251(.a(new_n346), .b(new_n345), .c(new_n344), .out0(\s[8] ));
  aoi012aa1n02x5               g252(.a(new_n118), .b(new_n107), .c(new_n108), .o1(new_n348));
  tech160nm_fiao0012aa1n02p5x5 g253(.a(new_n115), .b(new_n114), .c(new_n113), .o(new_n349));
  aoi112aa1n02x5               g254(.a(new_n124), .b(new_n349), .c(new_n117), .d(new_n120), .o1(new_n350));
  aboi22aa1n03x5               g255(.a(new_n348), .b(new_n350), .c(new_n123), .d(new_n124), .out0(\s[9] ));
endmodule


