// Benchmark "adder" written by ABC on Thu Jul 18 00:08:47 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n216, new_n217, new_n218, new_n219, new_n220, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n310, new_n311, new_n312, new_n314, new_n315, new_n318, new_n320,
    new_n321;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  and002aa1n24x5               g002(.a(\b[3] ), .b(\a[4] ), .o(new_n98));
  nand22aa1n06x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nand42aa1d28x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nor002aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  norb03aa1n12x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  nor002aa1d32x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n16x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb03aa1d24x5               g009(.a(new_n103), .b(new_n104), .c(new_n100), .out0(new_n105));
  oab012aa1n04x5               g010(.a(new_n103), .b(\a[4] ), .c(\b[3] ), .out0(new_n106));
  oaoi13aa1n12x5               g011(.a(new_n98), .b(new_n106), .c(new_n102), .d(new_n105), .o1(new_n107));
  nor002aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand42aa1d28x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  norb02aa1n06x4               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  nand42aa1d28x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  norp02aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  norb02aa1n03x4               g017(.a(new_n111), .b(new_n112), .out0(new_n113));
  tech160nm_fixnrc02aa1n05x5   g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  xnrc02aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .out0(new_n115));
  nano23aa1n09x5               g020(.a(new_n115), .b(new_n114), .c(new_n113), .d(new_n110), .out0(new_n116));
  nand22aa1n03x5               g021(.a(new_n107), .b(new_n116), .o1(new_n117));
  xorc02aa1n12x5               g022(.a(\a[7] ), .b(\b[6] ), .out0(new_n118));
  nano22aa1n03x7               g023(.a(new_n108), .b(new_n109), .c(new_n111), .out0(new_n119));
  oai022aa1d18x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  nor042aa1n04x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  inv030aa1n02x5               g026(.a(new_n121), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  aoi013aa1n02x4               g028(.a(new_n123), .b(new_n119), .c(new_n118), .d(new_n120), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n97), .b(new_n126), .c(new_n117), .d(new_n124), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xorc02aa1n12x5               g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  oaoi03aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n130));
  nor042aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nand22aa1n09x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  aoai13aa1n06x5               g038(.a(new_n133), .b(new_n130), .c(new_n127), .d(new_n129), .o1(new_n134));
  aoi112aa1n02x5               g039(.a(new_n133), .b(new_n130), .c(new_n127), .d(new_n129), .o1(new_n135));
  norb02aa1n02x7               g040(.a(new_n134), .b(new_n135), .out0(\s[11] ));
  inv040aa1n02x5               g041(.a(new_n131), .o1(new_n137));
  nor042aa1n04x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1d06x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aobi12aa1n02x7               g045(.a(new_n140), .b(new_n134), .c(new_n137), .out0(new_n141));
  nona22aa1n02x5               g046(.a(new_n134), .b(new_n140), .c(new_n131), .out0(new_n142));
  norb02aa1n03x4               g047(.a(new_n142), .b(new_n141), .out0(\s[12] ));
  nanp03aa1n06x5               g048(.a(new_n119), .b(new_n118), .c(new_n120), .o1(new_n144));
  nanb02aa1n09x5               g049(.a(new_n123), .b(new_n144), .out0(new_n145));
  nano23aa1d15x5               g050(.a(new_n131), .b(new_n138), .c(new_n139), .d(new_n132), .out0(new_n146));
  nanp03aa1d12x5               g051(.a(new_n146), .b(new_n125), .c(new_n129), .o1(new_n147));
  inv040aa1n02x5               g052(.a(new_n147), .o1(new_n148));
  aoai13aa1n06x5               g053(.a(new_n148), .b(new_n145), .c(new_n107), .d(new_n116), .o1(new_n149));
  oaoi03aa1n02x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .o1(new_n150));
  aoi012aa1n06x5               g055(.a(new_n150), .b(new_n146), .c(new_n130), .o1(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[12] ), .b(\a[13] ), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n149), .c(new_n151), .out0(\s[13] ));
  inv040aa1d32x5               g059(.a(\a[14] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n149), .b(new_n151), .o1(new_n156));
  nor042aa1d18x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n03x5               g062(.a(new_n157), .b(new_n156), .c(new_n153), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(new_n155), .out0(\s[14] ));
  xnrc02aa1n02x5               g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  nor002aa1n02x5               g065(.a(new_n160), .b(new_n152), .o1(new_n161));
  inv000aa1n02x5               g066(.a(new_n161), .o1(new_n162));
  inv040aa1d32x5               g067(.a(\b[13] ), .o1(new_n163));
  oao003aa1n09x5               g068(.a(new_n155), .b(new_n163), .c(new_n157), .carry(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n04x5               g070(.a(new_n165), .b(new_n162), .c(new_n149), .d(new_n151), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor022aa1n06x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n06x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nor042aa1n03x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand02aa1n06x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n168), .b(new_n172), .c(new_n166), .d(new_n169), .o1(new_n174));
  norb02aa1n02x7               g079(.a(new_n173), .b(new_n174), .out0(\s[16] ));
  nano23aa1d12x5               g080(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n176));
  nona22aa1n09x5               g081(.a(new_n176), .b(new_n160), .c(new_n152), .out0(new_n177));
  nor042aa1n06x5               g082(.a(new_n177), .b(new_n147), .o1(new_n178));
  aoai13aa1n12x5               g083(.a(new_n178), .b(new_n145), .c(new_n107), .d(new_n116), .o1(new_n179));
  tech160nm_fiaoi012aa1n03p5x5 g084(.a(new_n170), .b(new_n168), .c(new_n171), .o1(new_n180));
  aob012aa1d15x5               g085(.a(new_n180), .b(new_n176), .c(new_n164), .out0(new_n181));
  oab012aa1n12x5               g086(.a(new_n181), .b(new_n151), .c(new_n177), .out0(new_n182));
  nand02aa1d08x5               g087(.a(new_n179), .b(new_n182), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[18] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[17] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[16] ), .o1(new_n187));
  oaoi03aa1n03x5               g092(.a(new_n186), .b(new_n187), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  xroi22aa1d06x4               g094(.a(new_n186), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n190));
  oai022aa1d18x5               g095(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n191));
  oaib12aa1n18x5               g096(.a(new_n191), .b(new_n185), .c(\b[17] ), .out0(new_n192));
  inv040aa1n02x5               g097(.a(new_n192), .o1(new_n193));
  nor022aa1n16x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand02aa1d06x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n193), .c(new_n183), .d(new_n190), .o1(new_n197));
  aoi112aa1n02x5               g102(.a(new_n196), .b(new_n193), .c(new_n183), .d(new_n190), .o1(new_n198));
  norb02aa1n02x7               g103(.a(new_n197), .b(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  orn002aa1n02x5               g105(.a(\a[19] ), .b(\b[18] ), .o(new_n201));
  nor002aa1d32x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nand02aa1d06x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  aobi12aa1n06x5               g109(.a(new_n204), .b(new_n197), .c(new_n201), .out0(new_n205));
  nona22aa1n02x5               g110(.a(new_n197), .b(new_n204), .c(new_n194), .out0(new_n206));
  norb02aa1n03x4               g111(.a(new_n206), .b(new_n205), .out0(\s[20] ));
  nano23aa1n03x7               g112(.a(new_n194), .b(new_n202), .c(new_n203), .d(new_n195), .out0(new_n208));
  nanp02aa1n02x5               g113(.a(new_n190), .b(new_n208), .o1(new_n209));
  nona23aa1n09x5               g114(.a(new_n203), .b(new_n195), .c(new_n194), .d(new_n202), .out0(new_n210));
  tech160nm_fiaoi012aa1n05x5   g115(.a(new_n202), .b(new_n194), .c(new_n203), .o1(new_n211));
  oai012aa1n12x5               g116(.a(new_n211), .b(new_n210), .c(new_n192), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  aoai13aa1n04x5               g118(.a(new_n213), .b(new_n209), .c(new_n179), .d(new_n182), .o1(new_n214));
  xorb03aa1n02x5               g119(.a(new_n214), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  xorc02aa1n02x5               g121(.a(\a[21] ), .b(\b[20] ), .out0(new_n217));
  xorc02aa1n02x5               g122(.a(\a[22] ), .b(\b[21] ), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n216), .c(new_n214), .d(new_n217), .o1(new_n219));
  aoi112aa1n03x4               g124(.a(new_n216), .b(new_n218), .c(new_n214), .d(new_n217), .o1(new_n220));
  norb02aa1n02x7               g125(.a(new_n219), .b(new_n220), .out0(\s[22] ));
  inv000aa1d42x5               g126(.a(\a[21] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\a[22] ), .o1(new_n223));
  xroi22aa1d06x4               g128(.a(new_n222), .b(\b[20] ), .c(new_n223), .d(\b[21] ), .out0(new_n224));
  nanp03aa1n03x5               g129(.a(new_n224), .b(new_n190), .c(new_n208), .o1(new_n225));
  inv000aa1d42x5               g130(.a(\b[21] ), .o1(new_n226));
  oaoi03aa1n09x5               g131(.a(new_n223), .b(new_n226), .c(new_n216), .o1(new_n227));
  inv000aa1n02x5               g132(.a(new_n227), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n212), .c(new_n224), .o1(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n225), .c(new_n179), .d(new_n182), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .o1(new_n232));
  tech160nm_fixorc02aa1n02p5x5 g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  xorc02aa1n02x5               g138(.a(\a[24] ), .b(\b[23] ), .out0(new_n234));
  aoai13aa1n03x5               g139(.a(new_n234), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n232), .b(new_n234), .c(new_n230), .d(new_n233), .o1(new_n236));
  norb02aa1n02x7               g141(.a(new_n235), .b(new_n236), .out0(\s[24] ));
  and002aa1n06x5               g142(.a(new_n234), .b(new_n233), .o(new_n238));
  inv000aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  nano32aa1n02x4               g144(.a(new_n239), .b(new_n224), .c(new_n190), .d(new_n208), .out0(new_n240));
  inv020aa1n02x5               g145(.a(new_n211), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n224), .b(new_n241), .c(new_n208), .d(new_n193), .o1(new_n242));
  aoi112aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n243));
  oab012aa1n02x4               g148(.a(new_n243), .b(\a[24] ), .c(\b[23] ), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n239), .c(new_n242), .d(new_n227), .o1(new_n245));
  xorc02aa1n02x5               g150(.a(\a[25] ), .b(\b[24] ), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n245), .c(new_n183), .d(new_n240), .o1(new_n247));
  aoi112aa1n02x5               g152(.a(new_n246), .b(new_n245), .c(new_n183), .d(new_n240), .o1(new_n248));
  norb02aa1n02x7               g153(.a(new_n247), .b(new_n248), .out0(\s[25] ));
  nor042aa1n03x5               g154(.a(\b[24] ), .b(\a[25] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  xorc02aa1n02x5               g156(.a(\a[26] ), .b(\b[25] ), .out0(new_n252));
  aobi12aa1n06x5               g157(.a(new_n252), .b(new_n247), .c(new_n251), .out0(new_n253));
  nona22aa1n02x5               g158(.a(new_n247), .b(new_n252), .c(new_n250), .out0(new_n254));
  norb02aa1n03x4               g159(.a(new_n254), .b(new_n253), .out0(\s[26] ));
  inv000aa1d42x5               g160(.a(new_n98), .o1(new_n256));
  oaih12aa1n02x5               g161(.a(new_n106), .b(new_n102), .c(new_n105), .o1(new_n257));
  nanp02aa1n03x5               g162(.a(new_n257), .b(new_n256), .o1(new_n258));
  nanb02aa1n02x5               g163(.a(new_n108), .b(new_n109), .out0(new_n259));
  nona23aa1n02x4               g164(.a(new_n113), .b(new_n118), .c(new_n114), .d(new_n259), .out0(new_n260));
  oai012aa1n02x7               g165(.a(new_n124), .b(new_n258), .c(new_n260), .o1(new_n261));
  oabi12aa1n03x5               g166(.a(new_n181), .b(new_n151), .c(new_n177), .out0(new_n262));
  inv000aa1d42x5               g167(.a(\a[25] ), .o1(new_n263));
  inv020aa1n04x5               g168(.a(\a[26] ), .o1(new_n264));
  xroi22aa1d06x4               g169(.a(new_n263), .b(\b[24] ), .c(new_n264), .d(\b[25] ), .out0(new_n265));
  nano22aa1n03x7               g170(.a(new_n225), .b(new_n238), .c(new_n265), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n262), .c(new_n261), .d(new_n178), .o1(new_n267));
  oao003aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .c(new_n251), .carry(new_n268));
  aobi12aa1n06x5               g173(.a(new_n268), .b(new_n245), .c(new_n265), .out0(new_n269));
  xorc02aa1n12x5               g174(.a(\a[27] ), .b(\b[26] ), .out0(new_n270));
  xnbna2aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n267), .out0(\s[27] ));
  norp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  inv040aa1n03x5               g177(.a(new_n272), .o1(new_n273));
  inv020aa1n03x5               g178(.a(new_n266), .o1(new_n274));
  aoi012aa1n06x5               g179(.a(new_n274), .b(new_n179), .c(new_n182), .o1(new_n275));
  aoai13aa1n02x7               g180(.a(new_n238), .b(new_n228), .c(new_n212), .d(new_n224), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n265), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n268), .b(new_n277), .c(new_n276), .d(new_n244), .o1(new_n278));
  oaih12aa1n02x5               g183(.a(new_n270), .b(new_n278), .c(new_n275), .o1(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[27] ), .b(\a[28] ), .out0(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n279), .c(new_n273), .o1(new_n281));
  aobi12aa1n02x7               g186(.a(new_n270), .b(new_n269), .c(new_n267), .out0(new_n282));
  nano22aa1n03x5               g187(.a(new_n282), .b(new_n273), .c(new_n280), .out0(new_n283));
  norp02aa1n03x5               g188(.a(new_n281), .b(new_n283), .o1(\s[28] ));
  norb02aa1n02x5               g189(.a(new_n270), .b(new_n280), .out0(new_n285));
  oaih12aa1n02x5               g190(.a(new_n285), .b(new_n278), .c(new_n275), .o1(new_n286));
  oao003aa1n02x5               g191(.a(\a[28] ), .b(\b[27] ), .c(new_n273), .carry(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  tech160nm_fiaoi012aa1n02p5x5 g193(.a(new_n288), .b(new_n286), .c(new_n287), .o1(new_n289));
  aobi12aa1n02x7               g194(.a(new_n285), .b(new_n269), .c(new_n267), .out0(new_n290));
  nano22aa1n03x5               g195(.a(new_n290), .b(new_n287), .c(new_n288), .out0(new_n291));
  norp02aa1n03x5               g196(.a(new_n289), .b(new_n291), .o1(\s[29] ));
  xorb03aa1n02x5               g197(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g198(.a(new_n270), .b(new_n288), .c(new_n280), .out0(new_n294));
  oaih12aa1n02x5               g199(.a(new_n294), .b(new_n278), .c(new_n275), .o1(new_n295));
  oao003aa1n02x5               g200(.a(\a[29] ), .b(\b[28] ), .c(new_n287), .carry(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[29] ), .b(\a[30] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n295), .c(new_n296), .o1(new_n298));
  aobi12aa1n02x7               g203(.a(new_n294), .b(new_n269), .c(new_n267), .out0(new_n299));
  nano22aa1n03x5               g204(.a(new_n299), .b(new_n296), .c(new_n297), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n298), .b(new_n300), .o1(\s[30] ));
  norb02aa1n02x5               g206(.a(new_n294), .b(new_n297), .out0(new_n302));
  aobi12aa1n02x7               g207(.a(new_n302), .b(new_n269), .c(new_n267), .out0(new_n303));
  oao003aa1n02x5               g208(.a(\a[30] ), .b(\b[29] ), .c(new_n296), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[30] ), .b(\a[31] ), .out0(new_n305));
  nano22aa1n03x5               g210(.a(new_n303), .b(new_n304), .c(new_n305), .out0(new_n306));
  oaih12aa1n02x5               g211(.a(new_n302), .b(new_n278), .c(new_n275), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n305), .b(new_n307), .c(new_n304), .o1(new_n308));
  norp02aa1n03x5               g213(.a(new_n308), .b(new_n306), .o1(\s[31] ));
  norp02aa1n02x5               g214(.a(new_n102), .b(new_n105), .o1(new_n310));
  oai012aa1n02x5               g215(.a(new_n100), .b(new_n101), .c(new_n99), .o1(new_n311));
  oaib12aa1n02x5               g216(.a(new_n311), .b(new_n103), .c(new_n104), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n312), .b(new_n310), .out0(\s[3] ));
  xorc02aa1n02x5               g218(.a(\a[4] ), .b(\b[3] ), .out0(new_n314));
  norp03aa1n02x5               g219(.a(new_n310), .b(new_n314), .c(new_n103), .o1(new_n315));
  oaoi13aa1n02x5               g220(.a(new_n315), .b(new_n107), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g221(.a(new_n114), .b(new_n257), .c(new_n256), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g222(.a(\a[5] ), .b(\b[4] ), .c(new_n258), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi13aa1n02x5               g224(.a(new_n118), .b(new_n111), .c(new_n318), .d(new_n112), .o1(new_n320));
  oai112aa1n02x5               g225(.a(new_n111), .b(new_n118), .c(new_n318), .d(new_n112), .o1(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(\s[7] ));
  xnbna2aa1n03x5               g227(.a(new_n110), .b(new_n321), .c(new_n122), .out0(\s[8] ));
  xnbna2aa1n03x5               g228(.a(new_n125), .b(new_n117), .c(new_n124), .out0(\s[9] ));
endmodule


