// Benchmark "adder" written by ABC on Thu Jul 11 12:13:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n325, new_n327,
    new_n328, new_n329, new_n331, new_n332;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  160nm_ficinv00aa1n08x5       g004(.clk(\a[9] ), .clkout(new_n100));
  160nm_ficinv00aa1n08x5       g005(.clk(\b[8] ), .clkout(new_n101));
  nanp02aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[8] ), .b(\a[9] ), .o1(new_n103));
  160nm_ficinv00aa1n08x5       g008(.clk(\a[2] ), .clkout(new_n104));
  160nm_ficinv00aa1n08x5       g009(.clk(\b[1] ), .clkout(new_n105));
  nanp02aa1n02x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  oaoi03aa1n02x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nona23aa1n02x4               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  aoi012aa1n02x5               g017(.a(new_n108), .b(new_n110), .c(new_n109), .o1(new_n113));
  oai012aa1n02x5               g018(.a(new_n113), .b(new_n112), .c(new_n107), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  norp02aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  norp02aa1n02x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nona23aa1n02x4               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  xnrc02aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .out0(new_n123));
  norp03aa1n02x5               g028(.a(new_n122), .b(new_n123), .c(new_n117), .o1(new_n124));
  oai012aa1n02x5               g029(.a(new_n119), .b(new_n120), .c(new_n118), .o1(new_n125));
  orn002aa1n02x5               g030(.a(\a[5] ), .b(\b[4] ), .o(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[6] ), .b(\b[5] ), .c(new_n126), .o1(new_n127));
  oaib12aa1n02x5               g032(.a(new_n125), .b(new_n122), .c(new_n127), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n103), .b(new_n128), .c(new_n114), .d(new_n124), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n99), .b(new_n129), .c(new_n102), .out0(\s[10] ));
  160nm_ficinv00aa1n08x5       g035(.clk(new_n97), .clkout(new_n131));
  160nm_ficinv00aa1n08x5       g036(.clk(new_n98), .clkout(new_n132));
  aoai13aa1n02x5               g037(.a(new_n131), .b(new_n132), .c(new_n129), .d(new_n102), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  norp02aa1n02x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  norp02aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoi112aa1n02x5               g045(.a(new_n140), .b(new_n135), .c(new_n133), .d(new_n137), .o1(new_n141));
  aoai13aa1n02x5               g046(.a(new_n140), .b(new_n135), .c(new_n133), .d(new_n137), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(\s[12] ));
  oao003aa1n02x5               g048(.a(new_n104), .b(new_n105), .c(new_n106), .carry(new_n144));
  nano23aa1n02x4               g049(.a(new_n108), .b(new_n110), .c(new_n111), .d(new_n109), .out0(new_n145));
  aobi12aa1n02x5               g050(.a(new_n113), .b(new_n145), .c(new_n144), .out0(new_n146));
  nano23aa1n02x4               g051(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n147));
  nona22aa1n02x4               g052(.a(new_n147), .b(new_n123), .c(new_n117), .out0(new_n148));
  aobi12aa1n02x5               g053(.a(new_n125), .b(new_n147), .c(new_n127), .out0(new_n149));
  oai012aa1n02x5               g054(.a(new_n149), .b(new_n146), .c(new_n148), .o1(new_n150));
  nona23aa1n02x4               g055(.a(new_n139), .b(new_n136), .c(new_n135), .d(new_n138), .out0(new_n151));
  nano32aa1n02x4               g056(.a(new_n151), .b(new_n99), .c(new_n102), .d(new_n103), .out0(new_n152));
  oai012aa1n02x5               g057(.a(new_n139), .b(new_n138), .c(new_n135), .o1(new_n153));
  aoai13aa1n02x5               g058(.a(new_n98), .b(new_n97), .c(new_n100), .d(new_n101), .o1(new_n154));
  oai012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n155), .b(new_n150), .c(new_n152), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n02x5               g062(.a(\a[13] ), .b(\b[12] ), .c(new_n156), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  aoai13aa1n02x5               g064(.a(new_n152), .b(new_n128), .c(new_n114), .d(new_n124), .o1(new_n160));
  160nm_ficinv00aa1n08x5       g065(.clk(new_n155), .clkout(new_n161));
  norp02aa1n02x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nona23aa1n02x4               g070(.a(new_n165), .b(new_n163), .c(new_n162), .d(new_n164), .out0(new_n166));
  oai012aa1n02x5               g071(.a(new_n165), .b(new_n164), .c(new_n162), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n166), .c(new_n160), .d(new_n161), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  xorc02aa1n02x5               g075(.a(\a[15] ), .b(\b[14] ), .out0(new_n171));
  xorc02aa1n02x5               g076(.a(\a[16] ), .b(\b[15] ), .out0(new_n172));
  aoi112aa1n02x5               g077(.a(new_n172), .b(new_n170), .c(new_n168), .d(new_n171), .o1(new_n173));
  aoai13aa1n02x5               g078(.a(new_n172), .b(new_n170), .c(new_n168), .d(new_n171), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(\s[16] ));
  xorc02aa1n02x5               g080(.a(\a[9] ), .b(\b[8] ), .out0(new_n176));
  nanp03aa1n02x5               g081(.a(new_n137), .b(new_n99), .c(new_n140), .o1(new_n177));
  nano23aa1n02x4               g082(.a(new_n162), .b(new_n164), .c(new_n165), .d(new_n163), .out0(new_n178));
  nanp02aa1n02x5               g083(.a(new_n172), .b(new_n171), .o1(new_n179));
  nano23aa1n02x4               g084(.a(new_n179), .b(new_n177), .c(new_n178), .d(new_n176), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n128), .c(new_n114), .d(new_n124), .o1(new_n181));
  xnrc02aa1n02x5               g086(.a(\b[14] ), .b(\a[15] ), .out0(new_n182));
  xnrc02aa1n02x5               g087(.a(\b[15] ), .b(\a[16] ), .out0(new_n183));
  norp03aa1n02x5               g088(.a(new_n166), .b(new_n183), .c(new_n182), .o1(new_n184));
  aoi112aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n185));
  norp02aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  160nm_ficinv00aa1n08x5       g091(.clk(new_n186), .clkout(new_n187));
  oai013aa1n02x4               g092(.a(new_n187), .b(new_n182), .c(new_n183), .d(new_n167), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(new_n188), .b(new_n185), .c(new_n155), .d(new_n184), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n181), .b(new_n189), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g096(.clk(\a[18] ), .clkout(new_n192));
  160nm_ficinv00aa1n08x5       g097(.clk(\a[17] ), .clkout(new_n193));
  160nm_ficinv00aa1n08x5       g098(.clk(\b[16] ), .clkout(new_n194));
  oaoi03aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d04x5               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  160nm_ficinv00aa1n08x5       g102(.clk(new_n197), .clkout(new_n198));
  oai022aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n199));
  oaib12aa1n02x5               g104(.a(new_n199), .b(new_n192), .c(\b[17] ), .out0(new_n200));
  aoai13aa1n02x5               g105(.a(new_n200), .b(new_n198), .c(new_n181), .d(new_n189), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanp02aa1n02x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  160nm_ficinv00aa1n08x5       g110(.clk(\b[19] ), .clkout(new_n206));
  nanb02aa1n02x5               g111(.a(\a[20] ), .b(new_n206), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  aoi122aa1n02x5               g113(.a(new_n204), .b(new_n207), .c(new_n208), .d(new_n201), .e(new_n205), .o1(new_n209));
  160nm_ficinv00aa1n08x5       g114(.clk(new_n204), .clkout(new_n210));
  nanb02aa1n02x5               g115(.a(new_n204), .b(new_n205), .out0(new_n211));
  160nm_ficinv00aa1n08x5       g116(.clk(new_n211), .clkout(new_n212));
  nanp02aa1n02x5               g117(.a(new_n201), .b(new_n212), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(new_n207), .b(new_n208), .o1(new_n214));
  aoi012aa1n02x5               g119(.a(new_n214), .b(new_n213), .c(new_n210), .o1(new_n215));
  norp02aa1n02x5               g120(.a(new_n215), .b(new_n209), .o1(\s[20] ));
  norp02aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nona23aa1n02x4               g122(.a(new_n208), .b(new_n205), .c(new_n204), .d(new_n217), .out0(new_n218));
  160nm_ficinv00aa1n08x5       g123(.clk(new_n218), .clkout(new_n219));
  nanp02aa1n02x5               g124(.a(new_n197), .b(new_n219), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(new_n204), .b(new_n208), .o1(new_n221));
  norp03aa1n02x5               g126(.a(new_n200), .b(new_n211), .c(new_n214), .o1(new_n222));
  nano22aa1n02x4               g127(.a(new_n222), .b(new_n207), .c(new_n221), .out0(new_n223));
  aoai13aa1n02x5               g128(.a(new_n223), .b(new_n220), .c(new_n181), .d(new_n189), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  xorc02aa1n02x5               g131(.a(\a[21] ), .b(\b[20] ), .out0(new_n227));
  xorc02aa1n02x5               g132(.a(\a[22] ), .b(\b[21] ), .out0(new_n228));
  aoi112aa1n02x5               g133(.a(new_n226), .b(new_n228), .c(new_n224), .d(new_n227), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n228), .b(new_n226), .c(new_n224), .d(new_n227), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(\s[22] ));
  160nm_ficinv00aa1n08x5       g136(.clk(\a[21] ), .clkout(new_n232));
  160nm_ficinv00aa1n08x5       g137(.clk(\a[22] ), .clkout(new_n233));
  xroi22aa1d04x5               g138(.a(new_n232), .b(\b[20] ), .c(new_n233), .d(\b[21] ), .out0(new_n234));
  nanp03aa1n02x5               g139(.a(new_n234), .b(new_n197), .c(new_n219), .o1(new_n235));
  oai112aa1n02x5               g140(.a(new_n221), .b(new_n207), .c(new_n218), .d(new_n200), .o1(new_n236));
  160nm_ficinv00aa1n08x5       g141(.clk(\b[21] ), .clkout(new_n237));
  oaoi03aa1n02x5               g142(.a(new_n233), .b(new_n237), .c(new_n226), .o1(new_n238));
  160nm_ficinv00aa1n08x5       g143(.clk(new_n238), .clkout(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n236), .c(new_n234), .o1(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n235), .c(new_n181), .d(new_n189), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  xorc02aa1n02x5               g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  xorc02aa1n02x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoi112aa1n02x5               g150(.a(new_n243), .b(new_n245), .c(new_n241), .d(new_n244), .o1(new_n246));
  aoai13aa1n02x5               g151(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  nanp02aa1n02x5               g153(.a(new_n228), .b(new_n227), .o1(new_n249));
  xnrc02aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .out0(new_n250));
  xnrc02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .out0(new_n251));
  norp02aa1n02x5               g156(.a(new_n251), .b(new_n250), .o1(new_n252));
  nona23aa1n02x4               g157(.a(new_n197), .b(new_n252), .c(new_n249), .d(new_n218), .out0(new_n253));
  nano22aa1n02x4               g158(.a(new_n249), .b(new_n244), .c(new_n245), .out0(new_n254));
  160nm_ficinv00aa1n08x5       g159(.clk(\a[24] ), .clkout(new_n255));
  160nm_ficinv00aa1n08x5       g160(.clk(\b[23] ), .clkout(new_n256));
  oaoi03aa1n02x5               g161(.a(new_n255), .b(new_n256), .c(new_n243), .o1(new_n257));
  oai013aa1n02x4               g162(.a(new_n257), .b(new_n238), .c(new_n250), .d(new_n251), .o1(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(new_n236), .c(new_n254), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n259), .b(new_n253), .c(new_n181), .d(new_n189), .o1(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  xorc02aa1n02x5               g168(.a(\a[26] ), .b(\b[25] ), .out0(new_n264));
  aoi112aa1n02x5               g169(.a(new_n262), .b(new_n264), .c(new_n260), .d(new_n263), .o1(new_n265));
  aoai13aa1n02x5               g170(.a(new_n264), .b(new_n262), .c(new_n260), .d(new_n263), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n266), .b(new_n265), .out0(\s[26] ));
  nanp02aa1n02x5               g172(.a(new_n155), .b(new_n184), .o1(new_n268));
  nona22aa1n02x4               g173(.a(new_n268), .b(new_n188), .c(new_n185), .out0(new_n269));
  and002aa1n02x5               g174(.a(new_n264), .b(new_n263), .o(new_n270));
  nano32aa1n02x4               g175(.a(new_n220), .b(new_n270), .c(new_n234), .d(new_n252), .out0(new_n271));
  aoai13aa1n02x5               g176(.a(new_n271), .b(new_n269), .c(new_n150), .d(new_n180), .o1(new_n272));
  norp02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .o1(new_n273));
  160nm_ficinv00aa1n08x5       g178(.clk(new_n273), .clkout(new_n274));
  aoi112aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n275));
  160nm_ficinv00aa1n08x5       g180(.clk(new_n275), .clkout(new_n276));
  nanp02aa1n02x5               g181(.a(new_n234), .b(new_n252), .o1(new_n277));
  160nm_ficinv00aa1n08x5       g182(.clk(new_n257), .clkout(new_n278));
  aoi012aa1n02x5               g183(.a(new_n278), .b(new_n252), .c(new_n239), .o1(new_n279));
  160nm_ficinv00aa1n08x5       g184(.clk(new_n270), .clkout(new_n280));
  oaoi13aa1n02x5               g185(.a(new_n280), .b(new_n279), .c(new_n223), .d(new_n277), .o1(new_n281));
  nano22aa1n02x4               g186(.a(new_n281), .b(new_n274), .c(new_n276), .out0(new_n282));
  norp02aa1n02x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  norb02aa1n02x5               g189(.a(new_n284), .b(new_n283), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n282), .c(new_n272), .out0(\s[27] ));
  160nm_ficinv00aa1n08x5       g191(.clk(new_n283), .clkout(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[27] ), .b(\a[28] ), .out0(new_n288));
  aoai13aa1n02x5               g193(.a(new_n270), .b(new_n258), .c(new_n236), .d(new_n254), .o1(new_n289));
  nona22aa1n02x4               g194(.a(new_n289), .b(new_n275), .c(new_n273), .out0(new_n290));
  aoai13aa1n02x5               g195(.a(new_n284), .b(new_n290), .c(new_n190), .d(new_n271), .o1(new_n291));
  aoi012aa1n02x5               g196(.a(new_n288), .b(new_n291), .c(new_n287), .o1(new_n292));
  aobi12aa1n02x5               g197(.a(new_n284), .b(new_n282), .c(new_n272), .out0(new_n293));
  nano22aa1n02x4               g198(.a(new_n293), .b(new_n287), .c(new_n288), .out0(new_n294));
  norp02aa1n02x5               g199(.a(new_n292), .b(new_n294), .o1(\s[28] ));
  nano22aa1n02x4               g200(.a(new_n288), .b(new_n287), .c(new_n284), .out0(new_n296));
  aoai13aa1n02x5               g201(.a(new_n296), .b(new_n290), .c(new_n190), .d(new_n271), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .out0(new_n299));
  aoi012aa1n02x5               g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x5               g205(.a(new_n296), .b(new_n282), .c(new_n272), .out0(new_n301));
  nano22aa1n02x4               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n02x5               g207(.a(new_n300), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g209(.a(new_n285), .b(new_n299), .c(new_n288), .out0(new_n305));
  aoai13aa1n02x5               g210(.a(new_n305), .b(new_n290), .c(new_n190), .d(new_n271), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .out0(new_n308));
  aoi012aa1n02x5               g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  aobi12aa1n02x5               g214(.a(new_n305), .b(new_n282), .c(new_n272), .out0(new_n310));
  nano22aa1n02x4               g215(.a(new_n310), .b(new_n307), .c(new_n308), .out0(new_n311));
  norp02aa1n02x5               g216(.a(new_n309), .b(new_n311), .o1(\s[30] ));
  norb03aa1n02x5               g217(.a(new_n296), .b(new_n308), .c(new_n299), .out0(new_n313));
  aobi12aa1n02x5               g218(.a(new_n313), .b(new_n282), .c(new_n272), .out0(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  nano22aa1n02x4               g221(.a(new_n314), .b(new_n315), .c(new_n316), .out0(new_n317));
  aoai13aa1n02x5               g222(.a(new_n313), .b(new_n290), .c(new_n190), .d(new_n271), .o1(new_n318));
  aoi012aa1n02x5               g223(.a(new_n316), .b(new_n318), .c(new_n315), .o1(new_n319));
  norp02aa1n02x5               g224(.a(new_n319), .b(new_n317), .o1(\s[31] ));
  xnrb03aa1n02x5               g225(.a(new_n107), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g226(.a(\a[3] ), .b(\b[2] ), .c(new_n107), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g228(.a(new_n114), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g229(.a(\a[5] ), .b(\b[4] ), .c(new_n146), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g231(.a(new_n121), .b(new_n120), .out0(new_n327));
  oai112aa1n02x5               g232(.a(new_n327), .b(new_n116), .c(new_n325), .d(new_n115), .o1(new_n328));
  oaoi13aa1n02x5               g233(.a(new_n327), .b(new_n116), .c(new_n325), .d(new_n115), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n328), .b(new_n329), .out0(\s[7] ));
  norb02aa1n02x5               g235(.a(new_n119), .b(new_n118), .out0(new_n331));
  160nm_ficinv00aa1n08x5       g236(.clk(new_n120), .clkout(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n331), .b(new_n328), .c(new_n332), .out0(\s[8] ));
  xorb03aa1n02x5               g238(.a(new_n150), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


