// Benchmark "adder" written by ABC on Wed Jul 17 15:58:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n339, new_n341,
    new_n343, new_n345;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor002aa1n03x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n06x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nand02aa1n10x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  aoi012aa1n12x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nand02aa1d28x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand42aa1n04x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n09x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  aoi012aa1d24x5               g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1n09x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  xnrc02aa1n12x5               g017(.a(\b[5] ), .b(\a[6] ), .out0(new_n113));
  nand02aa1n06x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nanb02aa1n12x5               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  nor002aa1d32x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand22aa1n09x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand02aa1d04x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nor002aa1n20x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n119), .b(new_n118), .c(new_n120), .d(new_n117), .out0(new_n121));
  nor043aa1n06x5               g026(.a(new_n121), .b(new_n116), .c(new_n113), .o1(new_n122));
  inv040aa1d32x5               g027(.a(\a[6] ), .o1(new_n123));
  inv040aa1n16x5               g028(.a(\b[5] ), .o1(new_n124));
  tech160nm_fioaoi03aa1n02p5x5 g029(.a(new_n123), .b(new_n124), .c(new_n115), .o1(new_n125));
  tech160nm_fiaoi012aa1n03p5x5 g030(.a(new_n117), .b(new_n120), .c(new_n118), .o1(new_n126));
  tech160nm_fioai012aa1n05x5   g031(.a(new_n126), .b(new_n121), .c(new_n125), .o1(new_n127));
  nand42aa1n16x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n03x5               g034(.a(new_n129), .b(new_n127), .c(new_n112), .d(new_n122), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  nor002aa1n16x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand02aa1d16x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  nano23aa1n03x7               g039(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n135));
  nanb02aa1n06x5               g040(.a(new_n105), .b(new_n135), .out0(new_n136));
  nano23aa1n06x5               g041(.a(new_n120), .b(new_n117), .c(new_n118), .d(new_n119), .out0(new_n137));
  nona22aa1n02x4               g042(.a(new_n137), .b(new_n113), .c(new_n116), .out0(new_n138));
  oao003aa1n02x5               g043(.a(new_n123), .b(new_n124), .c(new_n115), .carry(new_n139));
  aobi12aa1n06x5               g044(.a(new_n126), .b(new_n137), .c(new_n139), .out0(new_n140));
  aoai13aa1n12x5               g045(.a(new_n140), .b(new_n138), .c(new_n136), .d(new_n111), .o1(new_n141));
  aoai13aa1n03x5               g046(.a(new_n98), .b(new_n100), .c(new_n141), .d(new_n128), .o1(new_n142));
  tech160nm_fioai012aa1n03p5x5 g047(.a(new_n142), .b(\b[9] ), .c(\a[10] ), .o1(new_n143));
  nand42aa1n02x5               g048(.a(new_n130), .b(new_n101), .o1(new_n144));
  oai012aa1n02x5               g049(.a(new_n98), .b(new_n144), .c(new_n97), .o1(new_n145));
  mtn022aa1n02x5               g050(.a(new_n143), .b(new_n145), .sa(new_n134), .o1(\s[11] ));
  nor002aa1n20x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1d28x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n03x5               g055(.a(new_n150), .b(new_n132), .c(new_n143), .d(new_n133), .o1(new_n151));
  aoai13aa1n03x5               g056(.a(new_n134), .b(new_n97), .c(new_n144), .d(new_n98), .o1(new_n152));
  nona22aa1n02x5               g057(.a(new_n152), .b(new_n150), .c(new_n132), .out0(new_n153));
  nanp02aa1n03x5               g058(.a(new_n151), .b(new_n153), .o1(\s[12] ));
  nano23aa1d15x5               g059(.a(new_n97), .b(new_n100), .c(new_n128), .d(new_n98), .out0(new_n155));
  nano23aa1d15x5               g060(.a(new_n132), .b(new_n147), .c(new_n148), .d(new_n133), .out0(new_n156));
  nand22aa1n12x5               g061(.a(new_n156), .b(new_n155), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n127), .c(new_n112), .d(new_n122), .o1(new_n159));
  nanb03aa1n09x5               g064(.a(new_n147), .b(new_n148), .c(new_n133), .out0(new_n160));
  oai122aa1n12x5               g065(.a(new_n98), .b(new_n97), .c(new_n100), .d(\b[10] ), .e(\a[11] ), .o1(new_n161));
  aoi012aa1d18x5               g066(.a(new_n147), .b(new_n132), .c(new_n148), .o1(new_n162));
  oai012aa1d24x5               g067(.a(new_n162), .b(new_n161), .c(new_n160), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  nor002aa1d32x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nanp02aa1n09x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n159), .c(new_n164), .out0(\s[13] ));
  nanp02aa1n02x5               g073(.a(new_n159), .b(new_n164), .o1(new_n169));
  aoi012aa1n02x5               g074(.a(new_n165), .b(new_n169), .c(new_n166), .o1(new_n170));
  xnrb03aa1n03x5               g075(.a(new_n170), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nand02aa1n06x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nano23aa1n03x7               g078(.a(new_n165), .b(new_n172), .c(new_n173), .d(new_n166), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n163), .c(new_n141), .d(new_n158), .o1(new_n175));
  tech160nm_fioai012aa1n05x5   g080(.a(new_n173), .b(new_n172), .c(new_n165), .o1(new_n176));
  nor042aa1d18x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand02aa1d28x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  norb02aa1n03x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n175), .c(new_n176), .out0(\s[15] ));
  nona23aa1n03x5               g085(.a(new_n173), .b(new_n166), .c(new_n165), .d(new_n172), .out0(new_n181));
  aoai13aa1n02x7               g086(.a(new_n176), .b(new_n181), .c(new_n159), .d(new_n164), .o1(new_n182));
  nor002aa1d32x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nand02aa1d08x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n183), .b(new_n184), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n177), .c(new_n182), .d(new_n178), .o1(new_n186));
  aoi112aa1n03x4               g091(.a(new_n177), .b(new_n185), .c(new_n182), .d(new_n178), .o1(new_n187));
  nanb02aa1n03x5               g092(.a(new_n187), .b(new_n186), .out0(\s[16] ));
  nano23aa1n03x7               g093(.a(new_n177), .b(new_n183), .c(new_n184), .d(new_n178), .out0(new_n189));
  nano22aa1d15x5               g094(.a(new_n157), .b(new_n174), .c(new_n189), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n127), .c(new_n112), .d(new_n122), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n183), .o1(new_n192));
  nano32aa1n06x5               g097(.a(new_n181), .b(new_n184), .c(new_n179), .d(new_n192), .out0(new_n193));
  nanb03aa1n03x5               g098(.a(new_n183), .b(new_n184), .c(new_n178), .out0(new_n194));
  tech160nm_fiaoi012aa1n02p5x5 g099(.a(new_n183), .b(new_n177), .c(new_n184), .o1(new_n195));
  oai013aa1n06x5               g100(.a(new_n195), .b(new_n194), .c(new_n176), .d(new_n177), .o1(new_n196));
  aoi012aa1d24x5               g101(.a(new_n196), .b(new_n163), .c(new_n193), .o1(new_n197));
  nand02aa1d08x5               g102(.a(new_n191), .b(new_n197), .o1(new_n198));
  xorc02aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  aoi112aa1n02x5               g104(.a(new_n199), .b(new_n196), .c(new_n163), .d(new_n193), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n198), .b(new_n199), .c(new_n191), .d(new_n200), .o1(\s[17] ));
  inv000aa1d42x5               g106(.a(\a[18] ), .o1(new_n202));
  nor002aa1n04x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  tech160nm_fiaoi012aa1n05x5   g108(.a(new_n203), .b(new_n198), .c(new_n199), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[17] ), .c(new_n202), .out0(\s[18] ));
  nand02aa1d06x5               g110(.a(new_n163), .b(new_n193), .o1(new_n206));
  nanb02aa1n12x5               g111(.a(new_n196), .b(new_n206), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  nor042aa1n02x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nanp02aa1n12x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nano23aa1n06x5               g115(.a(new_n203), .b(new_n209), .c(new_n210), .d(new_n208), .out0(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n207), .c(new_n141), .d(new_n190), .o1(new_n212));
  oa0012aa1n06x5               g117(.a(new_n210), .b(new_n209), .c(new_n203), .o(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nor042aa1n06x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand02aa1n08x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n09x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n03p5x5 g124(.a(new_n212), .b(new_n214), .o1(new_n220));
  nor042aa1d18x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1d12x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanb02aa1n02x5               g127(.a(new_n221), .b(new_n222), .out0(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n215), .c(new_n220), .d(new_n216), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n217), .b(new_n213), .c(new_n198), .d(new_n211), .o1(new_n225));
  nona22aa1n02x5               g130(.a(new_n225), .b(new_n223), .c(new_n215), .out0(new_n226));
  nanp02aa1n03x5               g131(.a(new_n224), .b(new_n226), .o1(\s[20] ));
  nano22aa1n03x7               g132(.a(new_n223), .b(new_n211), .c(new_n217), .out0(new_n228));
  inv030aa1n02x5               g133(.a(new_n228), .o1(new_n229));
  nanb03aa1d24x5               g134(.a(new_n221), .b(new_n222), .c(new_n216), .out0(new_n230));
  oai022aa1d24x5               g135(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n231));
  inv040aa1d30x5               g136(.a(\b[18] ), .o1(new_n232));
  nanb02aa1n12x5               g137(.a(\a[19] ), .b(new_n232), .out0(new_n233));
  nanp03aa1d12x5               g138(.a(new_n231), .b(new_n233), .c(new_n210), .o1(new_n234));
  aoi012aa1d24x5               g139(.a(new_n221), .b(new_n215), .c(new_n222), .o1(new_n235));
  oai012aa1d24x5               g140(.a(new_n235), .b(new_n234), .c(new_n230), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n237), .b(new_n229), .c(new_n191), .d(new_n197), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[20] ), .b(\a[21] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(new_n240), .b(new_n236), .c(new_n198), .d(new_n228), .o1(new_n241));
  aoi012aa1n02x5               g146(.a(new_n241), .b(new_n238), .c(new_n240), .o1(\s[21] ));
  nor002aa1n02x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[21] ), .b(\a[22] ), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n243), .c(new_n238), .d(new_n240), .o1(new_n245));
  aoi112aa1n03x4               g150(.a(new_n243), .b(new_n244), .c(new_n238), .d(new_n240), .o1(new_n246));
  nanb02aa1n03x5               g151(.a(new_n246), .b(new_n245), .out0(\s[22] ));
  nona32aa1n03x5               g152(.a(new_n198), .b(new_n244), .c(new_n239), .d(new_n229), .out0(new_n248));
  nor042aa1n06x5               g153(.a(new_n244), .b(new_n239), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\a[22] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[21] ), .o1(new_n251));
  oao003aa1n06x5               g156(.a(new_n250), .b(new_n251), .c(new_n243), .carry(new_n252));
  aoi012aa1n02x7               g157(.a(new_n252), .b(new_n236), .c(new_n249), .o1(new_n253));
  xorc02aa1n12x5               g158(.a(\a[23] ), .b(\b[22] ), .out0(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n248), .c(new_n253), .out0(\s[23] ));
  nand42aa1n02x5               g160(.a(new_n228), .b(new_n249), .o1(new_n256));
  aoai13aa1n04x5               g161(.a(new_n253), .b(new_n256), .c(new_n191), .d(new_n197), .o1(new_n257));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[23] ), .b(\a[24] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n258), .c(new_n257), .d(new_n254), .o1(new_n260));
  aoi112aa1n03x4               g165(.a(new_n258), .b(new_n259), .c(new_n257), .d(new_n254), .o1(new_n261));
  nanb02aa1n03x5               g166(.a(new_n261), .b(new_n260), .out0(\s[24] ));
  norb02aa1n03x5               g167(.a(new_n254), .b(new_n259), .out0(new_n263));
  nano22aa1n03x7               g168(.a(new_n229), .b(new_n249), .c(new_n263), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n207), .c(new_n141), .d(new_n190), .o1(new_n265));
  nano22aa1n02x4               g170(.a(new_n221), .b(new_n216), .c(new_n222), .out0(new_n266));
  oai012aa1n02x5               g171(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .o1(new_n267));
  oab012aa1n04x5               g172(.a(new_n267), .b(new_n203), .c(new_n209), .out0(new_n268));
  inv000aa1n02x5               g173(.a(new_n235), .o1(new_n269));
  aoai13aa1n06x5               g174(.a(new_n249), .b(new_n269), .c(new_n268), .d(new_n266), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n252), .o1(new_n271));
  nanb02aa1n02x5               g176(.a(new_n259), .b(new_n254), .out0(new_n272));
  aoi112aa1n02x5               g177(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n273));
  oab012aa1n02x4               g178(.a(new_n273), .b(\a[24] ), .c(\b[23] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .d(new_n271), .o1(new_n275));
  nanb02aa1n06x5               g180(.a(new_n275), .b(new_n265), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  aoai13aa1n04x5               g182(.a(new_n263), .b(new_n252), .c(new_n236), .d(new_n249), .o1(new_n278));
  nano22aa1n02x4               g183(.a(new_n277), .b(new_n278), .c(new_n274), .out0(new_n279));
  aoi022aa1n02x5               g184(.a(new_n276), .b(new_n277), .c(new_n265), .d(new_n279), .o1(\s[25] ));
  norp02aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .o1(new_n281));
  xnrc02aa1n12x5               g186(.a(\b[25] ), .b(\a[26] ), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n276), .d(new_n277), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n277), .b(new_n275), .c(new_n198), .d(new_n264), .o1(new_n284));
  nona22aa1n02x5               g189(.a(new_n284), .b(new_n282), .c(new_n281), .out0(new_n285));
  nanp02aa1n03x5               g190(.a(new_n283), .b(new_n285), .o1(\s[26] ));
  nanb02aa1n02x5               g191(.a(new_n282), .b(new_n277), .out0(new_n287));
  inv030aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nano32aa1n03x7               g193(.a(new_n229), .b(new_n288), .c(new_n249), .d(new_n263), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n207), .c(new_n141), .d(new_n190), .o1(new_n290));
  aoi112aa1n02x5               g195(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n291));
  oab012aa1n02x4               g196(.a(new_n291), .b(\a[26] ), .c(\b[25] ), .out0(new_n292));
  aobi12aa1n06x5               g197(.a(new_n292), .b(new_n275), .c(new_n288), .out0(new_n293));
  tech160nm_fixorc02aa1n03p5x5 g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(new_n290), .out0(\s[27] ));
  nand42aa1n02x5               g200(.a(new_n293), .b(new_n290), .o1(new_n296));
  norp02aa1n02x5               g201(.a(\b[26] ), .b(\a[27] ), .o1(new_n297));
  norp02aa1n02x5               g202(.a(\b[27] ), .b(\a[28] ), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(\b[27] ), .b(\a[28] ), .o1(new_n299));
  nanb02aa1n02x5               g204(.a(new_n298), .b(new_n299), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n297), .c(new_n296), .d(new_n294), .o1(new_n301));
  inv000aa1n02x5               g206(.a(new_n249), .o1(new_n302));
  nona23aa1n02x4               g207(.a(new_n228), .b(new_n288), .c(new_n302), .d(new_n272), .out0(new_n303));
  aoi012aa1n06x5               g208(.a(new_n303), .b(new_n191), .c(new_n197), .o1(new_n304));
  aoai13aa1n04x5               g209(.a(new_n292), .b(new_n287), .c(new_n278), .d(new_n274), .o1(new_n305));
  oaih12aa1n02x5               g210(.a(new_n294), .b(new_n305), .c(new_n304), .o1(new_n306));
  nona22aa1n02x5               g211(.a(new_n306), .b(new_n300), .c(new_n297), .out0(new_n307));
  nanp02aa1n03x5               g212(.a(new_n301), .b(new_n307), .o1(\s[28] ));
  xnrc02aa1n02x5               g213(.a(\b[28] ), .b(\a[29] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n294), .b(new_n300), .out0(new_n310));
  oaih12aa1n02x5               g215(.a(new_n310), .b(new_n305), .c(new_n304), .o1(new_n311));
  oai012aa1n02x5               g216(.a(new_n299), .b(new_n298), .c(new_n297), .o1(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n309), .b(new_n311), .c(new_n312), .o1(new_n313));
  inv000aa1n02x5               g218(.a(new_n310), .o1(new_n314));
  aoi012aa1n02x7               g219(.a(new_n314), .b(new_n293), .c(new_n290), .o1(new_n315));
  nano22aa1n02x4               g220(.a(new_n315), .b(new_n309), .c(new_n312), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n313), .b(new_n316), .o1(\s[29] ));
  xorb03aa1n02x5               g222(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g223(.a(new_n294), .b(new_n309), .c(new_n300), .out0(new_n319));
  oaih12aa1n02x5               g224(.a(new_n319), .b(new_n305), .c(new_n304), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .carry(new_n321));
  tech160nm_finand02aa1n03p5x5 g226(.a(new_n320), .b(new_n321), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  norb02aa1n02x5               g228(.a(new_n321), .b(new_n323), .out0(new_n324));
  aoi022aa1n02x7               g229(.a(new_n322), .b(new_n323), .c(new_n320), .d(new_n324), .o1(\s[30] ));
  nona23aa1n02x4               g230(.a(new_n294), .b(new_n323), .c(new_n309), .d(new_n300), .out0(new_n326));
  oabi12aa1n03x5               g231(.a(new_n326), .b(new_n305), .c(new_n304), .out0(new_n327));
  xorc02aa1n02x5               g232(.a(\a[31] ), .b(\b[30] ), .out0(new_n328));
  and002aa1n02x5               g233(.a(\b[29] ), .b(\a[30] ), .o(new_n329));
  oabi12aa1n02x5               g234(.a(new_n328), .b(\a[30] ), .c(\b[29] ), .out0(new_n330));
  oab012aa1n02x4               g235(.a(new_n330), .b(new_n321), .c(new_n329), .out0(new_n331));
  oao003aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n326), .c(new_n293), .d(new_n290), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n333), .b(new_n328), .c(new_n327), .d(new_n331), .o1(\s[31] ));
  xnrb03aa1n02x5               g239(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g240(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xobna2aa1n03x5               g242(.a(new_n116), .b(new_n136), .c(new_n111), .out0(\s[5] ));
  tech160nm_fiao0012aa1n03p5x5 g243(.a(new_n115), .b(new_n112), .c(new_n114), .o(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fioaoi03aa1n03p5x5 g245(.a(new_n123), .b(new_n124), .c(new_n339), .o1(new_n341));
  xnrb03aa1n02x5               g246(.a(new_n341), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n03x5               g247(.a(\a[7] ), .b(\b[6] ), .c(new_n341), .o1(new_n343));
  xorb03aa1n02x5               g248(.a(new_n343), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  aoi112aa1n02x5               g249(.a(new_n129), .b(new_n127), .c(new_n112), .d(new_n122), .o1(new_n345));
  aoi012aa1n02x5               g250(.a(new_n345), .b(new_n141), .c(new_n129), .o1(\s[9] ));
endmodule


