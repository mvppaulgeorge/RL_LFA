// Benchmark "adder" written by ABC on Thu Jul 18 03:11:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n330, new_n333,
    new_n334, new_n336, new_n337, new_n338, new_n340;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[1] ), .o1(new_n102));
  inv040aa1d32x5               g007(.a(\b[0] ), .o1(new_n103));
  norp02aa1n04x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand02aa1n03x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  oaoi13aa1n09x5               g010(.a(new_n104), .b(new_n105), .c(new_n102), .d(new_n103), .o1(new_n106));
  nand02aa1n08x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanp02aa1n09x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nona23aa1n09x5               g015(.a(new_n107), .b(new_n110), .c(new_n109), .d(new_n108), .out0(new_n111));
  tech160nm_fiaoi012aa1n05x5   g016(.a(new_n108), .b(new_n109), .c(new_n107), .o1(new_n112));
  oai012aa1n12x5               g017(.a(new_n112), .b(new_n111), .c(new_n106), .o1(new_n113));
  orn002aa1n03x5               g018(.a(\a[6] ), .b(\b[5] ), .o(new_n114));
  tech160nm_finand02aa1n05x5   g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand02aa1n04x5               g020(.a(new_n114), .b(new_n115), .o1(new_n116));
  nor022aa1n08x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand22aa1n09x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1n06x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nor022aa1n08x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n119), .b(new_n118), .c(new_n120), .d(new_n117), .out0(new_n121));
  tech160nm_fixnrc02aa1n04x5   g026(.a(\b[4] ), .b(\a[5] ), .out0(new_n122));
  nor043aa1n06x5               g027(.a(new_n121), .b(new_n122), .c(new_n116), .o1(new_n123));
  oai022aa1d24x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  nand42aa1n06x5               g029(.a(new_n124), .b(new_n115), .o1(new_n125));
  tech160nm_fiao0012aa1n02p5x5 g030(.a(new_n117), .b(new_n120), .c(new_n118), .o(new_n126));
  oabi12aa1n06x5               g031(.a(new_n126), .b(new_n121), .c(new_n125), .out0(new_n127));
  nand42aa1n16x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n03x5               g034(.a(new_n129), .b(new_n127), .c(new_n113), .d(new_n123), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  norp02aa1n02x5               g036(.a(new_n100), .b(new_n97), .o1(new_n132));
  aoi022aa1n03x5               g037(.a(new_n130), .b(new_n132), .c(\b[9] ), .d(\a[10] ), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv040aa1d32x5               g039(.a(\a[12] ), .o1(new_n135));
  inv040aa1d28x5               g040(.a(\b[11] ), .o1(new_n136));
  nand42aa1n04x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  nanp02aa1n04x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  inv040aa1d32x5               g043(.a(\a[11] ), .o1(new_n139));
  inv040aa1d32x5               g044(.a(\b[10] ), .o1(new_n140));
  oaoi03aa1n03x5               g045(.a(new_n139), .b(new_n140), .c(new_n133), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n137), .c(new_n138), .out0(\s[12] ));
  nanp02aa1n03x5               g047(.a(new_n113), .b(new_n123), .o1(new_n143));
  nano23aa1n02x5               g048(.a(new_n120), .b(new_n117), .c(new_n118), .d(new_n119), .out0(new_n144));
  inv000aa1n02x5               g049(.a(new_n125), .o1(new_n145));
  tech160nm_fiaoi012aa1n04x5   g050(.a(new_n126), .b(new_n144), .c(new_n145), .o1(new_n146));
  nand42aa1n06x5               g051(.a(new_n140), .b(new_n139), .o1(new_n147));
  nand42aa1n03x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n137), .b(new_n138), .o1(new_n150));
  nano23aa1n09x5               g055(.a(new_n97), .b(new_n100), .c(new_n128), .d(new_n98), .out0(new_n151));
  nona22aa1n12x5               g056(.a(new_n151), .b(new_n150), .c(new_n149), .out0(new_n152));
  tech160nm_fioai012aa1n05x5   g057(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(new_n153), .b(new_n147), .o1(new_n154));
  aoi022aa1d18x5               g059(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n155));
  aoi022aa1n02x5               g060(.a(new_n154), .b(new_n155), .c(new_n136), .d(new_n135), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n152), .c(new_n143), .d(new_n146), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1d28x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand42aa1n16x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1d15x5               g069(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n165));
  oa0012aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n159), .o(new_n166));
  nor042aa1d18x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nand22aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nanb02aa1d36x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n04x5               g075(.a(new_n170), .b(new_n166), .c(new_n157), .d(new_n165), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n170), .b(new_n166), .c(new_n157), .d(new_n165), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[15] ));
  nor042aa1n04x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1n08x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanb02aa1n06x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  oai112aa1n02x5               g081(.a(new_n171), .b(new_n176), .c(\b[14] ), .d(\a[15] ), .o1(new_n177));
  oaoi13aa1n02x5               g082(.a(new_n176), .b(new_n171), .c(\a[15] ), .d(\b[14] ), .o1(new_n178));
  norb02aa1n02x7               g083(.a(new_n177), .b(new_n178), .out0(\s[16] ));
  nona22aa1n09x5               g084(.a(new_n165), .b(new_n169), .c(new_n176), .out0(new_n180));
  nor042aa1n09x5               g085(.a(new_n180), .b(new_n152), .o1(new_n181));
  aoai13aa1n12x5               g086(.a(new_n181), .b(new_n127), .c(new_n113), .d(new_n123), .o1(new_n182));
  inv000aa1n02x5               g087(.a(new_n155), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n137), .b(new_n183), .c(new_n153), .d(new_n147), .o1(new_n184));
  oai112aa1n02x5               g089(.a(new_n164), .b(new_n168), .c(new_n163), .d(new_n159), .o1(new_n185));
  nona22aa1n03x5               g090(.a(new_n185), .b(new_n174), .c(new_n167), .out0(new_n186));
  aboi22aa1n12x5               g091(.a(new_n180), .b(new_n184), .c(new_n186), .d(new_n175), .out0(new_n187));
  nor042aa1n12x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  nanp02aa1n04x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  norb02aa1n15x5               g094(.a(new_n189), .b(new_n188), .out0(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n190), .b(new_n182), .c(new_n187), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(new_n188), .o1(new_n192));
  and002aa1n02x5               g097(.a(\b[0] ), .b(\a[1] ), .o(new_n193));
  oaoi03aa1n02x5               g098(.a(\a[2] ), .b(\b[1] ), .c(new_n193), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n107), .b(new_n108), .out0(new_n195));
  norb02aa1n02x7               g100(.a(new_n110), .b(new_n109), .out0(new_n196));
  nanp03aa1n02x5               g101(.a(new_n194), .b(new_n195), .c(new_n196), .o1(new_n197));
  nona22aa1n02x4               g102(.a(new_n144), .b(new_n122), .c(new_n116), .out0(new_n198));
  aoai13aa1n06x5               g103(.a(new_n146), .b(new_n198), .c(new_n197), .d(new_n112), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(new_n186), .b(new_n175), .o1(new_n200));
  oai012aa1n02x5               g105(.a(new_n200), .b(new_n156), .c(new_n180), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n190), .b(new_n201), .c(new_n199), .d(new_n181), .o1(new_n202));
  xnrc02aa1n12x5               g107(.a(\b[17] ), .b(\a[18] ), .out0(new_n203));
  xobna2aa1n03x5               g108(.a(new_n203), .b(new_n202), .c(new_n192), .out0(\s[18] ));
  nanp02aa1n06x5               g109(.a(new_n182), .b(new_n187), .o1(new_n205));
  nano22aa1n02x4               g110(.a(new_n203), .b(new_n192), .c(new_n189), .out0(new_n206));
  oaoi03aa1n02x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n207));
  nor002aa1d32x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nand42aa1d28x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nanb02aa1d24x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n207), .c(new_n205), .d(new_n206), .o1(new_n212));
  aoi112aa1n02x5               g117(.a(new_n211), .b(new_n207), .c(new_n205), .d(new_n206), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n212), .b(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand02aa1d28x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1d27x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  nona22aa1n06x5               g123(.a(new_n212), .b(new_n218), .c(new_n208), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n208), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n218), .o1(new_n221));
  tech160nm_fiaoi012aa1n05x5   g126(.a(new_n221), .b(new_n212), .c(new_n220), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n219), .b(new_n222), .out0(\s[20] ));
  nano23aa1d15x5               g128(.a(new_n210), .b(new_n203), .c(new_n190), .d(new_n218), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  nand02aa1n10x5               g130(.a(\b[17] ), .b(\a[18] ), .o1(new_n226));
  nanb03aa1d24x5               g131(.a(new_n208), .b(new_n209), .c(new_n226), .out0(new_n227));
  oai022aa1d24x5               g132(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n228));
  inv020aa1n02x5               g133(.a(new_n216), .o1(new_n229));
  nand23aa1n03x5               g134(.a(new_n228), .b(new_n229), .c(new_n217), .o1(new_n230));
  aoi012aa1n06x5               g135(.a(new_n216), .b(new_n208), .c(new_n217), .o1(new_n231));
  oai012aa1n12x5               g136(.a(new_n231), .b(new_n230), .c(new_n227), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n225), .c(new_n182), .d(new_n187), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  xorc02aa1n12x5               g141(.a(\a[21] ), .b(\b[20] ), .out0(new_n237));
  xorc02aa1n12x5               g142(.a(\a[22] ), .b(\b[21] ), .out0(new_n238));
  aoi112aa1n03x5               g143(.a(new_n236), .b(new_n238), .c(new_n234), .d(new_n237), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n238), .b(new_n236), .c(new_n234), .d(new_n237), .o1(new_n240));
  norb02aa1n02x7               g145(.a(new_n240), .b(new_n239), .out0(\s[22] ));
  inv000aa1d42x5               g146(.a(\a[21] ), .o1(new_n242));
  inv000aa1d42x5               g147(.a(\a[22] ), .o1(new_n243));
  xroi22aa1d04x5               g148(.a(new_n242), .b(\b[20] ), .c(new_n243), .d(\b[21] ), .out0(new_n244));
  nona23aa1n02x4               g149(.a(new_n244), .b(new_n206), .c(new_n210), .d(new_n221), .out0(new_n245));
  nano22aa1d15x5               g150(.a(new_n208), .b(new_n226), .c(new_n209), .out0(new_n246));
  nanp03aa1d12x5               g151(.a(new_n246), .b(new_n228), .c(new_n218), .o1(new_n247));
  nand22aa1n04x5               g152(.a(new_n238), .b(new_n237), .o1(new_n248));
  inv040aa1d28x5               g153(.a(\b[21] ), .o1(new_n249));
  oaoi03aa1n12x5               g154(.a(new_n243), .b(new_n249), .c(new_n236), .o1(new_n250));
  aoai13aa1n12x5               g155(.a(new_n250), .b(new_n248), .c(new_n247), .d(new_n231), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n245), .c(new_n182), .d(new_n187), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  xorc02aa1n12x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  aoi112aa1n03x5               g162(.a(new_n255), .b(new_n257), .c(new_n253), .d(new_n256), .o1(new_n258));
  aoai13aa1n03x5               g163(.a(new_n257), .b(new_n255), .c(new_n253), .d(new_n256), .o1(new_n259));
  norb02aa1n02x7               g164(.a(new_n259), .b(new_n258), .out0(\s[24] ));
  nand02aa1n02x5               g165(.a(new_n257), .b(new_n256), .o1(new_n261));
  nona22aa1n02x4               g166(.a(new_n224), .b(new_n248), .c(new_n261), .out0(new_n262));
  inv030aa1n02x5               g167(.a(new_n261), .o1(new_n263));
  inv000aa1d42x5               g168(.a(\a[24] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(\b[23] ), .o1(new_n265));
  oaoi03aa1n12x5               g170(.a(new_n264), .b(new_n265), .c(new_n255), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  tech160nm_fiaoi012aa1n05x5   g172(.a(new_n267), .b(new_n251), .c(new_n263), .o1(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n262), .c(new_n182), .d(new_n187), .o1(new_n269));
  xorb03aa1n02x5               g174(.a(new_n269), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xorc02aa1n12x5               g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  aoi112aa1n03x5               g178(.a(new_n271), .b(new_n273), .c(new_n269), .d(new_n272), .o1(new_n274));
  aoai13aa1n04x5               g179(.a(new_n273), .b(new_n271), .c(new_n269), .d(new_n272), .o1(new_n275));
  norb02aa1n03x4               g180(.a(new_n275), .b(new_n274), .out0(\s[26] ));
  nand42aa1n02x5               g181(.a(new_n273), .b(new_n272), .o1(new_n277));
  inv000aa1n04x5               g182(.a(new_n277), .o1(new_n278));
  nona23aa1d18x5               g183(.a(new_n224), .b(new_n278), .c(new_n261), .d(new_n248), .out0(new_n279));
  inv040aa1n06x5               g184(.a(new_n279), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n201), .c(new_n199), .d(new_n181), .o1(new_n281));
  aoai13aa1n12x5               g186(.a(new_n278), .b(new_n267), .c(new_n251), .d(new_n263), .o1(new_n282));
  aoi112aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n283));
  oab012aa1n09x5               g188(.a(new_n283), .b(\a[26] ), .c(\b[25] ), .out0(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  aoi013aa1n06x4               g191(.a(new_n286), .b(new_n281), .c(new_n282), .d(new_n284), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n250), .o1(new_n288));
  aoai13aa1n04x5               g193(.a(new_n263), .b(new_n288), .c(new_n232), .d(new_n244), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n284), .b(new_n277), .c(new_n289), .d(new_n266), .o1(new_n290));
  aoi112aa1n02x5               g195(.a(new_n290), .b(new_n285), .c(new_n205), .d(new_n280), .o1(new_n291));
  norp02aa1n02x5               g196(.a(new_n287), .b(new_n291), .o1(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  inv040aa1n03x5               g198(.a(new_n293), .o1(new_n294));
  tech160nm_fixnrc02aa1n04x5   g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  nano22aa1n03x7               g200(.a(new_n287), .b(new_n294), .c(new_n295), .out0(new_n296));
  aoi012aa1n06x5               g201(.a(new_n279), .b(new_n182), .c(new_n187), .o1(new_n297));
  oaih12aa1n02x5               g202(.a(new_n285), .b(new_n290), .c(new_n297), .o1(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n295), .b(new_n298), .c(new_n294), .o1(new_n299));
  norp02aa1n03x5               g204(.a(new_n299), .b(new_n296), .o1(\s[28] ));
  xnrc02aa1n02x5               g205(.a(\b[28] ), .b(\a[29] ), .out0(new_n301));
  norb02aa1n12x5               g206(.a(new_n285), .b(new_n295), .out0(new_n302));
  oai012aa1n03x5               g207(.a(new_n302), .b(new_n290), .c(new_n297), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n294), .carry(new_n304));
  tech160nm_fiaoi012aa1n02p5x5 g209(.a(new_n301), .b(new_n303), .c(new_n304), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n302), .o1(new_n306));
  aoi013aa1n02x5               g211(.a(new_n306), .b(new_n281), .c(new_n282), .d(new_n284), .o1(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n301), .c(new_n304), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n305), .b(new_n308), .o1(\s[29] ));
  xnrb03aa1n02x5               g214(.a(new_n193), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n09x5               g215(.a(new_n285), .b(new_n301), .c(new_n295), .out0(new_n311));
  oaih12aa1n02x5               g216(.a(new_n311), .b(new_n290), .c(new_n297), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[29] ), .b(\a[30] ), .out0(new_n314));
  tech160nm_fiaoi012aa1n02p5x5 g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  aoi013aa1n02x5               g221(.a(new_n316), .b(new_n281), .c(new_n282), .d(new_n284), .o1(new_n317));
  nano22aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n314), .out0(new_n318));
  norp02aa1n03x5               g223(.a(new_n315), .b(new_n318), .o1(\s[30] ));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  norb02aa1n03x5               g225(.a(new_n311), .b(new_n314), .out0(new_n321));
  inv000aa1n03x5               g226(.a(new_n321), .o1(new_n322));
  aoi013aa1n02x5               g227(.a(new_n322), .b(new_n281), .c(new_n282), .d(new_n284), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n324));
  nano22aa1n03x5               g229(.a(new_n323), .b(new_n320), .c(new_n324), .out0(new_n325));
  tech160nm_fioai012aa1n05x5   g230(.a(new_n321), .b(new_n290), .c(new_n297), .o1(new_n326));
  aoi012aa1n03x5               g231(.a(new_n320), .b(new_n326), .c(new_n324), .o1(new_n327));
  norp02aa1n03x5               g232(.a(new_n327), .b(new_n325), .o1(\s[31] ));
  xnrc02aa1n02x5               g233(.a(new_n106), .b(new_n196), .out0(\s[3] ));
  aoi112aa1n02x5               g234(.a(new_n109), .b(new_n195), .c(new_n194), .d(new_n196), .o1(new_n330));
  aoib12aa1n02x5               g235(.a(new_n330), .b(new_n113), .c(new_n108), .out0(\s[4] ));
  xorb03aa1n02x5               g236(.a(new_n113), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  orn002aa1n02x5               g237(.a(\a[5] ), .b(\b[4] ), .o(new_n333));
  nanb02aa1n02x5               g238(.a(new_n122), .b(new_n113), .out0(new_n334));
  xobna2aa1n03x5               g239(.a(new_n116), .b(new_n334), .c(new_n333), .out0(\s[6] ));
  nanb02aa1n02x5               g240(.a(new_n120), .b(new_n119), .out0(new_n336));
  norp02aa1n02x5               g241(.a(\b[4] ), .b(\a[5] ), .o1(new_n337));
  nona22aa1n02x4               g242(.a(new_n334), .b(new_n337), .c(new_n116), .out0(new_n338));
  xnbna2aa1n03x5               g243(.a(new_n336), .b(new_n338), .c(new_n115), .out0(\s[7] ));
  aoi013aa1n02x4               g244(.a(new_n120), .b(new_n338), .c(new_n115), .d(new_n119), .o1(new_n340));
  xnrb03aa1n02x5               g245(.a(new_n340), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g246(.a(new_n199), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


