// Benchmark "adder" written by ABC on Thu Jul 18 02:03:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n335, new_n337, new_n340,
    new_n341, new_n342, new_n344, new_n345, new_n346, new_n348, new_n349,
    new_n350, new_n351;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1d28x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  oai012aa1n06x5               g004(.a(new_n99), .b(\b[3] ), .c(\a[4] ), .o1(new_n100));
  nand42aa1n03x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nand42aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor042aa1n09x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nano23aa1n02x5               g008(.a(new_n100), .b(new_n103), .c(new_n101), .d(new_n102), .out0(new_n104));
  nanp02aa1n24x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nor042aa1n06x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nona22aa1n09x5               g011(.a(new_n99), .b(new_n106), .c(new_n105), .out0(new_n107));
  inv000aa1d42x5               g012(.a(\a[4] ), .o1(new_n108));
  inv040aa1d32x5               g013(.a(\b[3] ), .o1(new_n109));
  oao003aa1n03x5               g014(.a(new_n108), .b(new_n109), .c(new_n103), .carry(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .out0(new_n111));
  tech160nm_fixnrc02aa1n02p5x5 g016(.a(\b[4] ), .b(\a[5] ), .out0(new_n112));
  nor002aa1n10x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1d28x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1n12x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand02aa1n12x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n03x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nor043aa1n02x5               g022(.a(new_n117), .b(new_n112), .c(new_n111), .o1(new_n118));
  aoai13aa1n04x5               g023(.a(new_n118), .b(new_n110), .c(new_n104), .d(new_n107), .o1(new_n119));
  nano23aa1n09x5               g024(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n120));
  inv040aa1d32x5               g025(.a(\a[5] ), .o1(new_n121));
  inv040aa1n16x5               g026(.a(\b[4] ), .o1(new_n122));
  nanp02aa1n04x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  oaoi03aa1n12x5               g028(.a(\a[6] ), .b(\b[5] ), .c(new_n123), .o1(new_n124));
  oai022aa1n03x5               g029(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n125));
  aoi022aa1n12x5               g030(.a(new_n120), .b(new_n124), .c(new_n114), .d(new_n125), .o1(new_n126));
  xnrc02aa1n12x5               g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n98), .b(new_n127), .c(new_n119), .d(new_n126), .o1(new_n128));
  nor002aa1d24x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1n16x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n15x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  inv030aa1n02x5               g036(.a(new_n100), .o1(new_n132));
  nano22aa1n03x7               g037(.a(new_n103), .b(new_n101), .c(new_n102), .out0(new_n133));
  nanp03aa1n04x5               g038(.a(new_n133), .b(new_n107), .c(new_n132), .o1(new_n134));
  inv040aa1n02x5               g039(.a(new_n110), .o1(new_n135));
  tech160nm_fixorc02aa1n03p5x5 g040(.a(\a[6] ), .b(\b[5] ), .out0(new_n136));
  tech160nm_fixorc02aa1n04x5   g041(.a(\a[5] ), .b(\b[4] ), .out0(new_n137));
  nand03aa1n03x5               g042(.a(new_n120), .b(new_n136), .c(new_n137), .o1(new_n138));
  aoai13aa1n12x5               g043(.a(new_n126), .b(new_n138), .c(new_n134), .d(new_n135), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n127), .o1(new_n140));
  aoi112aa1n02x5               g045(.a(new_n131), .b(new_n97), .c(new_n139), .d(new_n140), .o1(new_n141));
  aoi012aa1n02x5               g046(.a(new_n141), .b(new_n128), .c(new_n131), .o1(\s[10] ));
  inv000aa1d42x5               g047(.a(new_n129), .o1(new_n143));
  aoai13aa1n06x5               g048(.a(new_n131), .b(new_n97), .c(new_n139), .d(new_n140), .o1(new_n144));
  xorc02aa1n12x5               g049(.a(\a[11] ), .b(\b[10] ), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n144), .c(new_n143), .out0(\s[11] ));
  aoai13aa1n02x5               g051(.a(new_n145), .b(new_n129), .c(new_n128), .d(new_n130), .o1(new_n147));
  xorc02aa1n12x5               g052(.a(\a[12] ), .b(\b[11] ), .out0(new_n148));
  nor042aa1d18x5               g053(.a(\b[10] ), .b(\a[11] ), .o1(new_n149));
  norp02aa1n02x5               g054(.a(new_n148), .b(new_n149), .o1(new_n150));
  inv000aa1n06x5               g055(.a(new_n149), .o1(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[10] ), .b(\a[11] ), .out0(new_n152));
  aoai13aa1n03x5               g057(.a(new_n151), .b(new_n152), .c(new_n144), .d(new_n143), .o1(new_n153));
  aoi022aa1n03x5               g058(.a(new_n153), .b(new_n148), .c(new_n147), .d(new_n150), .o1(\s[12] ));
  nona23aa1n09x5               g059(.a(new_n148), .b(new_n131), .c(new_n127), .d(new_n152), .out0(new_n155));
  xnrc02aa1n12x5               g060(.a(\b[11] ), .b(\a[12] ), .out0(new_n156));
  aoi012aa1n09x5               g061(.a(new_n129), .b(new_n97), .c(new_n130), .o1(new_n157));
  oao003aa1n06x5               g062(.a(\a[12] ), .b(\b[11] ), .c(new_n151), .carry(new_n158));
  oai013aa1d12x5               g063(.a(new_n158), .b(new_n156), .c(new_n152), .d(new_n157), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n155), .c(new_n119), .d(new_n126), .o1(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[12] ), .b(\a[13] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nano23aa1n03x7               g068(.a(new_n127), .b(new_n156), .c(new_n145), .d(new_n131), .out0(new_n164));
  aoi112aa1n02x5               g069(.a(new_n163), .b(new_n159), .c(new_n139), .d(new_n164), .o1(new_n165));
  aoi012aa1n02x5               g070(.a(new_n165), .b(new_n161), .c(new_n163), .o1(\s[13] ));
  orn002aa1n24x5               g071(.a(\a[13] ), .b(\b[12] ), .o(new_n167));
  aoai13aa1n03x5               g072(.a(new_n163), .b(new_n159), .c(new_n139), .d(new_n164), .o1(new_n168));
  xnrc02aa1n12x5               g073(.a(\b[13] ), .b(\a[14] ), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  xnbna2aa1n03x5               g075(.a(new_n170), .b(new_n168), .c(new_n167), .out0(\s[14] ));
  norp02aa1n02x5               g076(.a(new_n169), .b(new_n162), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n159), .c(new_n139), .d(new_n164), .o1(new_n173));
  oaoi03aa1n12x5               g078(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  nor002aa1d32x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nanp02aa1n04x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  norb02aa1n15x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  xnbna2aa1n03x5               g083(.a(new_n178), .b(new_n173), .c(new_n175), .out0(\s[15] ));
  aoai13aa1n02x5               g084(.a(new_n178), .b(new_n174), .c(new_n161), .d(new_n172), .o1(new_n180));
  nor022aa1n06x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nanp02aa1n04x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n182), .b(new_n181), .out0(new_n183));
  aoib12aa1n02x5               g088(.a(new_n176), .b(new_n182), .c(new_n181), .out0(new_n184));
  inv000aa1d42x5               g089(.a(new_n176), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n178), .o1(new_n186));
  aoai13aa1n03x5               g091(.a(new_n185), .b(new_n186), .c(new_n173), .d(new_n175), .o1(new_n187));
  aoi022aa1n02x7               g092(.a(new_n187), .b(new_n183), .c(new_n180), .d(new_n184), .o1(\s[16] ));
  nona23aa1n03x5               g093(.a(new_n182), .b(new_n177), .c(new_n176), .d(new_n181), .out0(new_n189));
  nor043aa1n02x5               g094(.a(new_n189), .b(new_n169), .c(new_n162), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n164), .b(new_n190), .o1(new_n191));
  oai012aa1n02x5               g096(.a(new_n182), .b(new_n181), .c(new_n176), .o1(new_n192));
  oaib12aa1n03x5               g097(.a(new_n192), .b(new_n189), .c(new_n174), .out0(new_n193));
  aoi012aa1n06x5               g098(.a(new_n193), .b(new_n159), .c(new_n190), .o1(new_n194));
  aoai13aa1n12x5               g099(.a(new_n194), .b(new_n191), .c(new_n119), .d(new_n126), .o1(new_n195));
  xorb03aa1n03x5               g100(.a(new_n195), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g101(.a(\a[17] ), .o1(new_n197));
  oaib12aa1n06x5               g102(.a(new_n195), .b(new_n197), .c(\b[16] ), .out0(new_n198));
  oaib12aa1n06x5               g103(.a(new_n198), .b(\b[16] ), .c(new_n197), .out0(new_n199));
  xorc02aa1n02x5               g104(.a(\a[18] ), .b(\b[17] ), .out0(new_n200));
  nor042aa1d18x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  norp02aa1n02x5               g106(.a(new_n200), .b(new_n201), .o1(new_n202));
  aoi022aa1n02x7               g107(.a(new_n199), .b(new_n200), .c(new_n198), .d(new_n202), .o1(\s[18] ));
  nano23aa1n06x5               g108(.a(new_n176), .b(new_n181), .c(new_n182), .d(new_n177), .out0(new_n204));
  nona22aa1n09x5               g109(.a(new_n204), .b(new_n169), .c(new_n162), .out0(new_n205));
  nor042aa1n03x5               g110(.a(new_n155), .b(new_n205), .o1(new_n206));
  nanb03aa1n02x5               g111(.a(new_n157), .b(new_n145), .c(new_n148), .out0(new_n207));
  aobi12aa1n06x5               g112(.a(new_n192), .b(new_n204), .c(new_n174), .out0(new_n208));
  aoai13aa1n09x5               g113(.a(new_n208), .b(new_n205), .c(new_n207), .d(new_n158), .o1(new_n209));
  inv040aa1d32x5               g114(.a(\a[18] ), .o1(new_n210));
  xroi22aa1d04x5               g115(.a(new_n197), .b(\b[16] ), .c(new_n210), .d(\b[17] ), .out0(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n209), .c(new_n139), .d(new_n206), .o1(new_n212));
  inv040aa1d32x5               g117(.a(\b[17] ), .o1(new_n213));
  oao003aa1n09x5               g118(.a(new_n210), .b(new_n213), .c(new_n201), .carry(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  xorc02aa1n12x5               g120(.a(\a[19] ), .b(\b[18] ), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n212), .c(new_n215), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g123(.a(new_n216), .b(new_n214), .c(new_n195), .d(new_n211), .o1(new_n219));
  xorc02aa1n03x5               g124(.a(\a[20] ), .b(\b[19] ), .out0(new_n220));
  inv000aa1d42x5               g125(.a(\a[19] ), .o1(new_n221));
  nanb02aa1d24x5               g126(.a(\b[18] ), .b(new_n221), .out0(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n220), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n216), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n222), .b(new_n224), .c(new_n212), .d(new_n215), .o1(new_n225));
  aoi022aa1n03x5               g130(.a(new_n225), .b(new_n220), .c(new_n219), .d(new_n223), .o1(\s[20] ));
  inv000aa1d42x5               g131(.a(\a[20] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n221), .b(\b[18] ), .c(new_n227), .d(\b[19] ), .out0(new_n228));
  and002aa1n02x5               g133(.a(new_n228), .b(new_n211), .o(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n209), .c(new_n139), .d(new_n206), .o1(new_n230));
  nand23aa1n06x5               g135(.a(new_n214), .b(new_n216), .c(new_n220), .o1(new_n231));
  oaoi03aa1n02x5               g136(.a(\a[20] ), .b(\b[19] ), .c(new_n222), .o1(new_n232));
  inv000aa1n06x5               g137(.a(new_n232), .o1(new_n233));
  nand02aa1d06x5               g138(.a(new_n231), .b(new_n233), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xorc02aa1n12x5               g140(.a(\a[21] ), .b(\b[20] ), .out0(new_n236));
  xnbna2aa1n03x5               g141(.a(new_n236), .b(new_n230), .c(new_n235), .out0(\s[21] ));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n234), .c(new_n195), .d(new_n229), .o1(new_n238));
  xorc02aa1n02x5               g143(.a(\a[22] ), .b(\b[21] ), .out0(new_n239));
  nor042aa1d18x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  norp02aa1n02x5               g145(.a(new_n239), .b(new_n240), .o1(new_n241));
  inv040aa1n08x5               g146(.a(new_n240), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[20] ), .b(\a[21] ), .out0(new_n243));
  aoai13aa1n03x5               g148(.a(new_n242), .b(new_n243), .c(new_n230), .d(new_n235), .o1(new_n244));
  aoi022aa1n03x5               g149(.a(new_n244), .b(new_n239), .c(new_n238), .d(new_n241), .o1(\s[22] ));
  xnrc02aa1n03x5               g150(.a(\b[21] ), .b(\a[22] ), .out0(new_n246));
  nor042aa1n03x5               g151(.a(new_n246), .b(new_n243), .o1(new_n247));
  and003aa1n02x5               g152(.a(new_n228), .b(new_n211), .c(new_n247), .o(new_n248));
  aoai13aa1n02x7               g153(.a(new_n248), .b(new_n209), .c(new_n139), .d(new_n206), .o1(new_n249));
  oaoi03aa1n03x5               g154(.a(\a[22] ), .b(\b[21] ), .c(new_n242), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n250), .b(new_n234), .c(new_n247), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n252), .c(new_n195), .d(new_n248), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n253), .b(new_n250), .c(new_n234), .d(new_n247), .o1(new_n255));
  aobi12aa1n02x7               g160(.a(new_n254), .b(new_n255), .c(new_n249), .out0(\s[23] ));
  xorc02aa1n12x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  nor002aa1d32x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  norp02aa1n02x5               g163(.a(new_n257), .b(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n258), .o1(new_n260));
  xnrc02aa1n02x5               g165(.a(\b[22] ), .b(\a[23] ), .out0(new_n261));
  aoai13aa1n03x5               g166(.a(new_n260), .b(new_n261), .c(new_n249), .d(new_n251), .o1(new_n262));
  aoi022aa1n03x5               g167(.a(new_n262), .b(new_n257), .c(new_n254), .d(new_n259), .o1(\s[24] ));
  xnrc02aa1n02x5               g168(.a(\b[23] ), .b(\a[24] ), .out0(new_n264));
  nona22aa1n09x5               g169(.a(new_n247), .b(new_n261), .c(new_n264), .out0(new_n265));
  nano22aa1n02x4               g170(.a(new_n265), .b(new_n211), .c(new_n228), .out0(new_n266));
  aoai13aa1n02x7               g171(.a(new_n266), .b(new_n209), .c(new_n139), .d(new_n206), .o1(new_n267));
  tech160nm_fioaoi03aa1n03p5x5 g172(.a(\a[24] ), .b(\b[23] ), .c(new_n260), .o1(new_n268));
  aoi013aa1n06x4               g173(.a(new_n268), .b(new_n250), .c(new_n253), .d(new_n257), .o1(new_n269));
  aoai13aa1n12x5               g174(.a(new_n269), .b(new_n265), .c(new_n231), .d(new_n233), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n270), .c(new_n195), .d(new_n266), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(new_n239), .b(new_n236), .o1(new_n273));
  nano22aa1n03x7               g178(.a(new_n273), .b(new_n253), .c(new_n257), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n232), .c(new_n214), .d(new_n228), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n271), .o1(new_n276));
  and003aa1n02x5               g181(.a(new_n275), .b(new_n276), .c(new_n269), .o(new_n277));
  aobi12aa1n02x7               g182(.a(new_n272), .b(new_n277), .c(new_n267), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  norp02aa1n02x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n270), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n280), .o1(new_n283));
  aoai13aa1n02x7               g188(.a(new_n283), .b(new_n276), .c(new_n267), .d(new_n282), .o1(new_n284));
  aoi022aa1n03x5               g189(.a(new_n284), .b(new_n279), .c(new_n272), .d(new_n281), .o1(\s[26] ));
  and002aa1n06x5               g190(.a(new_n279), .b(new_n271), .o(new_n286));
  nano32aa1n03x7               g191(.a(new_n265), .b(new_n286), .c(new_n211), .d(new_n228), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n287), .b(new_n209), .c(new_n139), .d(new_n206), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[25] ), .b(\a[26] ), .o1(new_n289));
  oai022aa1n02x5               g194(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n290));
  aoi022aa1n12x5               g195(.a(new_n270), .b(new_n286), .c(new_n289), .d(new_n290), .o1(new_n291));
  nor042aa1n03x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  and002aa1n24x5               g197(.a(\b[26] ), .b(\a[27] ), .o(new_n293));
  nor042aa1n03x5               g198(.a(new_n293), .b(new_n292), .o1(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n294), .b(new_n288), .c(new_n291), .out0(\s[27] ));
  inv000aa1n02x5               g200(.a(new_n286), .o1(new_n296));
  nanp02aa1n02x5               g201(.a(new_n290), .b(new_n289), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n296), .c(new_n275), .d(new_n269), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n293), .o1(new_n299));
  aoai13aa1n02x7               g204(.a(new_n299), .b(new_n298), .c(new_n195), .d(new_n287), .o1(new_n300));
  inv000aa1n03x5               g205(.a(new_n292), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n293), .c(new_n288), .d(new_n291), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(new_n303), .b(new_n292), .o1(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n300), .d(new_n304), .o1(\s[28] ));
  and002aa1n06x5               g210(.a(new_n303), .b(new_n294), .o(new_n306));
  aoai13aa1n02x7               g211(.a(new_n306), .b(new_n298), .c(new_n195), .d(new_n287), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n306), .o1(new_n308));
  oaoi03aa1n12x5               g213(.a(\a[28] ), .b(\b[27] ), .c(new_n301), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n308), .c(new_n288), .d(new_n291), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norp02aa1n02x5               g217(.a(new_n309), .b(new_n312), .o1(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n307), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g220(.a(new_n303), .b(new_n312), .c(new_n294), .o(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n298), .c(new_n195), .d(new_n287), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n316), .o1(new_n318));
  inv000aa1d42x5               g223(.a(\a[29] ), .o1(new_n319));
  inv000aa1d42x5               g224(.a(\b[28] ), .o1(new_n320));
  tech160nm_fioaoi03aa1n03p5x5 g225(.a(new_n319), .b(new_n320), .c(new_n309), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n318), .c(new_n288), .d(new_n291), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  oabi12aa1n02x5               g228(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n324), .b(new_n309), .c(new_n319), .d(new_n320), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n322), .b(new_n323), .c(new_n317), .d(new_n325), .o1(\s[30] ));
  nanp03aa1n02x5               g231(.a(new_n306), .b(new_n312), .c(new_n323), .o1(new_n327));
  inv000aa1n02x5               g232(.a(new_n327), .o1(new_n328));
  aoai13aa1n02x7               g233(.a(new_n328), .b(new_n298), .c(new_n195), .d(new_n287), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  oao003aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n331));
  norb02aa1n02x5               g236(.a(new_n331), .b(new_n330), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n331), .b(new_n327), .c(new_n288), .d(new_n291), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n333), .b(new_n330), .c(new_n329), .d(new_n332), .o1(\s[31] ));
  oai012aa1n02x5               g239(.a(new_n99), .b(new_n106), .c(new_n105), .o1(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g241(.a(\a[3] ), .b(\b[2] ), .c(new_n335), .o1(new_n337));
  xorb03aa1n02x5               g242(.a(new_n337), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnbna2aa1n03x5               g243(.a(new_n137), .b(new_n134), .c(new_n135), .out0(\s[5] ));
  nona22aa1n02x4               g244(.a(new_n134), .b(new_n110), .c(new_n112), .out0(new_n340));
  oaoi13aa1n02x5               g245(.a(new_n136), .b(new_n340), .c(new_n121), .d(new_n122), .o1(new_n341));
  oai112aa1n02x5               g246(.a(new_n340), .b(new_n136), .c(new_n122), .d(new_n121), .o1(new_n342));
  norb02aa1n02x5               g247(.a(new_n342), .b(new_n341), .out0(\s[6] ));
  norp02aa1n02x5               g248(.a(\b[5] ), .b(\a[6] ), .o1(new_n344));
  inv000aa1d42x5               g249(.a(new_n344), .o1(new_n345));
  norb02aa1n02x5               g250(.a(new_n116), .b(new_n115), .out0(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n342), .c(new_n345), .out0(\s[7] ));
  norb02aa1n02x5               g252(.a(new_n114), .b(new_n113), .out0(new_n348));
  aob012aa1n03x5               g253(.a(new_n346), .b(new_n342), .c(new_n345), .out0(new_n349));
  oai012aa1n02x5               g254(.a(new_n349), .b(\b[6] ), .c(\a[7] ), .o1(new_n350));
  aoib12aa1n02x5               g255(.a(new_n115), .b(new_n114), .c(new_n113), .out0(new_n351));
  aoi022aa1n02x5               g256(.a(new_n350), .b(new_n348), .c(new_n349), .d(new_n351), .o1(\s[8] ));
  xorb03aa1n02x5               g257(.a(new_n139), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


