// Benchmark "adder" written by ABC on Thu Jul 18 08:52:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n317,
    new_n320, new_n322, new_n323, new_n325, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n04x5   g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor002aa1d32x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[2] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[1] ), .o1(new_n101));
  nand22aa1n02x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  oaoi03aa1n03x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  norp02aa1n12x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor022aa1n08x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  inv000aa1d42x5               g013(.a(\a[3] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  aoai13aa1n04x5               g015(.a(new_n105), .b(new_n104), .c(new_n109), .d(new_n110), .o1(new_n111));
  oaih12aa1n06x5               g016(.a(new_n111), .b(new_n108), .c(new_n103), .o1(new_n112));
  nor042aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor042aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  tech160nm_finand02aa1n03p5x5 g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .out0(new_n118));
  xnrc02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .out0(new_n119));
  nor043aa1n03x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  orn002aa1n02x5               g025(.a(\a[5] ), .b(\b[4] ), .o(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  oai012aa1n02x5               g027(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n123));
  oaib12aa1n06x5               g028(.a(new_n123), .b(new_n117), .c(new_n122), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n112), .d(new_n120), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(\a[10] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(\b[9] ), .o1(new_n129));
  aoi012aa1n02x5               g034(.a(new_n98), .b(new_n128), .c(new_n129), .o1(new_n130));
  aoi022aa1n03x5               g035(.a(new_n126), .b(new_n130), .c(\b[9] ), .d(\a[10] ), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g037(.a(\a[11] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(\b[10] ), .o1(new_n134));
  oaoi03aa1n02x5               g039(.a(new_n133), .b(new_n134), .c(new_n131), .o1(new_n135));
  xnrb03aa1n02x5               g040(.a(new_n135), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nanp02aa1n03x5               g041(.a(new_n112), .b(new_n120), .o1(new_n137));
  nano23aa1n03x5               g042(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n138));
  aobi12aa1n03x5               g043(.a(new_n123), .b(new_n138), .c(new_n122), .out0(new_n139));
  nor022aa1n08x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nanp02aa1n12x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nor002aa1n16x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nano23aa1n09x5               g048(.a(new_n140), .b(new_n142), .c(new_n143), .d(new_n141), .out0(new_n144));
  nand23aa1n03x5               g049(.a(new_n144), .b(new_n97), .c(new_n125), .o1(new_n145));
  nona23aa1d18x5               g050(.a(new_n143), .b(new_n141), .c(new_n140), .d(new_n142), .out0(new_n146));
  oaoi03aa1n09x5               g051(.a(new_n128), .b(new_n129), .c(new_n98), .o1(new_n147));
  aoai13aa1n12x5               g052(.a(new_n143), .b(new_n142), .c(new_n133), .d(new_n134), .o1(new_n148));
  oai012aa1d24x5               g053(.a(new_n148), .b(new_n146), .c(new_n147), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n145), .c(new_n137), .d(new_n139), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g057(.a(\a[14] ), .o1(new_n153));
  nor042aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  tech160nm_fixorc02aa1n04x5   g059(.a(\a[13] ), .b(\b[12] ), .out0(new_n155));
  aoi012aa1n02x5               g060(.a(new_n154), .b(new_n151), .c(new_n155), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(new_n153), .out0(\s[14] ));
  xorc02aa1n02x5               g062(.a(\a[14] ), .b(\b[13] ), .out0(new_n158));
  and002aa1n02x5               g063(.a(new_n158), .b(new_n155), .o(new_n159));
  inv000aa1d42x5               g064(.a(\b[13] ), .o1(new_n160));
  oaoi03aa1n12x5               g065(.a(new_n153), .b(new_n160), .c(new_n154), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nor042aa1n04x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nand42aa1d28x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n162), .c(new_n151), .d(new_n159), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n165), .b(new_n162), .c(new_n151), .d(new_n159), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(\s[15] ));
  nor002aa1n03x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nand42aa1n16x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  oaoi13aa1n02x5               g077(.a(new_n172), .b(new_n166), .c(\a[15] ), .d(\b[14] ), .o1(new_n173));
  nona22aa1n02x4               g078(.a(new_n166), .b(new_n171), .c(new_n163), .out0(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(\s[16] ));
  nano23aa1n06x5               g080(.a(new_n163), .b(new_n169), .c(new_n170), .d(new_n164), .out0(new_n176));
  nand23aa1n03x5               g081(.a(new_n176), .b(new_n155), .c(new_n158), .o1(new_n177));
  nor042aa1n06x5               g082(.a(new_n177), .b(new_n145), .o1(new_n178));
  aoai13aa1n12x5               g083(.a(new_n178), .b(new_n124), .c(new_n112), .d(new_n120), .o1(new_n179));
  oai012aa1n02x5               g084(.a(new_n170), .b(new_n169), .c(new_n163), .o1(new_n180));
  oaib12aa1n02x5               g085(.a(new_n180), .b(new_n161), .c(new_n176), .out0(new_n181));
  aoib12aa1n12x5               g086(.a(new_n181), .b(new_n149), .c(new_n177), .out0(new_n182));
  nand02aa1d08x5               g087(.a(new_n179), .b(new_n182), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g089(.a(\a[18] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[17] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[16] ), .o1(new_n187));
  oaoi03aa1n02x5               g092(.a(new_n186), .b(new_n187), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  xroi22aa1d04x5               g094(.a(new_n186), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n190));
  nor002aa1n04x5               g095(.a(\b[17] ), .b(\a[18] ), .o1(new_n191));
  aoi112aa1n09x5               g096(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n192));
  nor042aa1n06x5               g097(.a(new_n192), .b(new_n191), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  nor022aa1n16x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand02aa1n04x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  norb02aa1n06x5               g101(.a(new_n196), .b(new_n195), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n194), .c(new_n183), .d(new_n190), .o1(new_n198));
  aoi112aa1n02x5               g103(.a(new_n197), .b(new_n194), .c(new_n183), .d(new_n190), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n20x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nand42aa1d28x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  norb02aa1n15x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  oaoi13aa1n06x5               g110(.a(new_n205), .b(new_n198), .c(\a[19] ), .d(\b[18] ), .o1(new_n206));
  nona22aa1n02x5               g111(.a(new_n198), .b(new_n204), .c(new_n195), .out0(new_n207));
  norb02aa1n03x4               g112(.a(new_n207), .b(new_n206), .out0(\s[20] ));
  nona23aa1n09x5               g113(.a(new_n203), .b(new_n196), .c(new_n195), .d(new_n202), .out0(new_n209));
  inv040aa1n03x5               g114(.a(new_n209), .o1(new_n210));
  nanp02aa1n02x5               g115(.a(new_n190), .b(new_n210), .o1(new_n211));
  oai012aa1n06x5               g116(.a(new_n203), .b(new_n202), .c(new_n195), .o1(new_n212));
  oai012aa1n18x5               g117(.a(new_n212), .b(new_n209), .c(new_n193), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  aoai13aa1n04x5               g119(.a(new_n214), .b(new_n211), .c(new_n179), .d(new_n182), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n16x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  xorc02aa1n12x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xorc02aa1n12x5               g123(.a(\a[22] ), .b(\b[21] ), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n215), .d(new_n218), .o1(new_n220));
  aoi112aa1n02x5               g125(.a(new_n217), .b(new_n219), .c(new_n215), .d(new_n218), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n220), .b(new_n221), .out0(\s[22] ));
  nand22aa1n12x5               g127(.a(new_n219), .b(new_n218), .o1(new_n223));
  nanb03aa1n06x5               g128(.a(new_n223), .b(new_n190), .c(new_n210), .out0(new_n224));
  oai112aa1n06x5               g129(.a(new_n197), .b(new_n204), .c(new_n192), .d(new_n191), .o1(new_n225));
  inv000aa1d42x5               g130(.a(\a[22] ), .o1(new_n226));
  inv020aa1d32x5               g131(.a(\b[21] ), .o1(new_n227));
  oaoi03aa1n12x5               g132(.a(new_n226), .b(new_n227), .c(new_n217), .o1(new_n228));
  aoai13aa1n12x5               g133(.a(new_n228), .b(new_n223), .c(new_n225), .d(new_n212), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n04x5               g135(.a(new_n230), .b(new_n224), .c(new_n179), .d(new_n182), .o1(new_n231));
  xorb03aa1n02x5               g136(.a(new_n231), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g137(.a(\b[22] ), .b(\a[23] ), .o1(new_n233));
  tech160nm_fixorc02aa1n02p5x5 g138(.a(\a[23] ), .b(\b[22] ), .out0(new_n234));
  xorc02aa1n02x5               g139(.a(\a[24] ), .b(\b[23] ), .out0(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n233), .c(new_n231), .d(new_n234), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(new_n233), .b(new_n235), .c(new_n231), .d(new_n234), .o1(new_n237));
  norb02aa1n03x4               g142(.a(new_n236), .b(new_n237), .out0(\s[24] ));
  and002aa1n02x5               g143(.a(new_n235), .b(new_n234), .o(new_n239));
  nona23aa1n02x4               g144(.a(new_n239), .b(new_n190), .c(new_n223), .d(new_n209), .out0(new_n240));
  inv000aa1d42x5               g145(.a(\a[24] ), .o1(new_n241));
  inv000aa1d42x5               g146(.a(\b[23] ), .o1(new_n242));
  oao003aa1n02x5               g147(.a(new_n241), .b(new_n242), .c(new_n233), .carry(new_n243));
  tech160nm_fiaoi012aa1n05x5   g148(.a(new_n243), .b(new_n229), .c(new_n239), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n240), .c(new_n179), .d(new_n182), .o1(new_n245));
  xorb03aa1n02x5               g150(.a(new_n245), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g151(.a(\b[24] ), .b(\a[25] ), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[25] ), .b(\b[24] ), .out0(new_n248));
  tech160nm_fixorc02aa1n04x5   g153(.a(\a[26] ), .b(\b[25] ), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n247), .c(new_n245), .d(new_n248), .o1(new_n250));
  aoi112aa1n03x5               g155(.a(new_n247), .b(new_n249), .c(new_n245), .d(new_n248), .o1(new_n251));
  norb02aa1n03x4               g156(.a(new_n250), .b(new_n251), .out0(\s[26] ));
  oao003aa1n02x5               g157(.a(new_n100), .b(new_n101), .c(new_n102), .carry(new_n253));
  nano23aa1n02x4               g158(.a(new_n104), .b(new_n106), .c(new_n107), .d(new_n105), .out0(new_n254));
  aobi12aa1n02x5               g159(.a(new_n111), .b(new_n254), .c(new_n253), .out0(new_n255));
  nona22aa1n02x4               g160(.a(new_n138), .b(new_n118), .c(new_n119), .out0(new_n256));
  oai012aa1n02x7               g161(.a(new_n139), .b(new_n255), .c(new_n256), .o1(new_n257));
  nanb02aa1n02x5               g162(.a(new_n147), .b(new_n144), .out0(new_n258));
  aobi12aa1n02x5               g163(.a(new_n180), .b(new_n162), .c(new_n176), .out0(new_n259));
  aoai13aa1n02x5               g164(.a(new_n259), .b(new_n177), .c(new_n258), .d(new_n148), .o1(new_n260));
  and002aa1n06x5               g165(.a(new_n249), .b(new_n248), .o(new_n261));
  nano22aa1n03x7               g166(.a(new_n224), .b(new_n239), .c(new_n261), .out0(new_n262));
  aoai13aa1n06x5               g167(.a(new_n262), .b(new_n260), .c(new_n257), .d(new_n178), .o1(new_n263));
  aoai13aa1n09x5               g168(.a(new_n261), .b(new_n243), .c(new_n229), .d(new_n239), .o1(new_n264));
  oai022aa1n02x5               g169(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n265));
  aob012aa1n02x5               g170(.a(new_n265), .b(\b[25] ), .c(\a[26] ), .out0(new_n266));
  xorc02aa1n12x5               g171(.a(\a[27] ), .b(\b[26] ), .out0(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoi013aa1n06x4               g173(.a(new_n268), .b(new_n263), .c(new_n264), .d(new_n266), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n262), .o1(new_n270));
  aoi012aa1n06x5               g175(.a(new_n270), .b(new_n179), .c(new_n182), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n223), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n228), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n239), .b(new_n273), .c(new_n213), .d(new_n272), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n243), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n261), .o1(new_n276));
  aoai13aa1n04x5               g181(.a(new_n266), .b(new_n276), .c(new_n274), .d(new_n275), .o1(new_n277));
  norp03aa1n02x5               g182(.a(new_n277), .b(new_n271), .c(new_n267), .o1(new_n278));
  norp02aa1n02x5               g183(.a(new_n269), .b(new_n278), .o1(\s[27] ));
  nor042aa1n03x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  oaih12aa1n02x5               g186(.a(new_n267), .b(new_n277), .c(new_n271), .o1(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n283), .b(new_n282), .c(new_n281), .o1(new_n284));
  nano22aa1n03x7               g189(.a(new_n269), .b(new_n281), .c(new_n283), .out0(new_n285));
  nor002aa1n02x5               g190(.a(new_n284), .b(new_n285), .o1(\s[28] ));
  norb02aa1n02x5               g191(.a(new_n267), .b(new_n283), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n277), .c(new_n271), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n281), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[28] ), .b(\a[29] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  inv000aa1n02x5               g196(.a(new_n287), .o1(new_n292));
  aoi013aa1n02x5               g197(.a(new_n292), .b(new_n263), .c(new_n264), .d(new_n266), .o1(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n290), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n291), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n06x5               g201(.a(new_n267), .b(new_n290), .c(new_n283), .out0(new_n297));
  oaih12aa1n02x5               g202(.a(new_n297), .b(new_n277), .c(new_n271), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[29] ), .b(\a[30] ), .out0(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n298), .c(new_n299), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n297), .o1(new_n302));
  aoi013aa1n02x5               g207(.a(new_n302), .b(new_n263), .c(new_n264), .d(new_n266), .o1(new_n303));
  nano22aa1n03x5               g208(.a(new_n303), .b(new_n299), .c(new_n300), .out0(new_n304));
  norp02aa1n03x5               g209(.a(new_n301), .b(new_n304), .o1(\s[30] ));
  norb02aa1n03x4               g210(.a(new_n297), .b(new_n300), .out0(new_n306));
  inv020aa1n02x5               g211(.a(new_n306), .o1(new_n307));
  aoi013aa1n02x5               g212(.a(new_n307), .b(new_n263), .c(new_n264), .d(new_n266), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  nano22aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n310), .out0(new_n311));
  oaih12aa1n02x5               g216(.a(new_n306), .b(new_n277), .c(new_n271), .o1(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n310), .b(new_n312), .c(new_n309), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n313), .b(new_n311), .o1(\s[31] ));
  xorb03aa1n02x5               g219(.a(new_n103), .b(\b[2] ), .c(new_n109), .out0(\s[3] ));
  nanb03aa1n02x5               g220(.a(new_n106), .b(new_n253), .c(new_n107), .out0(new_n316));
  aboi22aa1n03x5               g221(.a(new_n104), .b(new_n105), .c(new_n109), .d(new_n110), .out0(new_n317));
  aboi22aa1n03x5               g222(.a(new_n104), .b(new_n112), .c(new_n316), .d(new_n317), .out0(\s[4] ));
  xorb03aa1n02x5               g223(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g224(.a(\a[5] ), .b(\b[4] ), .c(new_n255), .o1(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oao003aa1n02x5               g226(.a(\a[5] ), .b(\b[4] ), .c(new_n255), .carry(new_n322));
  tech160nm_fioaoi03aa1n03p5x5 g227(.a(\a[6] ), .b(\b[5] ), .c(new_n322), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  inv000aa1d42x5               g229(.a(\a[8] ), .o1(new_n325));
  aoi012aa1n02x5               g230(.a(new_n115), .b(new_n323), .c(new_n116), .o1(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[7] ), .c(new_n325), .out0(\s[8] ));
  xnbna2aa1n03x5               g232(.a(new_n125), .b(new_n137), .c(new_n139), .out0(\s[9] ));
endmodule


