// Benchmark "adder" written by ABC on Thu Jul 18 08:58:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n321, new_n323, new_n325;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n02p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  and002aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[8] ), .o1(new_n100));
  nanb02aa1n03x5               g005(.a(\a[9] ), .b(new_n100), .out0(new_n101));
  xnrc02aa1n12x5               g006(.a(\b[7] ), .b(\a[8] ), .out0(new_n102));
  xnrc02aa1n12x5               g007(.a(\b[6] ), .b(\a[7] ), .out0(new_n103));
  oai022aa1d24x5               g008(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n104));
  aob012aa1d15x5               g009(.a(new_n104), .b(\b[5] ), .c(\a[6] ), .out0(new_n105));
  inv000aa1d42x5               g010(.a(\a[8] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[7] ), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  tech160nm_fioaoi03aa1n02p5x5 g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  oai013aa1n09x5               g014(.a(new_n109), .b(new_n105), .c(new_n102), .d(new_n103), .o1(new_n110));
  inv000aa1d42x5               g015(.a(new_n110), .o1(new_n111));
  norp02aa1n04x5               g016(.a(new_n103), .b(new_n102), .o1(new_n112));
  nor002aa1n02x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nor042aa1n12x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nona23aa1n03x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nand42aa1n02x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  nor042aa1n06x5               g023(.a(\b[1] ), .b(\a[2] ), .o1(new_n119));
  nand22aa1n06x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  oaih12aa1n06x5               g025(.a(new_n118), .b(new_n119), .c(new_n120), .o1(new_n121));
  inv040aa1n03x5               g026(.a(new_n115), .o1(new_n122));
  oaoi03aa1n09x5               g027(.a(\a[4] ), .b(\b[3] ), .c(new_n122), .o1(new_n123));
  oabi12aa1n02x7               g028(.a(new_n123), .b(new_n117), .c(new_n121), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[5] ), .b(\a[6] ), .out0(new_n125));
  xnrc02aa1n02x5               g030(.a(\b[4] ), .b(\a[5] ), .out0(new_n126));
  nor042aa1n02x5               g031(.a(new_n126), .b(new_n125), .o1(new_n127));
  nanp03aa1n03x5               g032(.a(new_n124), .b(new_n112), .c(new_n127), .o1(new_n128));
  nand23aa1n03x5               g033(.a(new_n128), .b(new_n101), .c(new_n111), .o1(new_n129));
  xobna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  tech160nm_fixorc02aa1n05x5   g035(.a(\a[11] ), .b(\b[10] ), .out0(new_n131));
  norp02aa1n02x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  aoai13aa1n06x5               g038(.a(new_n133), .b(new_n132), .c(new_n129), .d(new_n99), .o1(new_n134));
  xnrc02aa1n02x5               g039(.a(new_n134), .b(new_n131), .out0(\s[11] ));
  nor042aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  aoi012aa1n03x5               g041(.a(new_n132), .b(new_n129), .c(new_n99), .o1(new_n137));
  nano22aa1n03x7               g042(.a(new_n137), .b(new_n133), .c(new_n131), .out0(new_n138));
  xnrc02aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .out0(new_n139));
  oai012aa1n02x5               g044(.a(new_n139), .b(new_n138), .c(new_n136), .o1(new_n140));
  inv000aa1n02x5               g045(.a(new_n136), .o1(new_n141));
  xnrc02aa1n02x5               g046(.a(\b[10] ), .b(\a[11] ), .out0(new_n142));
  xorc02aa1n02x5               g047(.a(\a[12] ), .b(\b[11] ), .out0(new_n143));
  oai112aa1n02x5               g048(.a(new_n141), .b(new_n143), .c(new_n134), .d(new_n142), .o1(new_n144));
  nanp02aa1n02x5               g049(.a(new_n140), .b(new_n144), .o1(\s[12] ));
  oaoi03aa1n02x5               g050(.a(\a[10] ), .b(\b[9] ), .c(new_n101), .o1(new_n146));
  nand43aa1n02x5               g051(.a(new_n146), .b(new_n131), .c(new_n143), .o1(new_n147));
  oao003aa1n02x5               g052(.a(\a[12] ), .b(\b[11] ), .c(new_n141), .carry(new_n148));
  and002aa1n02x5               g053(.a(new_n147), .b(new_n148), .o(new_n149));
  xnrc02aa1n03x5               g054(.a(\b[8] ), .b(\a[9] ), .out0(new_n150));
  nona23aa1n03x5               g055(.a(new_n143), .b(new_n97), .c(new_n150), .d(new_n142), .out0(new_n151));
  aoai13aa1n02x5               g056(.a(new_n149), .b(new_n151), .c(new_n128), .d(new_n111), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d28x5               g058(.a(\a[14] ), .o1(new_n154));
  nor022aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  xnrc02aa1n12x5               g060(.a(\b[12] ), .b(\a[13] ), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoi012aa1n03x5               g062(.a(new_n155), .b(new_n152), .c(new_n157), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(new_n154), .out0(\s[14] ));
  nano23aa1n03x5               g064(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n160));
  inv020aa1n03x5               g065(.a(new_n121), .o1(new_n161));
  tech160nm_fiaoi012aa1n05x5   g066(.a(new_n123), .b(new_n160), .c(new_n161), .o1(new_n162));
  nano22aa1n03x7               g067(.a(new_n162), .b(new_n112), .c(new_n127), .out0(new_n163));
  oabi12aa1n03x5               g068(.a(new_n151), .b(new_n163), .c(new_n110), .out0(new_n164));
  xnrc02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .out0(new_n165));
  norp02aa1n02x5               g070(.a(new_n165), .b(new_n156), .o1(new_n166));
  inv000aa1n02x5               g071(.a(new_n166), .o1(new_n167));
  inv040aa1d32x5               g072(.a(\b[13] ), .o1(new_n168));
  oaoi03aa1n02x5               g073(.a(new_n154), .b(new_n168), .c(new_n155), .o1(new_n169));
  aoai13aa1n04x5               g074(.a(new_n169), .b(new_n167), .c(new_n164), .d(new_n149), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  nor002aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanp02aa1n04x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  aoai13aa1n03x5               g082(.a(new_n177), .b(new_n172), .c(new_n170), .d(new_n174), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(new_n170), .b(new_n174), .o1(new_n179));
  nona22aa1n02x4               g084(.a(new_n179), .b(new_n177), .c(new_n172), .out0(new_n180));
  nanp02aa1n02x5               g085(.a(new_n180), .b(new_n178), .o1(\s[16] ));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  nano23aa1n09x5               g087(.a(new_n172), .b(new_n175), .c(new_n176), .d(new_n173), .out0(new_n183));
  oao003aa1n02x5               g088(.a(new_n154), .b(new_n168), .c(new_n155), .carry(new_n184));
  oa0012aa1n02x5               g089(.a(new_n176), .b(new_n175), .c(new_n172), .o(new_n185));
  tech160nm_fiaoi012aa1n03p5x5 g090(.a(new_n185), .b(new_n183), .c(new_n184), .o1(new_n186));
  nona22aa1n03x5               g091(.a(new_n183), .b(new_n165), .c(new_n156), .out0(new_n187));
  aoai13aa1n06x5               g092(.a(new_n186), .b(new_n187), .c(new_n147), .d(new_n148), .o1(new_n188));
  nor042aa1n03x5               g093(.a(new_n151), .b(new_n187), .o1(new_n189));
  oaoi13aa1n12x5               g094(.a(new_n188), .b(new_n189), .c(new_n163), .d(new_n110), .o1(new_n190));
  xorb03aa1n03x5               g095(.a(new_n190), .b(\b[16] ), .c(new_n182), .out0(\s[17] ));
  oaoi03aa1n03x5               g096(.a(\a[17] ), .b(\b[16] ), .c(new_n190), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g098(.a(\a[18] ), .o1(new_n194));
  xroi22aa1d06x4               g099(.a(new_n182), .b(\b[16] ), .c(new_n194), .d(\b[17] ), .out0(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  oai022aa1n02x7               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oaib12aa1n09x5               g102(.a(new_n197), .b(new_n194), .c(\b[17] ), .out0(new_n198));
  tech160nm_fioai012aa1n05x5   g103(.a(new_n198), .b(new_n190), .c(new_n196), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n20x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1n08x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  nor022aa1n16x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand02aa1n08x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  aoai13aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n199), .d(new_n204), .o1(new_n208));
  aoi013aa1n06x4               g113(.a(new_n110), .b(new_n124), .c(new_n112), .d(new_n127), .o1(new_n209));
  inv000aa1n02x5               g114(.a(new_n189), .o1(new_n210));
  oabi12aa1n06x5               g115(.a(new_n188), .b(new_n209), .c(new_n210), .out0(new_n211));
  nanb02aa1n02x5               g116(.a(\b[16] ), .b(new_n182), .out0(new_n212));
  oaoi03aa1n02x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n212), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n204), .b(new_n213), .c(new_n211), .d(new_n195), .o1(new_n214));
  nona22aa1n03x5               g119(.a(new_n214), .b(new_n207), .c(new_n202), .out0(new_n215));
  nanp02aa1n03x5               g120(.a(new_n208), .b(new_n215), .o1(\s[20] ));
  nona23aa1d18x5               g121(.a(new_n206), .b(new_n203), .c(new_n202), .d(new_n205), .out0(new_n217));
  oa0012aa1n03x5               g122(.a(new_n206), .b(new_n205), .c(new_n202), .o(new_n218));
  oabi12aa1n18x5               g123(.a(new_n218), .b(new_n198), .c(new_n217), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  xorc02aa1n02x5               g125(.a(\a[17] ), .b(\b[16] ), .out0(new_n221));
  xnrc02aa1n02x5               g126(.a(\b[17] ), .b(\a[18] ), .out0(new_n222));
  norb03aa1d15x5               g127(.a(new_n221), .b(new_n217), .c(new_n222), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  tech160nm_fioai012aa1n05x5   g129(.a(new_n220), .b(new_n190), .c(new_n224), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[20] ), .b(\a[21] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  tech160nm_fixnrc02aa1n05x5   g134(.a(\b[21] ), .b(\a[22] ), .out0(new_n230));
  aoai13aa1n03x5               g135(.a(new_n230), .b(new_n227), .c(new_n225), .d(new_n229), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n229), .b(new_n219), .c(new_n211), .d(new_n223), .o1(new_n232));
  nona22aa1n02x4               g137(.a(new_n232), .b(new_n230), .c(new_n227), .out0(new_n233));
  nanp02aa1n03x5               g138(.a(new_n231), .b(new_n233), .o1(\s[22] ));
  nor042aa1n09x5               g139(.a(new_n230), .b(new_n228), .o1(new_n235));
  inv000aa1d42x5               g140(.a(\a[22] ), .o1(new_n236));
  inv040aa1d32x5               g141(.a(\b[21] ), .o1(new_n237));
  oao003aa1n12x5               g142(.a(new_n236), .b(new_n237), .c(new_n227), .carry(new_n238));
  aoi012aa1d24x5               g143(.a(new_n238), .b(new_n219), .c(new_n235), .o1(new_n239));
  nano23aa1d18x5               g144(.a(new_n202), .b(new_n205), .c(new_n206), .d(new_n203), .out0(new_n240));
  nand23aa1d12x5               g145(.a(new_n195), .b(new_n235), .c(new_n240), .o1(new_n241));
  tech160nm_fioai012aa1n05x5   g146(.a(new_n239), .b(new_n190), .c(new_n241), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[23] ), .b(\a[24] ), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n244), .c(new_n242), .d(new_n245), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n239), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n241), .o1(new_n249));
  aoai13aa1n02x5               g154(.a(new_n245), .b(new_n248), .c(new_n211), .d(new_n249), .o1(new_n250));
  nona22aa1n03x5               g155(.a(new_n250), .b(new_n246), .c(new_n244), .out0(new_n251));
  nanp02aa1n02x5               g156(.a(new_n247), .b(new_n251), .o1(\s[24] ));
  norb02aa1n03x5               g157(.a(new_n245), .b(new_n246), .out0(new_n253));
  inv040aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  nano32aa1n03x7               g159(.a(new_n254), .b(new_n195), .c(new_n235), .d(new_n240), .out0(new_n255));
  inv020aa1n02x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n235), .b(new_n218), .c(new_n240), .d(new_n213), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n238), .o1(new_n258));
  oai022aa1n02x5               g163(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n259));
  aob012aa1n02x5               g164(.a(new_n259), .b(\b[23] ), .c(\a[24] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n254), .c(new_n257), .d(new_n258), .o1(new_n261));
  inv030aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  tech160nm_fioai012aa1n05x5   g167(.a(new_n262), .b(new_n190), .c(new_n256), .o1(new_n263));
  xorb03aa1n02x5               g168(.a(new_n263), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  tech160nm_fixorc02aa1n04x5   g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  tech160nm_fixnrc02aa1n02p5x5 g171(.a(\b[25] ), .b(\a[26] ), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n265), .c(new_n263), .d(new_n266), .o1(new_n268));
  aoai13aa1n02x5               g173(.a(new_n266), .b(new_n261), .c(new_n211), .d(new_n255), .o1(new_n269));
  nona22aa1n03x5               g174(.a(new_n269), .b(new_n267), .c(new_n265), .out0(new_n270));
  nanp02aa1n03x5               g175(.a(new_n268), .b(new_n270), .o1(\s[26] ));
  nanp02aa1n02x5               g176(.a(\b[25] ), .b(\a[26] ), .o1(new_n272));
  norb02aa1n06x5               g177(.a(new_n266), .b(new_n267), .out0(new_n273));
  oai022aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n274));
  aoi022aa1n06x5               g179(.a(new_n261), .b(new_n273), .c(new_n272), .d(new_n274), .o1(new_n275));
  nano22aa1d15x5               g180(.a(new_n241), .b(new_n253), .c(new_n273), .out0(new_n276));
  inv020aa1n03x5               g181(.a(new_n276), .o1(new_n277));
  oai012aa1n12x5               g182(.a(new_n275), .b(new_n190), .c(new_n277), .o1(new_n278));
  xorb03aa1n02x5               g183(.a(new_n278), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  xorc02aa1n02x5               g185(.a(\a[27] ), .b(\b[26] ), .out0(new_n281));
  xnrc02aa1n02x5               g186(.a(\b[27] ), .b(\a[28] ), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n282), .b(new_n280), .c(new_n278), .d(new_n281), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n253), .b(new_n238), .c(new_n219), .d(new_n235), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n273), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n274), .b(new_n272), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n285), .c(new_n284), .d(new_n260), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n281), .b(new_n287), .c(new_n211), .d(new_n276), .o1(new_n288));
  nona22aa1n02x5               g193(.a(new_n288), .b(new_n282), .c(new_n280), .out0(new_n289));
  nanp02aa1n03x5               g194(.a(new_n283), .b(new_n289), .o1(\s[28] ));
  norb02aa1n02x5               g195(.a(new_n281), .b(new_n282), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n287), .c(new_n211), .d(new_n276), .o1(new_n292));
  inv000aa1n03x5               g197(.a(new_n280), .o1(new_n293));
  oaoi03aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n293), .o1(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  nona22aa1n02x5               g200(.a(new_n292), .b(new_n294), .c(new_n295), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n295), .b(new_n294), .c(new_n278), .d(new_n291), .o1(new_n297));
  nanp02aa1n03x5               g202(.a(new_n297), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g204(.a(new_n281), .b(new_n295), .c(new_n282), .out0(new_n300));
  oao003aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n293), .carry(new_n301));
  oaoi03aa1n02x5               g206(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .o1(new_n302));
  tech160nm_fixorc02aa1n03p5x5 g207(.a(\a[30] ), .b(\b[29] ), .out0(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n302), .c(new_n278), .d(new_n300), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n300), .b(new_n287), .c(new_n211), .d(new_n276), .o1(new_n306));
  nona22aa1n02x5               g211(.a(new_n306), .b(new_n302), .c(new_n304), .out0(new_n307));
  nanp02aa1n03x5               g212(.a(new_n305), .b(new_n307), .o1(\s[30] ));
  nanp02aa1n02x5               g213(.a(new_n302), .b(new_n303), .o1(new_n309));
  oai012aa1n02x5               g214(.a(new_n309), .b(\b[29] ), .c(\a[30] ), .o1(new_n310));
  nano23aa1n02x4               g215(.a(new_n295), .b(new_n282), .c(new_n303), .d(new_n281), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n287), .c(new_n211), .d(new_n276), .o1(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[30] ), .b(\a[31] ), .out0(new_n313));
  nona22aa1n02x5               g218(.a(new_n312), .b(new_n313), .c(new_n310), .out0(new_n314));
  aoai13aa1n03x5               g219(.a(new_n313), .b(new_n310), .c(new_n278), .d(new_n311), .o1(new_n315));
  nanp02aa1n03x5               g220(.a(new_n315), .b(new_n314), .o1(\s[31] ));
  xnbna2aa1n03x5               g221(.a(new_n121), .b(new_n122), .c(new_n116), .out0(\s[3] ));
  oaoi03aa1n02x5               g222(.a(\a[3] ), .b(\b[2] ), .c(new_n121), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g224(.a(new_n124), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g225(.a(\a[5] ), .b(\b[4] ), .c(new_n162), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaib12aa1n02x5               g227(.a(new_n105), .b(new_n162), .c(new_n127), .out0(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoib12aa1n02x5               g229(.a(new_n108), .b(new_n323), .c(new_n103), .out0(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[7] ), .c(new_n106), .out0(\s[8] ));
  xobna2aa1n03x5               g231(.a(new_n150), .b(new_n128), .c(new_n111), .out0(\s[9] ));
endmodule


