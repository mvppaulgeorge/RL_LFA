// Benchmark "adder" written by ABC on Wed Jul 17 21:57:02 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n349, new_n351, new_n353,
    new_n355, new_n357, new_n358, new_n360;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n12x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor042aa1n06x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  xorc02aa1n12x5               g005(.a(\a[4] ), .b(\b[3] ), .out0(new_n101));
  nand42aa1n06x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nor042aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano22aa1n03x7               g009(.a(new_n103), .b(new_n102), .c(new_n104), .out0(new_n105));
  nand22aa1n04x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nona22aa1n09x5               g012(.a(new_n102), .b(new_n107), .c(new_n106), .out0(new_n108));
  inv000aa1d42x5               g013(.a(\a[4] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[3] ), .o1(new_n110));
  oaoi03aa1n09x5               g015(.a(new_n109), .b(new_n110), .c(new_n103), .o1(new_n111));
  inv000aa1n02x5               g016(.a(new_n111), .o1(new_n112));
  aoi013aa1n06x4               g017(.a(new_n112), .b(new_n108), .c(new_n105), .d(new_n101), .o1(new_n113));
  nor042aa1d18x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  norb02aa1n12x5               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nand02aa1d06x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nor002aa1d24x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nanb02aa1n03x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  xorc02aa1n06x5               g025(.a(\a[8] ), .b(\b[7] ), .out0(new_n121));
  nona23aa1n09x5               g026(.a(new_n121), .b(new_n116), .c(new_n117), .d(new_n120), .out0(new_n122));
  inv000aa1d42x5               g027(.a(\a[8] ), .o1(new_n123));
  oai022aa1d18x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  aoai13aa1n03x5               g029(.a(new_n115), .b(new_n114), .c(new_n124), .d(new_n118), .o1(new_n125));
  oaib12aa1n03x5               g030(.a(new_n125), .b(\b[7] ), .c(new_n123), .out0(new_n126));
  oaib12aa1n12x5               g031(.a(new_n126), .b(new_n123), .c(\b[7] ), .out0(new_n127));
  oai012aa1n18x5               g032(.a(new_n127), .b(new_n113), .c(new_n122), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n99), .b(new_n100), .c(new_n128), .d(new_n129), .o1(new_n130));
  xnrc02aa1n02x5               g035(.a(\b[3] ), .b(\a[4] ), .out0(new_n131));
  nanb03aa1n02x5               g036(.a(new_n103), .b(new_n104), .c(new_n102), .out0(new_n132));
  norb03aa1n03x5               g037(.a(new_n102), .b(new_n107), .c(new_n106), .out0(new_n133));
  oai013aa1n03x5               g038(.a(new_n111), .b(new_n133), .c(new_n132), .d(new_n131), .o1(new_n134));
  tech160nm_fixorc02aa1n03p5x5 g039(.a(\a[5] ), .b(\b[4] ), .out0(new_n135));
  nanp02aa1n02x5               g040(.a(new_n135), .b(new_n116), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n119), .o1(new_n137));
  nano32aa1n03x5               g042(.a(new_n136), .b(new_n121), .c(new_n118), .d(new_n137), .out0(new_n138));
  oaoi03aa1n02x5               g043(.a(\a[8] ), .b(\b[7] ), .c(new_n125), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n129), .b(new_n139), .c(new_n134), .d(new_n138), .o1(new_n140));
  norb03aa1n02x5               g045(.a(new_n98), .b(new_n97), .c(new_n100), .out0(new_n141));
  nand42aa1n03x5               g046(.a(new_n140), .b(new_n141), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(new_n130), .b(new_n142), .o1(\s[10] ));
  nand42aa1n08x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nor002aa1d32x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  nanb03aa1n02x5               g050(.a(new_n145), .b(new_n98), .c(new_n144), .out0(new_n146));
  nanb02aa1n02x5               g051(.a(new_n146), .b(new_n142), .out0(new_n147));
  inv030aa1n04x5               g052(.a(new_n145), .o1(new_n148));
  aoi022aa1n02x5               g053(.a(new_n142), .b(new_n98), .c(new_n148), .d(new_n144), .o1(new_n149));
  norb02aa1n02x7               g054(.a(new_n147), .b(new_n149), .out0(\s[11] ));
  nor002aa1d32x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nand02aa1d16x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  norb02aa1n06x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n151), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n145), .b(new_n154), .c(new_n152), .o1(new_n155));
  aoai13aa1n02x5               g060(.a(new_n148), .b(new_n146), .c(new_n140), .d(new_n141), .o1(new_n156));
  aoi022aa1n02x5               g061(.a(new_n147), .b(new_n155), .c(new_n156), .d(new_n153), .o1(\s[12] ));
  nanb02aa1n12x5               g062(.a(new_n145), .b(new_n144), .out0(new_n158));
  nona23aa1d24x5               g063(.a(new_n153), .b(new_n129), .c(new_n99), .d(new_n158), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n139), .c(new_n134), .d(new_n138), .o1(new_n161));
  nanb03aa1n06x5               g066(.a(new_n151), .b(new_n152), .c(new_n144), .out0(new_n162));
  oai112aa1n04x5               g067(.a(new_n148), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n163));
  aoi012aa1n06x5               g068(.a(new_n151), .b(new_n145), .c(new_n152), .o1(new_n164));
  oai012aa1n12x5               g069(.a(new_n164), .b(new_n163), .c(new_n162), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  nor042aa1n06x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  nand42aa1n06x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n161), .c(new_n166), .out0(\s[13] ));
  nanp02aa1n06x5               g075(.a(new_n161), .b(new_n166), .o1(new_n171));
  nor042aa1n06x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nand42aa1n16x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  aoi112aa1n02x5               g079(.a(new_n167), .b(new_n174), .c(new_n171), .d(new_n169), .o1(new_n175));
  aoai13aa1n02x5               g080(.a(new_n174), .b(new_n167), .c(new_n171), .d(new_n168), .o1(new_n176));
  norb02aa1n03x4               g081(.a(new_n176), .b(new_n175), .out0(\s[14] ));
  nano23aa1n09x5               g082(.a(new_n167), .b(new_n172), .c(new_n173), .d(new_n168), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n165), .c(new_n128), .d(new_n160), .o1(new_n179));
  oai012aa1n18x5               g084(.a(new_n173), .b(new_n172), .c(new_n167), .o1(new_n180));
  xnrc02aa1n12x5               g085(.a(\b[14] ), .b(\a[15] ), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n179), .c(new_n180), .out0(\s[15] ));
  inv000aa1d42x5               g088(.a(new_n180), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n182), .b(new_n184), .c(new_n171), .d(new_n178), .o1(new_n185));
  xnrc02aa1n12x5               g090(.a(\b[15] ), .b(\a[16] ), .out0(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  nor042aa1n06x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  norb02aa1n02x5               g093(.a(new_n186), .b(new_n188), .out0(new_n189));
  inv000aa1d42x5               g094(.a(new_n188), .o1(new_n190));
  aoai13aa1n02x5               g095(.a(new_n190), .b(new_n181), .c(new_n179), .d(new_n180), .o1(new_n191));
  aoi022aa1n03x5               g096(.a(new_n191), .b(new_n187), .c(new_n185), .d(new_n189), .o1(\s[16] ));
  nor042aa1n06x5               g097(.a(new_n186), .b(new_n181), .o1(new_n193));
  nano22aa1d15x5               g098(.a(new_n159), .b(new_n178), .c(new_n193), .out0(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n139), .c(new_n134), .d(new_n138), .o1(new_n195));
  aoai13aa1n06x5               g100(.a(new_n193), .b(new_n184), .c(new_n165), .d(new_n178), .o1(new_n196));
  oao003aa1n02x5               g101(.a(\a[16] ), .b(\b[15] ), .c(new_n190), .carry(new_n197));
  nanp03aa1d12x5               g102(.a(new_n195), .b(new_n196), .c(new_n197), .o1(new_n198));
  xorc02aa1n12x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  nano22aa1n02x4               g104(.a(new_n199), .b(new_n196), .c(new_n197), .out0(new_n200));
  aoi022aa1n02x5               g105(.a(new_n198), .b(new_n199), .c(new_n200), .d(new_n195), .o1(\s[17] ));
  inv000aa1d42x5               g106(.a(\a[17] ), .o1(new_n202));
  nanb02aa1n02x5               g107(.a(\b[16] ), .b(new_n202), .out0(new_n203));
  inv000aa1n02x5               g108(.a(new_n193), .o1(new_n204));
  nano22aa1n03x5               g109(.a(new_n151), .b(new_n144), .c(new_n152), .out0(new_n205));
  oai012aa1n02x5               g110(.a(new_n98), .b(\b[10] ), .c(\a[11] ), .o1(new_n206));
  oab012aa1n02x4               g111(.a(new_n206), .b(new_n97), .c(new_n100), .out0(new_n207));
  inv020aa1n02x5               g112(.a(new_n164), .o1(new_n208));
  aoai13aa1n04x5               g113(.a(new_n178), .b(new_n208), .c(new_n207), .d(new_n205), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n197), .b(new_n204), .c(new_n209), .d(new_n180), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n199), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n211));
  nor002aa1n20x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nanp02aa1n24x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  norb02aa1n06x4               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  xnbna2aa1n03x5               g119(.a(new_n214), .b(new_n211), .c(new_n203), .out0(\s[18] ));
  and002aa1n02x5               g120(.a(new_n199), .b(new_n214), .o(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n217));
  oaoi03aa1n02x5               g122(.a(\a[18] ), .b(\b[17] ), .c(new_n203), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  nor042aa1d18x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nand42aa1n10x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n12x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n217), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n06x5               g129(.a(new_n222), .b(new_n218), .c(new_n198), .d(new_n216), .o1(new_n225));
  nor042aa1n06x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  nand42aa1d28x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n227), .b(new_n226), .out0(new_n228));
  inv000aa1d42x5               g133(.a(\a[19] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\b[18] ), .o1(new_n230));
  aboi22aa1n03x5               g135(.a(new_n226), .b(new_n227), .c(new_n229), .d(new_n230), .out0(new_n231));
  inv030aa1n08x5               g136(.a(new_n220), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n222), .o1(new_n233));
  aoai13aa1n02x5               g138(.a(new_n232), .b(new_n233), .c(new_n217), .d(new_n219), .o1(new_n234));
  aoi022aa1n03x5               g139(.a(new_n234), .b(new_n228), .c(new_n225), .d(new_n231), .o1(\s[20] ));
  nano32aa1n03x7               g140(.a(new_n233), .b(new_n199), .c(new_n228), .d(new_n214), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n237));
  nanb03aa1n12x5               g142(.a(new_n226), .b(new_n227), .c(new_n221), .out0(new_n238));
  nor042aa1n06x5               g143(.a(\b[16] ), .b(\a[17] ), .o1(new_n239));
  oai112aa1n06x5               g144(.a(new_n232), .b(new_n213), .c(new_n212), .d(new_n239), .o1(new_n240));
  aoi012aa1n12x5               g145(.a(new_n226), .b(new_n220), .c(new_n227), .o1(new_n241));
  oai012aa1d24x5               g146(.a(new_n241), .b(new_n240), .c(new_n238), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  nor042aa1d18x5               g148(.a(\b[20] ), .b(\a[21] ), .o1(new_n244));
  nand42aa1n16x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  norb02aa1n03x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  xnbna2aa1n03x5               g151(.a(new_n246), .b(new_n237), .c(new_n243), .out0(\s[21] ));
  aoai13aa1n03x5               g152(.a(new_n246), .b(new_n242), .c(new_n198), .d(new_n236), .o1(new_n248));
  nor042aa1n09x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  nand42aa1d28x5               g154(.a(\b[21] ), .b(\a[22] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n250), .b(new_n249), .out0(new_n251));
  aoib12aa1n02x5               g156(.a(new_n244), .b(new_n250), .c(new_n249), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n244), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n246), .o1(new_n254));
  aoai13aa1n02x5               g159(.a(new_n253), .b(new_n254), .c(new_n237), .d(new_n243), .o1(new_n255));
  aoi022aa1n03x5               g160(.a(new_n255), .b(new_n251), .c(new_n248), .d(new_n252), .o1(\s[22] ));
  inv020aa1n02x5               g161(.a(new_n236), .o1(new_n257));
  nano22aa1n03x7               g162(.a(new_n257), .b(new_n246), .c(new_n251), .out0(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n259));
  nano23aa1d15x5               g164(.a(new_n244), .b(new_n249), .c(new_n250), .d(new_n245), .out0(new_n260));
  aoi012aa1d24x5               g165(.a(new_n249), .b(new_n244), .c(new_n250), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoi012aa1d18x5               g167(.a(new_n262), .b(new_n242), .c(new_n260), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(new_n259), .b(new_n263), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[23] ), .b(\b[22] ), .out0(new_n265));
  aoi112aa1n02x5               g170(.a(new_n265), .b(new_n262), .c(new_n242), .d(new_n260), .o1(new_n266));
  aoi022aa1n02x5               g171(.a(new_n264), .b(new_n265), .c(new_n259), .d(new_n266), .o1(\s[23] ));
  inv000aa1d42x5               g172(.a(new_n263), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n265), .b(new_n268), .c(new_n198), .d(new_n258), .o1(new_n269));
  tech160nm_fixorc02aa1n02p5x5 g174(.a(\a[24] ), .b(\b[23] ), .out0(new_n270));
  nor042aa1n09x5               g175(.a(\b[22] ), .b(\a[23] ), .o1(new_n271));
  norp02aa1n02x5               g176(.a(new_n270), .b(new_n271), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n265), .o1(new_n274));
  aoai13aa1n04x5               g179(.a(new_n273), .b(new_n274), .c(new_n259), .d(new_n263), .o1(new_n275));
  aoi022aa1n02x7               g180(.a(new_n275), .b(new_n270), .c(new_n269), .d(new_n272), .o1(\s[24] ));
  and002aa1n12x5               g181(.a(new_n270), .b(new_n265), .o(new_n277));
  nano22aa1n03x7               g182(.a(new_n257), .b(new_n277), .c(new_n260), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n279));
  nano22aa1n02x4               g184(.a(new_n226), .b(new_n221), .c(new_n227), .out0(new_n280));
  tech160nm_fioai012aa1n03p5x5 g185(.a(new_n213), .b(\b[18] ), .c(\a[19] ), .o1(new_n281));
  oab012aa1n02x4               g186(.a(new_n281), .b(new_n239), .c(new_n212), .out0(new_n282));
  inv020aa1n03x5               g187(.a(new_n241), .o1(new_n283));
  aoai13aa1n04x5               g188(.a(new_n260), .b(new_n283), .c(new_n282), .d(new_n280), .o1(new_n284));
  inv000aa1n06x5               g189(.a(new_n277), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[24] ), .b(\b[23] ), .c(new_n273), .carry(new_n286));
  aoai13aa1n12x5               g191(.a(new_n286), .b(new_n285), .c(new_n284), .d(new_n261), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(new_n279), .b(new_n288), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[25] ), .b(\b[24] ), .out0(new_n290));
  aoai13aa1n06x5               g195(.a(new_n277), .b(new_n262), .c(new_n242), .d(new_n260), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n290), .o1(new_n292));
  and003aa1n02x5               g197(.a(new_n291), .b(new_n292), .c(new_n286), .o(new_n293));
  aoi022aa1n02x5               g198(.a(new_n289), .b(new_n290), .c(new_n279), .d(new_n293), .o1(\s[25] ));
  aoai13aa1n03x5               g199(.a(new_n290), .b(new_n287), .c(new_n198), .d(new_n278), .o1(new_n295));
  tech160nm_fixorc02aa1n02p5x5 g200(.a(\a[26] ), .b(\b[25] ), .out0(new_n296));
  nor042aa1n06x5               g201(.a(\b[24] ), .b(\a[25] ), .o1(new_n297));
  norp02aa1n02x5               g202(.a(new_n296), .b(new_n297), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n297), .o1(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n292), .c(new_n279), .d(new_n288), .o1(new_n300));
  aoi022aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n298), .o1(\s[26] ));
  and002aa1n12x5               g206(.a(new_n296), .b(new_n290), .o(new_n302));
  nano32aa1n03x7               g207(.a(new_n257), .b(new_n302), .c(new_n260), .d(new_n277), .out0(new_n303));
  aoai13aa1n06x5               g208(.a(new_n303), .b(new_n210), .c(new_n128), .d(new_n194), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[26] ), .b(\b[25] ), .c(new_n299), .carry(new_n305));
  inv000aa1d42x5               g210(.a(new_n305), .o1(new_n306));
  aoi012aa1d18x5               g211(.a(new_n306), .b(new_n287), .c(new_n302), .o1(new_n307));
  nanp02aa1n02x5               g212(.a(new_n304), .b(new_n307), .o1(new_n308));
  xorc02aa1n12x5               g213(.a(\a[27] ), .b(\b[26] ), .out0(new_n309));
  aoi112aa1n02x5               g214(.a(new_n309), .b(new_n306), .c(new_n287), .d(new_n302), .o1(new_n310));
  aoi022aa1n02x7               g215(.a(new_n308), .b(new_n309), .c(new_n304), .d(new_n310), .o1(\s[27] ));
  inv000aa1d42x5               g216(.a(new_n302), .o1(new_n312));
  aoai13aa1n04x5               g217(.a(new_n305), .b(new_n312), .c(new_n291), .d(new_n286), .o1(new_n313));
  aoai13aa1n02x5               g218(.a(new_n309), .b(new_n313), .c(new_n198), .d(new_n303), .o1(new_n314));
  tech160nm_fixorc02aa1n03p5x5 g219(.a(\a[28] ), .b(\b[27] ), .out0(new_n315));
  norp02aa1n02x5               g220(.a(\b[26] ), .b(\a[27] ), .o1(new_n316));
  norp02aa1n02x5               g221(.a(new_n315), .b(new_n316), .o1(new_n317));
  inv000aa1n03x5               g222(.a(new_n316), .o1(new_n318));
  inv000aa1n02x5               g223(.a(new_n309), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n318), .b(new_n319), .c(new_n304), .d(new_n307), .o1(new_n320));
  aoi022aa1n03x5               g225(.a(new_n320), .b(new_n315), .c(new_n314), .d(new_n317), .o1(\s[28] ));
  and002aa1n02x5               g226(.a(new_n315), .b(new_n309), .o(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n313), .c(new_n198), .d(new_n303), .o1(new_n323));
  tech160nm_fixorc02aa1n02p5x5 g228(.a(\a[29] ), .b(\b[28] ), .out0(new_n324));
  oao003aa1n02x5               g229(.a(\a[28] ), .b(\b[27] ), .c(new_n318), .carry(new_n325));
  norb02aa1n02x5               g230(.a(new_n325), .b(new_n324), .out0(new_n326));
  inv000aa1d42x5               g231(.a(new_n322), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n325), .b(new_n327), .c(new_n304), .d(new_n307), .o1(new_n328));
  aoi022aa1n03x5               g233(.a(new_n328), .b(new_n324), .c(new_n323), .d(new_n326), .o1(\s[29] ));
  xorb03aa1n02x5               g234(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g235(.a(new_n319), .b(new_n315), .c(new_n324), .out0(new_n331));
  aoai13aa1n02x5               g236(.a(new_n331), .b(new_n313), .c(new_n198), .d(new_n303), .o1(new_n332));
  xorc02aa1n02x5               g237(.a(\a[30] ), .b(\b[29] ), .out0(new_n333));
  oao003aa1n02x5               g238(.a(\a[29] ), .b(\b[28] ), .c(new_n325), .carry(new_n334));
  norb02aa1n02x5               g239(.a(new_n334), .b(new_n333), .out0(new_n335));
  inv000aa1d42x5               g240(.a(new_n331), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n334), .b(new_n336), .c(new_n304), .d(new_n307), .o1(new_n337));
  aoi022aa1n03x5               g242(.a(new_n337), .b(new_n333), .c(new_n332), .d(new_n335), .o1(\s[30] ));
  nano32aa1n06x5               g243(.a(new_n319), .b(new_n333), .c(new_n315), .d(new_n324), .out0(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n313), .c(new_n198), .d(new_n303), .o1(new_n340));
  xorc02aa1n02x5               g245(.a(\a[31] ), .b(\b[30] ), .out0(new_n341));
  and002aa1n02x5               g246(.a(\b[29] ), .b(\a[30] ), .o(new_n342));
  oabi12aa1n02x5               g247(.a(new_n341), .b(\a[30] ), .c(\b[29] ), .out0(new_n343));
  oab012aa1n02x4               g248(.a(new_n343), .b(new_n334), .c(new_n342), .out0(new_n344));
  inv000aa1d42x5               g249(.a(new_n339), .o1(new_n345));
  oao003aa1n02x5               g250(.a(\a[30] ), .b(\b[29] ), .c(new_n334), .carry(new_n346));
  aoai13aa1n03x5               g251(.a(new_n346), .b(new_n345), .c(new_n304), .d(new_n307), .o1(new_n347));
  aoi022aa1n03x5               g252(.a(new_n347), .b(new_n341), .c(new_n340), .d(new_n344), .o1(\s[31] ));
  oai012aa1n02x5               g253(.a(new_n102), .b(new_n107), .c(new_n106), .o1(new_n349));
  xnrb03aa1n02x5               g254(.a(new_n349), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g255(.a(\a[3] ), .b(\b[2] ), .c(new_n349), .o1(new_n351));
  xorb03aa1n02x5               g256(.a(new_n351), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  aoi113aa1n02x5               g257(.a(new_n112), .b(new_n135), .c(new_n108), .d(new_n105), .e(new_n101), .o1(new_n353));
  aoi012aa1n02x5               g258(.a(new_n353), .b(new_n134), .c(new_n135), .o1(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g259(.a(\a[5] ), .b(\b[4] ), .c(new_n113), .o1(new_n355));
  xorb03aa1n02x5               g260(.a(new_n355), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g261(.a(new_n116), .b(new_n119), .c(new_n355), .d(new_n118), .o1(new_n357));
  aoi112aa1n02x5               g262(.a(new_n119), .b(new_n116), .c(new_n355), .d(new_n118), .o1(new_n358));
  norb02aa1n02x5               g263(.a(new_n357), .b(new_n358), .out0(\s[7] ));
  inv000aa1d42x5               g264(.a(new_n114), .o1(new_n360));
  xnbna2aa1n03x5               g265(.a(new_n121), .b(new_n357), .c(new_n360), .out0(\s[8] ));
  xorb03aa1n02x5               g266(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


