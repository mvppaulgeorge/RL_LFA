// Benchmark "adder" written by ABC on Thu Jul 18 11:18:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n343, new_n345,
    new_n348, new_n349, new_n350, new_n351, new_n353, new_n355, new_n356,
    new_n357, new_n359, new_n360, new_n361;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\a[9] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\b[8] ), .b(new_n98), .out0(new_n99));
  inv000aa1d42x5               g004(.a(\a[2] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[1] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  tech160nm_finand02aa1n05x5   g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  aob012aa1n06x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .out0(new_n105));
  nor042aa1n03x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nand42aa1n04x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  norb02aa1n03x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  norp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nand42aa1n03x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  norb02aa1n06x4               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  nanp03aa1n09x5               g016(.a(new_n105), .b(new_n108), .c(new_n111), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[3] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[2] ), .o1(new_n114));
  aoai13aa1n09x5               g019(.a(new_n107), .b(new_n106), .c(new_n113), .d(new_n114), .o1(new_n115));
  nor042aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  norb02aa1n06x5               g022(.a(new_n117), .b(new_n116), .out0(new_n118));
  xorc02aa1n12x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nand02aa1n04x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nor002aa1n20x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nor042aa1n06x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  nand02aa1n04x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  nano23aa1n06x5               g028(.a(new_n122), .b(new_n121), .c(new_n123), .d(new_n120), .out0(new_n124));
  nand03aa1n03x5               g029(.a(new_n124), .b(new_n118), .c(new_n119), .o1(new_n125));
  nanb03aa1n03x5               g030(.a(new_n116), .b(new_n123), .c(new_n117), .out0(new_n126));
  nor042aa1n02x5               g031(.a(\b[4] ), .b(\a[5] ), .o1(new_n127));
  inv000aa1n02x5               g032(.a(new_n122), .o1(new_n128));
  aoai13aa1n04x5               g033(.a(new_n128), .b(new_n121), .c(new_n127), .d(new_n120), .o1(new_n129));
  aoi012aa1n06x5               g034(.a(new_n122), .b(new_n116), .c(new_n123), .o1(new_n130));
  inv000aa1n02x5               g035(.a(new_n130), .o1(new_n131));
  oab012aa1n06x5               g036(.a(new_n131), .b(new_n129), .c(new_n126), .out0(new_n132));
  aoai13aa1n12x5               g037(.a(new_n132), .b(new_n125), .c(new_n112), .d(new_n115), .o1(new_n133));
  tech160nm_fixorc02aa1n02p5x5 g038(.a(\a[9] ), .b(\b[8] ), .out0(new_n134));
  nand22aa1n03x5               g039(.a(new_n133), .b(new_n134), .o1(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n97), .b(new_n135), .c(new_n99), .out0(\s[10] ));
  nanp02aa1n02x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nand42aa1n06x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norp02aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  oa0022aa1n03x5               g045(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n141));
  nanp02aa1n03x5               g046(.a(new_n135), .b(new_n141), .o1(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n140), .b(new_n142), .c(new_n137), .out0(\s[11] ));
  nano22aa1n02x4               g048(.a(new_n139), .b(new_n137), .c(new_n138), .out0(new_n144));
  tech160nm_fiaoi012aa1n05x5   g049(.a(new_n139), .b(new_n142), .c(new_n144), .o1(new_n145));
  xnrb03aa1n03x5               g050(.a(new_n145), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n03x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand42aa1n08x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nano23aa1n02x5               g053(.a(new_n147), .b(new_n139), .c(new_n148), .d(new_n138), .out0(new_n149));
  and003aa1n02x5               g054(.a(new_n149), .b(new_n134), .c(new_n97), .o(new_n150));
  nand22aa1n03x5               g055(.a(new_n133), .b(new_n150), .o1(new_n151));
  nano22aa1n03x7               g056(.a(new_n147), .b(new_n138), .c(new_n148), .out0(new_n152));
  nona23aa1d18x5               g057(.a(new_n152), .b(new_n137), .c(new_n141), .d(new_n139), .out0(new_n153));
  aoi012aa1d18x5               g058(.a(new_n147), .b(new_n139), .c(new_n148), .o1(new_n154));
  nand02aa1d06x5               g059(.a(new_n153), .b(new_n154), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nanp02aa1n03x5               g061(.a(new_n151), .b(new_n156), .o1(new_n157));
  xorc02aa1n12x5               g062(.a(\a[13] ), .b(\b[12] ), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  and003aa1n02x5               g064(.a(new_n153), .b(new_n159), .c(new_n154), .o(new_n160));
  aoi022aa1n02x5               g065(.a(new_n157), .b(new_n158), .c(new_n151), .d(new_n160), .o1(\s[13] ));
  inv000aa1d42x5               g066(.a(\a[14] ), .o1(new_n162));
  norp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  tech160nm_fiaoi012aa1n05x5   g068(.a(new_n163), .b(new_n157), .c(new_n158), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(new_n162), .out0(\s[14] ));
  tech160nm_fixorc02aa1n04x5   g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  and002aa1n02x5               g071(.a(new_n166), .b(new_n158), .o(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n155), .c(new_n133), .d(new_n150), .o1(new_n168));
  inv000aa1d42x5               g073(.a(\b[13] ), .o1(new_n169));
  oao003aa1n02x5               g074(.a(new_n162), .b(new_n169), .c(new_n163), .carry(new_n170));
  nanb02aa1n02x5               g075(.a(new_n170), .b(new_n168), .out0(new_n171));
  norp02aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  oai022aa1n02x5               g079(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n175));
  oaoi13aa1n02x5               g080(.a(new_n174), .b(new_n175), .c(new_n162), .d(new_n169), .o1(new_n176));
  aoi022aa1n02x5               g081(.a(new_n171), .b(new_n174), .c(new_n168), .d(new_n176), .o1(\s[15] ));
  nor042aa1n02x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand42aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n03x5               g085(.a(new_n180), .b(new_n172), .c(new_n171), .d(new_n173), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n174), .b(new_n170), .c(new_n157), .d(new_n167), .o1(new_n182));
  nona22aa1n02x4               g087(.a(new_n182), .b(new_n180), .c(new_n172), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n181), .b(new_n183), .o1(\s[16] ));
  nano23aa1n06x5               g089(.a(new_n172), .b(new_n178), .c(new_n179), .d(new_n173), .out0(new_n185));
  nand23aa1d12x5               g090(.a(new_n185), .b(new_n158), .c(new_n166), .o1(new_n186));
  nano32aa1d12x5               g091(.a(new_n186), .b(new_n149), .c(new_n134), .d(new_n97), .out0(new_n187));
  nanp02aa1n06x5               g092(.a(new_n133), .b(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n186), .o1(new_n189));
  nanb03aa1n02x5               g094(.a(new_n178), .b(new_n179), .c(new_n173), .out0(new_n190));
  oai122aa1n02x7               g095(.a(new_n175), .b(\a[15] ), .c(\b[14] ), .d(new_n162), .e(new_n169), .o1(new_n191));
  aoi012aa1n02x5               g096(.a(new_n178), .b(new_n172), .c(new_n179), .o1(new_n192));
  oa0012aa1n06x5               g097(.a(new_n192), .b(new_n191), .c(new_n190), .o(new_n193));
  aobi12aa1n06x5               g098(.a(new_n193), .b(new_n155), .c(new_n189), .out0(new_n194));
  nand02aa1d10x5               g099(.a(new_n188), .b(new_n194), .o1(new_n195));
  xorc02aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  norb02aa1n02x5               g101(.a(new_n192), .b(new_n196), .out0(new_n197));
  oai012aa1n02x5               g102(.a(new_n197), .b(new_n191), .c(new_n190), .o1(new_n198));
  aoi012aa1n02x5               g103(.a(new_n198), .b(new_n155), .c(new_n189), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n195), .b(new_n196), .c(new_n188), .d(new_n199), .o1(\s[17] ));
  inv040aa1d32x5               g105(.a(\a[18] ), .o1(new_n201));
  nor022aa1n04x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  tech160nm_fiaoi012aa1n05x5   g107(.a(new_n202), .b(new_n195), .c(new_n196), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[17] ), .c(new_n201), .out0(\s[18] ));
  aoai13aa1n12x5               g109(.a(new_n193), .b(new_n186), .c(new_n153), .d(new_n154), .o1(new_n205));
  inv000aa1d42x5               g110(.a(\a[17] ), .o1(new_n206));
  xroi22aa1d06x4               g111(.a(new_n206), .b(\b[16] ), .c(new_n201), .d(\b[17] ), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n205), .c(new_n133), .d(new_n187), .o1(new_n208));
  nand42aa1n02x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  oab012aa1n02x4               g114(.a(new_n202), .b(\a[18] ), .c(\b[17] ), .out0(new_n210));
  norb02aa1n02x5               g115(.a(new_n209), .b(new_n210), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor022aa1n04x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nanp02aa1n04x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n06x4               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n208), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n06x5               g122(.a(new_n208), .b(new_n212), .o1(new_n218));
  nor042aa1n04x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand42aa1n06x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nanb02aa1n02x5               g125(.a(new_n219), .b(new_n220), .out0(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n213), .c(new_n218), .d(new_n214), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(new_n218), .b(new_n215), .o1(new_n223));
  nona22aa1n02x4               g128(.a(new_n223), .b(new_n221), .c(new_n213), .out0(new_n224));
  nanp02aa1n02x5               g129(.a(new_n224), .b(new_n222), .o1(\s[20] ));
  nanb03aa1d18x5               g130(.a(new_n221), .b(new_n207), .c(new_n215), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n205), .c(new_n133), .d(new_n187), .o1(new_n228));
  nanb03aa1n02x5               g133(.a(new_n219), .b(new_n220), .c(new_n214), .out0(new_n229));
  oai022aa1n02x5               g134(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n230));
  oai112aa1n02x5               g135(.a(new_n230), .b(new_n209), .c(\b[18] ), .d(\a[19] ), .o1(new_n231));
  aoi012aa1n12x5               g136(.a(new_n219), .b(new_n213), .c(new_n220), .o1(new_n232));
  tech160nm_fioai012aa1n03p5x5 g137(.a(new_n232), .b(new_n231), .c(new_n229), .o1(new_n233));
  nanb02aa1n03x5               g138(.a(new_n233), .b(new_n228), .out0(new_n234));
  tech160nm_fixorc02aa1n03p5x5 g139(.a(\a[21] ), .b(\b[20] ), .out0(new_n235));
  nano22aa1n02x4               g140(.a(new_n219), .b(new_n214), .c(new_n220), .out0(new_n236));
  oai012aa1n02x5               g141(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .o1(new_n237));
  norp02aa1n02x5               g142(.a(new_n210), .b(new_n237), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n232), .o1(new_n239));
  aoi112aa1n02x5               g144(.a(new_n239), .b(new_n235), .c(new_n238), .d(new_n236), .o1(new_n240));
  aoi022aa1n02x5               g145(.a(new_n234), .b(new_n235), .c(new_n228), .d(new_n240), .o1(\s[21] ));
  nor042aa1n03x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  tech160nm_fixnrc02aa1n05x5   g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n242), .c(new_n234), .d(new_n235), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n235), .b(new_n233), .c(new_n195), .d(new_n227), .o1(new_n245));
  nona22aa1n03x5               g150(.a(new_n245), .b(new_n243), .c(new_n242), .out0(new_n246));
  nanp02aa1n03x5               g151(.a(new_n244), .b(new_n246), .o1(\s[22] ));
  xnrc02aa1n02x5               g152(.a(\b[20] ), .b(\a[21] ), .out0(new_n248));
  nor002aa1n03x5               g153(.a(new_n243), .b(new_n248), .o1(new_n249));
  nano32aa1n02x5               g154(.a(new_n221), .b(new_n207), .c(new_n249), .d(new_n215), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n205), .c(new_n133), .d(new_n187), .o1(new_n251));
  nona22aa1n02x4               g156(.a(new_n236), .b(new_n210), .c(new_n237), .out0(new_n252));
  nanb02aa1n03x5               g157(.a(new_n243), .b(new_n235), .out0(new_n253));
  inv000aa1d42x5               g158(.a(\a[22] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\b[21] ), .o1(new_n255));
  oao003aa1n06x5               g160(.a(new_n254), .b(new_n255), .c(new_n242), .carry(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  aoai13aa1n02x5               g162(.a(new_n257), .b(new_n253), .c(new_n252), .d(new_n232), .o1(new_n258));
  nanb02aa1n03x5               g163(.a(new_n258), .b(new_n251), .out0(new_n259));
  xorc02aa1n12x5               g164(.a(\a[23] ), .b(\b[22] ), .out0(new_n260));
  aoi112aa1n02x5               g165(.a(new_n260), .b(new_n256), .c(new_n233), .d(new_n249), .o1(new_n261));
  aoi022aa1n02x5               g166(.a(new_n259), .b(new_n260), .c(new_n251), .d(new_n261), .o1(\s[23] ));
  nor002aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  tech160nm_fixnrc02aa1n04x5   g168(.a(\b[23] ), .b(\a[24] ), .out0(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n263), .c(new_n259), .d(new_n260), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n260), .b(new_n258), .c(new_n195), .d(new_n250), .o1(new_n266));
  nona22aa1n03x5               g171(.a(new_n266), .b(new_n264), .c(new_n263), .out0(new_n267));
  nanp02aa1n03x5               g172(.a(new_n265), .b(new_n267), .o1(\s[24] ));
  norb02aa1n06x5               g173(.a(new_n260), .b(new_n264), .out0(new_n269));
  nano22aa1n03x7               g174(.a(new_n226), .b(new_n249), .c(new_n269), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n205), .c(new_n133), .d(new_n187), .o1(new_n271));
  aoai13aa1n03x5               g176(.a(new_n249), .b(new_n239), .c(new_n238), .d(new_n236), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n269), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\a[24] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(\b[23] ), .o1(new_n275));
  oao003aa1n02x5               g180(.a(new_n274), .b(new_n275), .c(new_n263), .carry(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n273), .c(new_n272), .d(new_n257), .o1(new_n278));
  nanb02aa1n06x5               g183(.a(new_n278), .b(new_n271), .out0(new_n279));
  xorc02aa1n12x5               g184(.a(\a[25] ), .b(\b[24] ), .out0(new_n280));
  aoi112aa1n02x5               g185(.a(new_n280), .b(new_n276), .c(new_n258), .d(new_n269), .o1(new_n281));
  aoi022aa1n02x5               g186(.a(new_n279), .b(new_n280), .c(new_n271), .d(new_n281), .o1(\s[25] ));
  norp02aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  tech160nm_fixnrc02aa1n04x5   g188(.a(\b[25] ), .b(\a[26] ), .out0(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n283), .c(new_n279), .d(new_n280), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n280), .b(new_n278), .c(new_n195), .d(new_n270), .o1(new_n286));
  nona22aa1n03x5               g191(.a(new_n286), .b(new_n284), .c(new_n283), .out0(new_n287));
  nanp02aa1n02x5               g192(.a(new_n285), .b(new_n287), .o1(\s[26] ));
  norb02aa1n03x5               g193(.a(new_n280), .b(new_n284), .out0(new_n289));
  nano32aa1n03x7               g194(.a(new_n226), .b(new_n289), .c(new_n249), .d(new_n269), .out0(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n205), .c(new_n133), .d(new_n187), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\a[26] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\b[25] ), .o1(new_n293));
  oao003aa1n02x5               g198(.a(new_n292), .b(new_n293), .c(new_n283), .carry(new_n294));
  aoi012aa1n03x5               g199(.a(new_n294), .b(new_n278), .c(new_n289), .o1(new_n295));
  tech160nm_fixorc02aa1n05x5   g200(.a(\a[27] ), .b(\b[26] ), .out0(new_n296));
  xnbna2aa1n03x5               g201(.a(new_n296), .b(new_n295), .c(new_n291), .out0(\s[27] ));
  aoai13aa1n02x5               g202(.a(new_n289), .b(new_n276), .c(new_n258), .d(new_n269), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n294), .o1(new_n299));
  nanp03aa1n06x5               g204(.a(new_n291), .b(new_n298), .c(new_n299), .o1(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  norp02aa1n02x5               g206(.a(\b[27] ), .b(\a[28] ), .o1(new_n302));
  nanp02aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .o1(new_n303));
  nanb02aa1n02x5               g208(.a(new_n302), .b(new_n303), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n300), .d(new_n296), .o1(new_n305));
  aoai13aa1n02x5               g210(.a(new_n269), .b(new_n256), .c(new_n233), .d(new_n249), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n289), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n299), .b(new_n307), .c(new_n306), .d(new_n277), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n296), .b(new_n308), .c(new_n195), .d(new_n290), .o1(new_n309));
  nona22aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n301), .out0(new_n310));
  nanp02aa1n03x5               g215(.a(new_n305), .b(new_n310), .o1(\s[28] ));
  norb02aa1n09x5               g216(.a(new_n296), .b(new_n304), .out0(new_n312));
  aoai13aa1n02x5               g217(.a(new_n312), .b(new_n308), .c(new_n195), .d(new_n290), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .out0(new_n314));
  aoi012aa1n02x5               g219(.a(new_n302), .b(new_n301), .c(new_n303), .o1(new_n315));
  norb02aa1n02x5               g220(.a(new_n315), .b(new_n314), .out0(new_n316));
  inv000aa1d42x5               g221(.a(new_n312), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n315), .b(new_n317), .c(new_n295), .d(new_n291), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n313), .d(new_n316), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g225(.a(new_n304), .b(new_n314), .c(new_n296), .out0(new_n321));
  nanb02aa1n03x5               g226(.a(new_n321), .b(new_n300), .out0(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  inv000aa1d42x5               g228(.a(\a[29] ), .o1(new_n324));
  inv000aa1d42x5               g229(.a(\b[28] ), .o1(new_n325));
  oaib12aa1n02x5               g230(.a(new_n315), .b(\b[28] ), .c(new_n324), .out0(new_n326));
  oaoi13aa1n02x5               g231(.a(new_n323), .b(new_n326), .c(new_n324), .d(new_n325), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n326), .b(new_n325), .c(\a[29] ), .out0(new_n328));
  aoai13aa1n02x7               g233(.a(new_n328), .b(new_n321), .c(new_n295), .d(new_n291), .o1(new_n329));
  aoi022aa1n03x5               g234(.a(new_n329), .b(new_n323), .c(new_n322), .d(new_n327), .o1(\s[30] ));
  nano22aa1n06x5               g235(.a(new_n317), .b(new_n314), .c(new_n323), .out0(new_n331));
  aoai13aa1n03x5               g236(.a(new_n331), .b(new_n308), .c(new_n195), .d(new_n290), .o1(new_n332));
  aoi022aa1n02x5               g237(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n333));
  norb02aa1n02x5               g238(.a(\b[30] ), .b(\a[31] ), .out0(new_n334));
  obai22aa1n02x7               g239(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n335));
  aoi112aa1n02x5               g240(.a(new_n335), .b(new_n334), .c(new_n326), .d(new_n333), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n331), .o1(new_n337));
  norp02aa1n02x5               g242(.a(\b[29] ), .b(\a[30] ), .o1(new_n338));
  aoi012aa1n02x5               g243(.a(new_n338), .b(new_n326), .c(new_n333), .o1(new_n339));
  aoai13aa1n02x7               g244(.a(new_n339), .b(new_n337), .c(new_n295), .d(new_n291), .o1(new_n340));
  xorc02aa1n02x5               g245(.a(\a[31] ), .b(\b[30] ), .out0(new_n341));
  aoi022aa1n02x7               g246(.a(new_n340), .b(new_n341), .c(new_n336), .d(new_n332), .o1(\s[31] ));
  nanp03aa1n02x5               g247(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n111), .b(new_n343), .c(new_n102), .out0(\s[3] ));
  oaoi03aa1n02x5               g249(.a(new_n113), .b(new_n114), .c(new_n105), .o1(new_n345));
  xnrc02aa1n02x5               g250(.a(new_n345), .b(new_n108), .out0(\s[4] ));
  xnbna2aa1n03x5               g251(.a(new_n119), .b(new_n112), .c(new_n115), .out0(\s[5] ));
  nanp02aa1n02x5               g252(.a(new_n112), .b(new_n115), .o1(new_n348));
  norb02aa1n02x5               g253(.a(new_n120), .b(new_n121), .out0(new_n349));
  aoai13aa1n03x5               g254(.a(new_n349), .b(new_n127), .c(new_n348), .d(new_n119), .o1(new_n350));
  aoi112aa1n02x5               g255(.a(new_n127), .b(new_n349), .c(new_n348), .d(new_n119), .o1(new_n351));
  norb02aa1n02x5               g256(.a(new_n350), .b(new_n351), .out0(\s[6] ));
  inv000aa1d42x5               g257(.a(new_n121), .o1(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n118), .b(new_n350), .c(new_n353), .out0(\s[7] ));
  orn002aa1n02x5               g259(.a(\a[7] ), .b(\b[6] ), .o(new_n355));
  norb02aa1n02x5               g260(.a(new_n123), .b(new_n122), .out0(new_n356));
  aob012aa1n02x5               g261(.a(new_n118), .b(new_n350), .c(new_n353), .out0(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n356), .b(new_n357), .c(new_n355), .out0(\s[8] ));
  aoi012aa1n02x5               g263(.a(new_n125), .b(new_n112), .c(new_n115), .o1(new_n359));
  norp02aa1n02x5               g264(.a(new_n129), .b(new_n126), .o1(new_n360));
  norp03aa1n02x5               g265(.a(new_n360), .b(new_n131), .c(new_n134), .o1(new_n361));
  aboi22aa1n03x5               g266(.a(new_n359), .b(new_n361), .c(new_n133), .d(new_n134), .out0(\s[9] ));
endmodule


