// Benchmark "adder" written by ABC on Wed Jul 17 18:47:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n355, new_n357, new_n358, new_n360,
    new_n362, new_n363, new_n364, new_n366, new_n367, new_n369, new_n370,
    new_n371, new_n373;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[8] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\a[9] ), .b(new_n97), .out0(new_n98));
  norp02aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aob012aa1n06x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  nor002aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n06x4               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor042aa1n04x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanp02aa1n04x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n06x4               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nand23aa1n06x5               g014(.a(new_n103), .b(new_n106), .c(new_n109), .o1(new_n110));
  tech160nm_fiaoi012aa1n05x5   g015(.a(new_n104), .b(new_n107), .c(new_n105), .o1(new_n111));
  nor042aa1n12x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand42aa1n10x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor042aa1n03x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand02aa1d04x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nor042aa1n03x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand02aa1d24x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nor002aa1n12x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nanp02aa1n12x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nano23aa1n02x5               g025(.a(new_n117), .b(new_n119), .c(new_n120), .d(new_n118), .out0(new_n121));
  nand02aa1n02x5               g026(.a(new_n121), .b(new_n116), .o1(new_n122));
  norb02aa1n06x4               g027(.a(new_n118), .b(new_n117), .out0(new_n123));
  nano22aa1n03x7               g028(.a(new_n119), .b(new_n113), .c(new_n120), .out0(new_n124));
  oai022aa1n03x5               g029(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n125));
  inv040aa1n02x5               g030(.a(new_n119), .o1(new_n126));
  oaoi03aa1n09x5               g031(.a(\a[8] ), .b(\b[7] ), .c(new_n126), .o1(new_n127));
  aoi013aa1n06x4               g032(.a(new_n127), .b(new_n124), .c(new_n125), .d(new_n123), .o1(new_n128));
  aoai13aa1n12x5               g033(.a(new_n128), .b(new_n122), .c(new_n110), .d(new_n111), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  nanp02aa1n02x5               g035(.a(new_n129), .b(new_n130), .o1(new_n131));
  xorc02aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n131), .c(new_n98), .out0(\s[10] ));
  and002aa1n02x5               g038(.a(new_n132), .b(new_n130), .o(new_n134));
  nanp02aa1n06x5               g039(.a(new_n129), .b(new_n134), .o1(new_n135));
  nanp02aa1n04x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  oai022aa1d24x5               g041(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n137));
  nanp02aa1n02x5               g042(.a(new_n137), .b(new_n136), .o1(new_n138));
  nor042aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1n04x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n135), .c(new_n138), .out0(\s[11] ));
  aob012aa1n03x5               g047(.a(new_n141), .b(new_n135), .c(new_n138), .out0(new_n143));
  nor042aa1n06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand02aa1d16x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  aoib12aa1n02x5               g051(.a(new_n139), .b(new_n145), .c(new_n144), .out0(new_n147));
  oai012aa1n03x5               g052(.a(new_n143), .b(\b[10] ), .c(\a[11] ), .o1(new_n148));
  aoi022aa1n03x5               g053(.a(new_n148), .b(new_n146), .c(new_n143), .d(new_n147), .o1(\s[12] ));
  nano23aa1n06x5               g054(.a(new_n139), .b(new_n144), .c(new_n145), .d(new_n140), .out0(new_n150));
  nand23aa1n06x5               g055(.a(new_n150), .b(new_n130), .c(new_n132), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(new_n129), .b(new_n152), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n99), .b(new_n101), .c(new_n102), .o1(new_n154));
  nona23aa1n02x4               g059(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n155));
  tech160nm_fioai012aa1n03p5x5 g060(.a(new_n111), .b(new_n155), .c(new_n154), .o1(new_n156));
  nanb02aa1n06x5               g061(.a(new_n122), .b(new_n156), .out0(new_n157));
  nano22aa1n09x5               g062(.a(new_n144), .b(new_n140), .c(new_n145), .out0(new_n158));
  oai112aa1n06x5               g063(.a(new_n137), .b(new_n136), .c(\b[10] ), .d(\a[11] ), .o1(new_n159));
  aoi012aa1d18x5               g064(.a(new_n144), .b(new_n139), .c(new_n145), .o1(new_n160));
  oaib12aa1n18x5               g065(.a(new_n160), .b(new_n159), .c(new_n158), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n151), .c(new_n157), .d(new_n128), .o1(new_n163));
  nor042aa1n04x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nand02aa1d04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  nanb02aa1n06x5               g071(.a(new_n159), .b(new_n158), .out0(new_n167));
  nano22aa1n02x4               g072(.a(new_n166), .b(new_n167), .c(new_n160), .out0(new_n168));
  aoi022aa1n02x5               g073(.a(new_n163), .b(new_n166), .c(new_n153), .d(new_n168), .o1(\s[13] ));
  orn002aa1n02x5               g074(.a(\a[13] ), .b(\b[12] ), .o(new_n170));
  aoai13aa1n03x5               g075(.a(new_n166), .b(new_n161), .c(new_n129), .d(new_n152), .o1(new_n171));
  nor022aa1n08x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nand02aa1d06x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n171), .c(new_n170), .out0(\s[14] ));
  nano23aa1n06x5               g080(.a(new_n164), .b(new_n172), .c(new_n173), .d(new_n165), .out0(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n161), .c(new_n129), .d(new_n152), .o1(new_n177));
  tech160nm_fioaoi03aa1n03p5x5 g082(.a(\a[14] ), .b(\b[13] ), .c(new_n170), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  nor042aa1d18x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  nanp02aa1n04x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  norb02aa1d21x5               g086(.a(new_n181), .b(new_n180), .out0(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n177), .c(new_n179), .out0(\s[15] ));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n178), .c(new_n163), .d(new_n176), .o1(new_n184));
  xorc02aa1n02x5               g089(.a(\a[16] ), .b(\b[15] ), .out0(new_n185));
  inv000aa1d42x5               g090(.a(\a[16] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[15] ), .o1(new_n187));
  nanp02aa1n02x5               g092(.a(new_n187), .b(new_n186), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  aoi012aa1n02x5               g094(.a(new_n180), .b(new_n188), .c(new_n189), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n180), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n182), .o1(new_n192));
  aoai13aa1n03x5               g097(.a(new_n191), .b(new_n192), .c(new_n177), .d(new_n179), .o1(new_n193));
  aoi022aa1n02x7               g098(.a(new_n193), .b(new_n185), .c(new_n184), .d(new_n190), .o1(\s[16] ));
  nand23aa1n04x5               g099(.a(new_n176), .b(new_n182), .c(new_n185), .o1(new_n195));
  nor042aa1n09x5               g100(.a(new_n195), .b(new_n151), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n129), .b(new_n196), .o1(new_n197));
  nona23aa1n02x4               g102(.a(new_n173), .b(new_n165), .c(new_n164), .d(new_n172), .out0(new_n198));
  nano32aa1n03x7               g103(.a(new_n198), .b(new_n189), .c(new_n182), .d(new_n188), .out0(new_n199));
  nand03aa1n02x5               g104(.a(new_n199), .b(new_n134), .c(new_n150), .o1(new_n200));
  nanp03aa1n02x5               g105(.a(new_n188), .b(new_n181), .c(new_n189), .o1(new_n201));
  oai112aa1n06x5               g106(.a(new_n191), .b(new_n173), .c(new_n172), .d(new_n164), .o1(new_n202));
  tech160nm_fioaoi03aa1n03p5x5 g107(.a(new_n186), .b(new_n187), .c(new_n180), .o1(new_n203));
  oai012aa1n06x5               g108(.a(new_n203), .b(new_n202), .c(new_n201), .o1(new_n204));
  tech160nm_fiaoi012aa1n05x5   g109(.a(new_n204), .b(new_n161), .c(new_n199), .o1(new_n205));
  aoai13aa1n04x5               g110(.a(new_n205), .b(new_n200), .c(new_n157), .d(new_n128), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[17] ), .b(\b[16] ), .out0(new_n207));
  norp02aa1n02x5               g112(.a(new_n202), .b(new_n201), .o1(new_n208));
  nanb02aa1n02x5               g113(.a(new_n207), .b(new_n203), .out0(new_n209));
  aoi112aa1n02x5               g114(.a(new_n209), .b(new_n208), .c(new_n161), .d(new_n199), .o1(new_n210));
  aoi022aa1n02x5               g115(.a(new_n206), .b(new_n207), .c(new_n197), .d(new_n210), .o1(\s[17] ));
  inv000aa1d42x5               g116(.a(\a[17] ), .o1(new_n212));
  nanb02aa1n02x5               g117(.a(\b[16] ), .b(new_n212), .out0(new_n213));
  inv000aa1n02x5               g118(.a(new_n204), .o1(new_n214));
  aoai13aa1n12x5               g119(.a(new_n214), .b(new_n195), .c(new_n167), .d(new_n160), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n207), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n216));
  xorc02aa1n02x5               g121(.a(\a[18] ), .b(\b[17] ), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n216), .c(new_n213), .out0(\s[18] ));
  inv000aa1d42x5               g123(.a(\a[18] ), .o1(new_n219));
  xroi22aa1d04x5               g124(.a(new_n212), .b(\b[16] ), .c(new_n219), .d(\b[17] ), .out0(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n221));
  oaoi03aa1n02x5               g126(.a(\a[18] ), .b(\b[17] ), .c(new_n213), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  nor002aa1n20x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  nand42aa1n04x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  norb02aa1n02x5               g130(.a(new_n225), .b(new_n224), .out0(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n221), .c(new_n223), .out0(\s[19] ));
  xnrc02aa1n02x5               g132(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g133(.a(new_n226), .b(new_n222), .c(new_n206), .d(new_n220), .o1(new_n229));
  nor042aa1n04x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nand42aa1n20x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(\a[19] ), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\b[18] ), .o1(new_n234));
  aboi22aa1n03x5               g139(.a(new_n230), .b(new_n231), .c(new_n233), .d(new_n234), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n224), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n226), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n237), .c(new_n221), .d(new_n223), .o1(new_n238));
  aoi022aa1n03x5               g143(.a(new_n238), .b(new_n232), .c(new_n229), .d(new_n235), .o1(\s[20] ));
  nano23aa1n02x5               g144(.a(new_n224), .b(new_n230), .c(new_n231), .d(new_n225), .out0(new_n240));
  and003aa1n02x5               g145(.a(new_n240), .b(new_n217), .c(new_n207), .o(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n242));
  oaih22aa1n04x5               g147(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n243));
  nano22aa1n03x7               g148(.a(new_n230), .b(new_n225), .c(new_n231), .out0(new_n244));
  aoi012aa1n09x5               g149(.a(new_n224), .b(\a[18] ), .c(\b[17] ), .o1(new_n245));
  nanp03aa1d12x5               g150(.a(new_n244), .b(new_n243), .c(new_n245), .o1(new_n246));
  aoi012aa1d18x5               g151(.a(new_n230), .b(new_n224), .c(new_n231), .o1(new_n247));
  nand22aa1n12x5               g152(.a(new_n246), .b(new_n247), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(new_n242), .b(new_n249), .o1(new_n250));
  nor042aa1d18x5               g155(.a(\b[20] ), .b(\a[21] ), .o1(new_n251));
  nand42aa1d28x5               g156(.a(\b[20] ), .b(\a[21] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  nanb03aa1n02x5               g158(.a(new_n230), .b(new_n231), .c(new_n225), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n254), .b(new_n245), .c(new_n243), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n253), .o1(new_n256));
  nano22aa1n02x4               g161(.a(new_n255), .b(new_n247), .c(new_n256), .out0(new_n257));
  aoi022aa1n02x5               g162(.a(new_n250), .b(new_n253), .c(new_n242), .d(new_n257), .o1(\s[21] ));
  aoai13aa1n03x5               g163(.a(new_n253), .b(new_n248), .c(new_n206), .d(new_n241), .o1(new_n259));
  nor042aa1n04x5               g164(.a(\b[21] ), .b(\a[22] ), .o1(new_n260));
  nand42aa1d28x5               g165(.a(\b[21] ), .b(\a[22] ), .o1(new_n261));
  norb02aa1n02x5               g166(.a(new_n261), .b(new_n260), .out0(new_n262));
  aoib12aa1n02x5               g167(.a(new_n251), .b(new_n261), .c(new_n260), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n251), .o1(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n256), .c(new_n242), .d(new_n249), .o1(new_n265));
  aoi022aa1n03x5               g170(.a(new_n265), .b(new_n262), .c(new_n259), .d(new_n263), .o1(\s[22] ));
  nano23aa1d15x5               g171(.a(new_n251), .b(new_n260), .c(new_n261), .d(new_n252), .out0(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  nano32aa1n02x4               g173(.a(new_n268), .b(new_n240), .c(new_n217), .d(new_n207), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n270));
  oai022aa1d24x5               g175(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n271));
  aoi022aa1n12x5               g176(.a(new_n248), .b(new_n267), .c(new_n261), .d(new_n271), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(new_n270), .b(new_n272), .o1(new_n273));
  nor002aa1n16x5               g178(.a(\b[22] ), .b(\a[23] ), .o1(new_n274));
  nand02aa1n03x5               g179(.a(\b[22] ), .b(\a[23] ), .o1(new_n275));
  norb02aa1n15x5               g180(.a(new_n275), .b(new_n274), .out0(new_n276));
  aoi122aa1n02x5               g181(.a(new_n276), .b(new_n261), .c(new_n271), .d(new_n248), .e(new_n267), .o1(new_n277));
  aoi022aa1n02x5               g182(.a(new_n273), .b(new_n276), .c(new_n270), .d(new_n277), .o1(\s[23] ));
  inv000aa1n02x5               g183(.a(new_n272), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n276), .b(new_n279), .c(new_n206), .d(new_n269), .o1(new_n280));
  tech160nm_fixorc02aa1n04x5   g185(.a(\a[24] ), .b(\b[23] ), .out0(new_n281));
  orn002aa1n02x7               g186(.a(\a[24] ), .b(\b[23] ), .o(new_n282));
  nanp02aa1n02x5               g187(.a(\b[23] ), .b(\a[24] ), .o1(new_n283));
  aoi012aa1n02x5               g188(.a(new_n274), .b(new_n282), .c(new_n283), .o1(new_n284));
  inv000aa1n02x5               g189(.a(new_n274), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n276), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n285), .b(new_n286), .c(new_n270), .d(new_n272), .o1(new_n287));
  aoi022aa1n03x5               g192(.a(new_n287), .b(new_n281), .c(new_n280), .d(new_n284), .o1(\s[24] ));
  nand23aa1d12x5               g193(.a(new_n267), .b(new_n276), .c(new_n281), .o1(new_n289));
  nano32aa1n02x4               g194(.a(new_n289), .b(new_n240), .c(new_n217), .d(new_n207), .out0(new_n290));
  aoai13aa1n04x5               g195(.a(new_n290), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n291));
  nanp03aa1n02x5               g196(.a(new_n282), .b(new_n275), .c(new_n283), .o1(new_n292));
  nano32aa1n02x4               g197(.a(new_n292), .b(new_n271), .c(new_n285), .d(new_n261), .out0(new_n293));
  aob012aa1n02x5               g198(.a(new_n282), .b(new_n274), .c(new_n283), .out0(new_n294));
  nor042aa1n04x5               g199(.a(new_n293), .b(new_n294), .o1(new_n295));
  aoai13aa1n12x5               g200(.a(new_n295), .b(new_n289), .c(new_n246), .d(new_n247), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n296), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(new_n291), .b(new_n297), .o1(new_n298));
  xorc02aa1n12x5               g203(.a(\a[25] ), .b(\b[24] ), .out0(new_n299));
  nanb02aa1n06x5               g204(.a(new_n289), .b(new_n248), .out0(new_n300));
  inv000aa1d42x5               g205(.a(new_n299), .o1(new_n301));
  nano23aa1n02x4               g206(.a(new_n294), .b(new_n293), .c(new_n300), .d(new_n301), .out0(new_n302));
  aoi022aa1n02x5               g207(.a(new_n298), .b(new_n299), .c(new_n291), .d(new_n302), .o1(\s[25] ));
  aoai13aa1n03x5               g208(.a(new_n299), .b(new_n296), .c(new_n206), .d(new_n290), .o1(new_n304));
  tech160nm_fixorc02aa1n02p5x5 g209(.a(\a[26] ), .b(\b[25] ), .out0(new_n305));
  nor042aa1n03x5               g210(.a(\b[24] ), .b(\a[25] ), .o1(new_n306));
  norp02aa1n02x5               g211(.a(new_n305), .b(new_n306), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n306), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n301), .c(new_n291), .d(new_n297), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n304), .d(new_n307), .o1(\s[26] ));
  nand22aa1n06x5               g215(.a(new_n305), .b(new_n299), .o1(new_n311));
  nano23aa1n06x5               g216(.a(new_n311), .b(new_n289), .c(new_n220), .d(new_n240), .out0(new_n312));
  aoai13aa1n12x5               g217(.a(new_n312), .b(new_n215), .c(new_n129), .d(new_n196), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n311), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[26] ), .b(\b[25] ), .c(new_n308), .carry(new_n315));
  aobi12aa1n12x5               g220(.a(new_n315), .b(new_n296), .c(new_n314), .out0(new_n316));
  nanp02aa1n03x5               g221(.a(new_n313), .b(new_n316), .o1(new_n317));
  xorc02aa1n12x5               g222(.a(\a[27] ), .b(\b[26] ), .out0(new_n318));
  inv000aa1n02x5               g223(.a(new_n318), .o1(new_n319));
  oai112aa1n02x5               g224(.a(new_n315), .b(new_n319), .c(new_n297), .d(new_n311), .o1(new_n320));
  aboi22aa1n03x5               g225(.a(new_n320), .b(new_n313), .c(new_n317), .d(new_n318), .out0(\s[27] ));
  aoai13aa1n04x5               g226(.a(new_n315), .b(new_n311), .c(new_n300), .d(new_n295), .o1(new_n322));
  aoai13aa1n02x5               g227(.a(new_n318), .b(new_n322), .c(new_n206), .d(new_n312), .o1(new_n323));
  tech160nm_fixorc02aa1n03p5x5 g228(.a(\a[28] ), .b(\b[27] ), .out0(new_n324));
  norp02aa1n02x5               g229(.a(\b[26] ), .b(\a[27] ), .o1(new_n325));
  norp02aa1n02x5               g230(.a(new_n324), .b(new_n325), .o1(new_n326));
  inv000aa1n03x5               g231(.a(new_n325), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n319), .c(new_n313), .d(new_n316), .o1(new_n328));
  aoi022aa1n03x5               g233(.a(new_n328), .b(new_n324), .c(new_n323), .d(new_n326), .o1(\s[28] ));
  and002aa1n02x5               g234(.a(new_n324), .b(new_n318), .o(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n322), .c(new_n206), .d(new_n312), .o1(new_n331));
  inv000aa1d42x5               g236(.a(new_n330), .o1(new_n332));
  oao003aa1n02x5               g237(.a(\a[28] ), .b(\b[27] ), .c(new_n327), .carry(new_n333));
  aoai13aa1n03x5               g238(.a(new_n333), .b(new_n332), .c(new_n313), .d(new_n316), .o1(new_n334));
  tech160nm_fixorc02aa1n03p5x5 g239(.a(\a[29] ), .b(\b[28] ), .out0(new_n335));
  norb02aa1n02x5               g240(.a(new_n333), .b(new_n335), .out0(new_n336));
  aoi022aa1n03x5               g241(.a(new_n334), .b(new_n335), .c(new_n331), .d(new_n336), .o1(\s[29] ));
  xorb03aa1n02x5               g242(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g243(.a(new_n319), .b(new_n324), .c(new_n335), .out0(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n322), .c(new_n206), .d(new_n312), .o1(new_n340));
  inv000aa1d42x5               g245(.a(new_n339), .o1(new_n341));
  oao003aa1n02x5               g246(.a(\a[29] ), .b(\b[28] ), .c(new_n333), .carry(new_n342));
  aoai13aa1n03x5               g247(.a(new_n342), .b(new_n341), .c(new_n313), .d(new_n316), .o1(new_n343));
  tech160nm_fixorc02aa1n03p5x5 g248(.a(\a[30] ), .b(\b[29] ), .out0(new_n344));
  norb02aa1n02x5               g249(.a(new_n342), .b(new_n344), .out0(new_n345));
  aoi022aa1n03x5               g250(.a(new_n343), .b(new_n344), .c(new_n340), .d(new_n345), .o1(\s[30] ));
  nano32aa1n02x5               g251(.a(new_n319), .b(new_n344), .c(new_n324), .d(new_n335), .out0(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n322), .c(new_n206), .d(new_n312), .o1(new_n348));
  xorc02aa1n02x5               g253(.a(\a[31] ), .b(\b[30] ), .out0(new_n349));
  oao003aa1n02x5               g254(.a(\a[30] ), .b(\b[29] ), .c(new_n342), .carry(new_n350));
  norb02aa1n02x5               g255(.a(new_n350), .b(new_n349), .out0(new_n351));
  inv000aa1d42x5               g256(.a(new_n347), .o1(new_n352));
  aoai13aa1n03x5               g257(.a(new_n350), .b(new_n352), .c(new_n313), .d(new_n316), .o1(new_n353));
  aoi022aa1n03x5               g258(.a(new_n353), .b(new_n349), .c(new_n348), .d(new_n351), .o1(\s[31] ));
  aoi112aa1n02x5               g259(.a(new_n109), .b(new_n99), .c(new_n101), .d(new_n102), .o1(new_n355));
  aoi012aa1n02x5               g260(.a(new_n355), .b(new_n103), .c(new_n109), .o1(\s[3] ));
  oaoi03aa1n02x5               g261(.a(\a[3] ), .b(\b[2] ), .c(new_n154), .o1(new_n357));
  aoi112aa1n02x5               g262(.a(new_n107), .b(new_n106), .c(new_n103), .d(new_n108), .o1(new_n358));
  aoi012aa1n02x5               g263(.a(new_n358), .b(new_n106), .c(new_n357), .o1(\s[4] ));
  norb02aa1n02x5               g264(.a(new_n115), .b(new_n114), .out0(new_n360));
  xnbna2aa1n03x5               g265(.a(new_n360), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  norb02aa1n02x5               g266(.a(new_n113), .b(new_n112), .out0(new_n362));
  aoai13aa1n02x5               g267(.a(new_n362), .b(new_n114), .c(new_n156), .d(new_n115), .o1(new_n363));
  aoi112aa1n02x5               g268(.a(new_n114), .b(new_n362), .c(new_n156), .d(new_n360), .o1(new_n364));
  norb02aa1n02x5               g269(.a(new_n363), .b(new_n364), .out0(\s[6] ));
  inv000aa1d42x5               g270(.a(new_n112), .o1(new_n366));
  norb02aa1n02x5               g271(.a(new_n120), .b(new_n119), .out0(new_n367));
  xnbna2aa1n03x5               g272(.a(new_n367), .b(new_n363), .c(new_n366), .out0(\s[7] ));
  aob012aa1n02x5               g273(.a(new_n367), .b(new_n363), .c(new_n366), .out0(new_n369));
  nanp02aa1n02x5               g274(.a(new_n369), .b(new_n126), .o1(new_n370));
  aoib12aa1n02x5               g275(.a(new_n119), .b(new_n118), .c(new_n117), .out0(new_n371));
  aoi022aa1n02x5               g276(.a(new_n370), .b(new_n123), .c(new_n369), .d(new_n371), .o1(\s[8] ));
  aoi113aa1n02x5               g277(.a(new_n130), .b(new_n127), .c(new_n124), .d(new_n125), .e(new_n123), .o1(new_n373));
  aoi022aa1n02x5               g278(.a(new_n129), .b(new_n130), .c(new_n157), .d(new_n373), .o1(\s[9] ));
endmodule


