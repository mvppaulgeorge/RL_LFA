// Benchmark "adder" written by ABC on Wed Jul 17 16:58:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n358,
    new_n359, new_n360, new_n361, new_n363, new_n364, new_n366, new_n368,
    new_n369, new_n370, new_n372, new_n373, new_n375, new_n376, new_n378,
    new_n379;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1n20x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand22aa1n12x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oaoi03aa1n12x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nand02aa1d28x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand02aa1d16x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1d18x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  aoi012aa1n12x5               g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1d24x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  nanp02aa1n24x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand02aa1n06x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n113), .b(new_n116), .c(new_n115), .d(new_n114), .out0(new_n117));
  xnrc02aa1n12x5               g022(.a(\b[7] ), .b(\a[8] ), .out0(new_n118));
  xnrc02aa1n12x5               g023(.a(\b[6] ), .b(\a[7] ), .out0(new_n119));
  nor043aa1n09x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\a[8] ), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\b[7] ), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  inv040aa1d32x5               g028(.a(\a[7] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[6] ), .o1(new_n125));
  nand42aa1n02x5               g030(.a(new_n125), .b(new_n124), .o1(new_n126));
  tech160nm_fioai012aa1n03p5x5 g031(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n127));
  aoi022aa1d24x5               g032(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n128));
  inv030aa1n02x5               g033(.a(new_n128), .o1(new_n129));
  aoai13aa1n09x5               g034(.a(new_n123), .b(new_n129), .c(new_n127), .d(new_n126), .o1(new_n130));
  nanp02aa1n09x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n100), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n130), .c(new_n112), .d(new_n120), .o1(new_n133));
  xobna2aa1n03x5               g038(.a(new_n99), .b(new_n133), .c(new_n101), .out0(\s[10] ));
  nand42aa1n20x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor002aa1d32x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  inv040aa1n03x5               g042(.a(new_n104), .o1(new_n138));
  oaoi03aa1n12x5               g043(.a(\a[2] ), .b(\b[1] ), .c(new_n138), .o1(new_n139));
  nano23aa1n09x5               g044(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n140));
  nanp02aa1n06x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  nano23aa1n02x4               g046(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n142));
  nona22aa1n03x5               g047(.a(new_n142), .b(new_n118), .c(new_n119), .out0(new_n143));
  nand02aa1n02x5               g048(.a(new_n127), .b(new_n126), .o1(new_n144));
  aoi022aa1n03x5               g049(.a(new_n144), .b(new_n128), .c(new_n122), .d(new_n121), .o1(new_n145));
  aoai13aa1n04x5               g050(.a(new_n145), .b(new_n143), .c(new_n141), .d(new_n111), .o1(new_n146));
  oaih22aa1d12x5               g051(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n147));
  aoai13aa1n02x5               g052(.a(new_n98), .b(new_n147), .c(new_n146), .d(new_n132), .o1(new_n148));
  nano22aa1n02x4               g053(.a(new_n136), .b(new_n98), .c(new_n135), .out0(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n147), .c(new_n146), .d(new_n132), .o1(new_n150));
  aobi12aa1n02x5               g055(.a(new_n150), .b(new_n148), .c(new_n137), .out0(\s[11] ));
  inv000aa1d42x5               g056(.a(new_n136), .o1(new_n152));
  nor002aa1d32x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  nand42aa1d28x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  norb03aa1n12x5               g060(.a(new_n154), .b(new_n136), .c(new_n153), .out0(new_n156));
  nanp02aa1n02x5               g061(.a(new_n150), .b(new_n156), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n155), .c(new_n150), .d(new_n152), .o1(\s[12] ));
  nano23aa1n09x5               g063(.a(new_n153), .b(new_n136), .c(new_n154), .d(new_n135), .out0(new_n159));
  nano23aa1n09x5               g064(.a(new_n97), .b(new_n100), .c(new_n131), .d(new_n98), .out0(new_n160));
  nanp02aa1n03x5               g065(.a(new_n160), .b(new_n159), .o1(new_n161));
  inv000aa1n02x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n130), .c(new_n112), .d(new_n120), .o1(new_n163));
  aoi022aa1n06x5               g068(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n164));
  aoi012aa1d18x5               g069(.a(new_n153), .b(new_n136), .c(new_n154), .o1(new_n165));
  inv000aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  aoi013aa1n03x5               g071(.a(new_n166), .b(new_n156), .c(new_n164), .d(new_n147), .o1(new_n167));
  tech160nm_finand02aa1n05x5   g072(.a(new_n163), .b(new_n167), .o1(new_n168));
  nor002aa1d32x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nand42aa1d28x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  aoi113aa1n02x5               g076(.a(new_n171), .b(new_n166), .c(new_n156), .d(new_n164), .e(new_n147), .o1(new_n172));
  aoi022aa1n02x5               g077(.a(new_n168), .b(new_n171), .c(new_n163), .d(new_n172), .o1(\s[13] ));
  aoi012aa1n02x5               g078(.a(new_n169), .b(new_n168), .c(new_n170), .o1(new_n174));
  nor002aa1d32x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nand42aa1d28x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  nand23aa1n06x5               g082(.a(new_n156), .b(new_n147), .c(new_n164), .o1(new_n178));
  nand22aa1n03x5               g083(.a(new_n178), .b(new_n165), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n171), .b(new_n179), .c(new_n146), .d(new_n162), .o1(new_n180));
  nona23aa1n02x4               g085(.a(new_n180), .b(new_n176), .c(new_n175), .d(new_n169), .out0(new_n181));
  oai012aa1n02x5               g086(.a(new_n181), .b(new_n174), .c(new_n177), .o1(\s[14] ));
  nano23aa1d15x5               g087(.a(new_n169), .b(new_n175), .c(new_n176), .d(new_n170), .out0(new_n183));
  oai012aa1d24x5               g088(.a(new_n176), .b(new_n175), .c(new_n169), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n184), .o1(new_n185));
  xorc02aa1n12x5               g090(.a(\a[15] ), .b(\b[14] ), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n185), .c(new_n168), .d(new_n183), .o1(new_n187));
  aoi112aa1n02x5               g092(.a(new_n186), .b(new_n185), .c(new_n168), .d(new_n183), .o1(new_n188));
  norb02aa1n02x5               g093(.a(new_n187), .b(new_n188), .out0(\s[15] ));
  orn002aa1n24x5               g094(.a(\a[15] ), .b(\b[14] ), .o(new_n190));
  nor042aa1d18x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  and002aa1n12x5               g096(.a(\b[15] ), .b(\a[16] ), .o(new_n192));
  nor042aa1n06x5               g097(.a(new_n192), .b(new_n191), .o1(new_n193));
  oai022aa1n02x5               g098(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n194));
  nona22aa1n03x5               g099(.a(new_n187), .b(new_n192), .c(new_n194), .out0(new_n195));
  aoai13aa1n02x5               g100(.a(new_n195), .b(new_n193), .c(new_n190), .d(new_n187), .o1(\s[16] ));
  nand23aa1n06x5               g101(.a(new_n183), .b(new_n186), .c(new_n193), .o1(new_n197));
  nor042aa1n06x5               g102(.a(new_n197), .b(new_n161), .o1(new_n198));
  aoai13aa1n12x5               g103(.a(new_n198), .b(new_n130), .c(new_n112), .d(new_n120), .o1(new_n199));
  nona23aa1n02x5               g104(.a(new_n176), .b(new_n170), .c(new_n169), .d(new_n175), .out0(new_n200));
  nanp02aa1n02x5               g105(.a(\b[14] ), .b(\a[15] ), .o1(new_n201));
  nano32aa1n06x5               g106(.a(new_n200), .b(new_n193), .c(new_n190), .d(new_n201), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n191), .o1(new_n203));
  aob012aa1n02x5               g108(.a(new_n201), .b(\b[15] ), .c(\a[16] ), .out0(new_n204));
  aoai13aa1n09x5               g109(.a(new_n203), .b(new_n204), .c(new_n184), .d(new_n190), .o1(new_n205));
  aoi012aa1n12x5               g110(.a(new_n205), .b(new_n179), .c(new_n202), .o1(new_n206));
  nanp02aa1n12x5               g111(.a(new_n199), .b(new_n206), .o1(new_n207));
  nor002aa1d32x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  nand42aa1n16x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi012aa1n02x5               g115(.a(new_n204), .b(new_n184), .c(new_n190), .o1(new_n211));
  oaib12aa1n02x5               g116(.a(new_n203), .b(new_n208), .c(new_n209), .out0(new_n212));
  aoi112aa1n02x5               g117(.a(new_n212), .b(new_n211), .c(new_n179), .d(new_n202), .o1(new_n213));
  aoi022aa1n02x5               g118(.a(new_n207), .b(new_n210), .c(new_n199), .d(new_n213), .o1(\s[17] ));
  inv000aa1d42x5               g119(.a(new_n208), .o1(new_n215));
  oabi12aa1n03x5               g120(.a(new_n205), .b(new_n167), .c(new_n197), .out0(new_n216));
  aoai13aa1n03x5               g121(.a(new_n210), .b(new_n216), .c(new_n146), .d(new_n198), .o1(new_n217));
  nor042aa1d18x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  nand42aa1d28x5               g123(.a(\b[17] ), .b(\a[18] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  nona23aa1n02x4               g125(.a(new_n217), .b(new_n219), .c(new_n218), .d(new_n208), .out0(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n220), .c(new_n215), .d(new_n217), .o1(\s[18] ));
  nano23aa1d15x5               g127(.a(new_n208), .b(new_n218), .c(new_n219), .d(new_n209), .out0(new_n223));
  oaoi03aa1n02x5               g128(.a(\a[18] ), .b(\b[17] ), .c(new_n215), .o1(new_n224));
  nor042aa1d18x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  nand22aa1n06x5               g130(.a(\b[18] ), .b(\a[19] ), .o1(new_n226));
  norb02aa1n09x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n207), .d(new_n223), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n227), .b(new_n224), .c(new_n207), .d(new_n223), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n228), .b(new_n229), .out0(\s[19] ));
  xnrc02aa1n02x5               g135(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n02x5               g136(.a(new_n225), .o1(new_n232));
  nor002aa1n20x5               g137(.a(\b[19] ), .b(\a[20] ), .o1(new_n233));
  nand22aa1n12x5               g138(.a(\b[19] ), .b(\a[20] ), .o1(new_n234));
  norb02aa1n12x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  norb03aa1n02x5               g140(.a(new_n234), .b(new_n225), .c(new_n233), .out0(new_n236));
  tech160nm_finand02aa1n03p5x5 g141(.a(new_n228), .b(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n235), .c(new_n232), .d(new_n228), .o1(\s[20] ));
  nand23aa1n09x5               g143(.a(new_n223), .b(new_n227), .c(new_n235), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nanb03aa1n06x5               g145(.a(new_n233), .b(new_n234), .c(new_n226), .out0(new_n241));
  oai112aa1n06x5               g146(.a(new_n232), .b(new_n219), .c(new_n218), .d(new_n208), .o1(new_n242));
  aoi012aa1d24x5               g147(.a(new_n233), .b(new_n225), .c(new_n234), .o1(new_n243));
  oai012aa1n06x5               g148(.a(new_n243), .b(new_n242), .c(new_n241), .o1(new_n244));
  nor042aa1n12x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  nand42aa1n02x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  norb02aa1n02x5               g151(.a(new_n246), .b(new_n245), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n244), .c(new_n207), .d(new_n240), .o1(new_n248));
  nano22aa1n03x7               g153(.a(new_n233), .b(new_n226), .c(new_n234), .out0(new_n249));
  tech160nm_fioai012aa1n03p5x5 g154(.a(new_n219), .b(\b[18] ), .c(\a[19] ), .o1(new_n250));
  oab012aa1n06x5               g155(.a(new_n250), .b(new_n208), .c(new_n218), .out0(new_n251));
  inv000aa1n02x5               g156(.a(new_n243), .o1(new_n252));
  aoi112aa1n02x5               g157(.a(new_n252), .b(new_n247), .c(new_n251), .d(new_n249), .o1(new_n253));
  aobi12aa1n02x5               g158(.a(new_n253), .b(new_n207), .c(new_n240), .out0(new_n254));
  norb02aa1n03x4               g159(.a(new_n248), .b(new_n254), .out0(\s[21] ));
  inv000aa1d42x5               g160(.a(new_n245), .o1(new_n256));
  nor042aa1n03x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  nand02aa1d08x5               g162(.a(\b[21] ), .b(\a[22] ), .o1(new_n258));
  norb02aa1n02x5               g163(.a(new_n258), .b(new_n257), .out0(new_n259));
  norb03aa1n02x5               g164(.a(new_n258), .b(new_n245), .c(new_n257), .out0(new_n260));
  tech160nm_finand02aa1n03p5x5 g165(.a(new_n248), .b(new_n260), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n259), .c(new_n256), .d(new_n248), .o1(\s[22] ));
  nano23aa1n06x5               g167(.a(new_n245), .b(new_n257), .c(new_n258), .d(new_n246), .out0(new_n263));
  norb02aa1n02x5               g168(.a(new_n263), .b(new_n239), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n263), .b(new_n252), .c(new_n251), .d(new_n249), .o1(new_n265));
  aoi012aa1n12x5               g170(.a(new_n257), .b(new_n245), .c(new_n258), .o1(new_n266));
  nanp02aa1n02x5               g171(.a(new_n265), .b(new_n266), .o1(new_n267));
  nor042aa1d18x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  nanp02aa1n04x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  norb02aa1n02x5               g174(.a(new_n269), .b(new_n268), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n267), .c(new_n207), .d(new_n264), .o1(new_n271));
  inv000aa1n02x5               g176(.a(new_n266), .o1(new_n272));
  nona22aa1n02x4               g177(.a(new_n265), .b(new_n272), .c(new_n270), .out0(new_n273));
  aoi012aa1n02x5               g178(.a(new_n273), .b(new_n207), .c(new_n264), .o1(new_n274));
  norb02aa1n03x4               g179(.a(new_n271), .b(new_n274), .out0(\s[23] ));
  inv040aa1d28x5               g180(.a(new_n268), .o1(new_n276));
  nor042aa1n04x5               g181(.a(\b[23] ), .b(\a[24] ), .o1(new_n277));
  and002aa1n12x5               g182(.a(\b[23] ), .b(\a[24] ), .o(new_n278));
  norp02aa1n02x5               g183(.a(new_n278), .b(new_n277), .o1(new_n279));
  norp03aa1n02x5               g184(.a(new_n278), .b(new_n277), .c(new_n268), .o1(new_n280));
  tech160nm_finand02aa1n03p5x5 g185(.a(new_n271), .b(new_n280), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n279), .c(new_n276), .d(new_n271), .o1(\s[24] ));
  nano32aa1n02x5               g187(.a(new_n239), .b(new_n279), .c(new_n263), .d(new_n270), .out0(new_n283));
  nano23aa1d15x5               g188(.a(new_n278), .b(new_n277), .c(new_n276), .d(new_n269), .out0(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  oab012aa1n04x5               g190(.a(new_n277), .b(new_n276), .c(new_n278), .out0(new_n286));
  aoai13aa1n04x5               g191(.a(new_n286), .b(new_n285), .c(new_n265), .d(new_n266), .o1(new_n287));
  xorc02aa1n12x5               g192(.a(\a[25] ), .b(\b[24] ), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n287), .c(new_n207), .d(new_n283), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n284), .b(new_n272), .c(new_n244), .d(new_n263), .o1(new_n290));
  nanb03aa1n02x5               g195(.a(new_n288), .b(new_n290), .c(new_n286), .out0(new_n291));
  aoi012aa1n02x5               g196(.a(new_n291), .b(new_n207), .c(new_n283), .o1(new_n292));
  norb02aa1n03x4               g197(.a(new_n289), .b(new_n292), .out0(\s[25] ));
  nor042aa1n04x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  nor042aa1n04x5               g200(.a(\b[25] ), .b(\a[26] ), .o1(new_n296));
  and002aa1n12x5               g201(.a(\b[25] ), .b(\a[26] ), .o(new_n297));
  nor042aa1n04x5               g202(.a(new_n297), .b(new_n296), .o1(new_n298));
  norp03aa1n02x5               g203(.a(new_n297), .b(new_n296), .c(new_n294), .o1(new_n299));
  tech160nm_finand02aa1n03p5x5 g204(.a(new_n289), .b(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n298), .c(new_n295), .d(new_n289), .o1(\s[26] ));
  nand42aa1n06x5               g206(.a(new_n288), .b(new_n298), .o1(new_n302));
  nano23aa1n06x5               g207(.a(new_n239), .b(new_n302), .c(new_n284), .d(new_n263), .out0(new_n303));
  aoai13aa1n06x5               g208(.a(new_n303), .b(new_n216), .c(new_n146), .d(new_n198), .o1(new_n304));
  aobi12aa1n06x5               g209(.a(new_n303), .b(new_n199), .c(new_n206), .out0(new_n305));
  oab012aa1n09x5               g210(.a(new_n296), .b(new_n295), .c(new_n297), .out0(new_n306));
  aoai13aa1n04x5               g211(.a(new_n306), .b(new_n302), .c(new_n290), .d(new_n286), .o1(new_n307));
  xorc02aa1n12x5               g212(.a(\a[27] ), .b(\b[26] ), .out0(new_n308));
  oai012aa1n06x5               g213(.a(new_n308), .b(new_n307), .c(new_n305), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n302), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n306), .o1(new_n311));
  aoi112aa1n02x5               g216(.a(new_n308), .b(new_n311), .c(new_n287), .d(new_n310), .o1(new_n312));
  aobi12aa1n02x7               g217(.a(new_n309), .b(new_n312), .c(new_n304), .out0(\s[27] ));
  nor042aa1d18x5               g218(.a(\b[26] ), .b(\a[27] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .out0(new_n316));
  tech160nm_fiaoi012aa1n05x5   g221(.a(new_n311), .b(new_n287), .c(new_n310), .o1(new_n317));
  inv000aa1n03x5               g222(.a(new_n308), .o1(new_n318));
  inv000aa1d42x5               g223(.a(\a[28] ), .o1(new_n319));
  inv000aa1d42x5               g224(.a(\b[27] ), .o1(new_n320));
  aoi012aa1d24x5               g225(.a(new_n314), .b(new_n319), .c(new_n320), .o1(new_n321));
  oa0012aa1n02x5               g226(.a(new_n321), .b(new_n320), .c(new_n319), .o(new_n322));
  aoai13aa1n02x7               g227(.a(new_n322), .b(new_n318), .c(new_n317), .d(new_n304), .o1(new_n323));
  aoai13aa1n03x5               g228(.a(new_n323), .b(new_n316), .c(new_n309), .d(new_n315), .o1(\s[28] ));
  and002aa1n02x5               g229(.a(new_n316), .b(new_n308), .o(new_n325));
  oaih12aa1n02x5               g230(.a(new_n325), .b(new_n307), .c(new_n305), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n325), .o1(new_n327));
  oaoi03aa1n02x5               g232(.a(new_n319), .b(new_n320), .c(new_n314), .o1(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n327), .c(new_n317), .d(new_n304), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[29] ), .b(\b[28] ), .out0(new_n330));
  inv000aa1d42x5               g235(.a(new_n321), .o1(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n330), .b(new_n331), .c(new_n319), .d(new_n320), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n329), .b(new_n330), .c(new_n326), .d(new_n332), .o1(\s[29] ));
  xorb03aa1n02x5               g238(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g239(.a(new_n318), .b(new_n316), .c(new_n330), .out0(new_n335));
  oaih12aa1n02x5               g240(.a(new_n335), .b(new_n307), .c(new_n305), .o1(new_n336));
  inv000aa1n02x5               g241(.a(new_n335), .o1(new_n337));
  aoi022aa1n03x5               g242(.a(\b[28] ), .b(\a[29] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n338));
  obai22aa1n06x5               g243(.a(new_n338), .b(new_n321), .c(\a[29] ), .d(\b[28] ), .out0(new_n339));
  inv000aa1d42x5               g244(.a(new_n339), .o1(new_n340));
  aoai13aa1n03x5               g245(.a(new_n340), .b(new_n337), .c(new_n317), .d(new_n304), .o1(new_n341));
  xorc02aa1n02x5               g246(.a(\a[30] ), .b(\b[29] ), .out0(new_n342));
  norp02aa1n02x5               g247(.a(\b[28] ), .b(\a[29] ), .o1(new_n343));
  aoi112aa1n02x5               g248(.a(new_n343), .b(new_n342), .c(new_n331), .d(new_n338), .o1(new_n344));
  aoi022aa1n03x5               g249(.a(new_n341), .b(new_n342), .c(new_n336), .d(new_n344), .o1(\s[30] ));
  nano32aa1n02x4               g250(.a(new_n318), .b(new_n342), .c(new_n316), .d(new_n330), .out0(new_n346));
  oaih12aa1n02x5               g251(.a(new_n346), .b(new_n307), .c(new_n305), .o1(new_n347));
  inv000aa1d42x5               g252(.a(\a[30] ), .o1(new_n348));
  inv000aa1d42x5               g253(.a(\b[29] ), .o1(new_n349));
  aboi22aa1n03x5               g254(.a(\b[30] ), .b(\a[31] ), .c(new_n348), .d(new_n349), .out0(new_n350));
  oaib12aa1n02x5               g255(.a(new_n350), .b(\a[31] ), .c(\b[30] ), .out0(new_n351));
  oaoi13aa1n02x5               g256(.a(new_n351), .b(new_n339), .c(new_n348), .d(new_n349), .o1(new_n352));
  xorc02aa1n02x5               g257(.a(\a[31] ), .b(\b[30] ), .out0(new_n353));
  inv000aa1n02x5               g258(.a(new_n346), .o1(new_n354));
  oaoi03aa1n02x5               g259(.a(new_n348), .b(new_n349), .c(new_n339), .o1(new_n355));
  aoai13aa1n03x5               g260(.a(new_n355), .b(new_n354), .c(new_n317), .d(new_n304), .o1(new_n356));
  aoi022aa1n03x5               g261(.a(new_n356), .b(new_n353), .c(new_n347), .d(new_n352), .o1(\s[31] ));
  aoi022aa1n02x5               g262(.a(new_n103), .b(new_n102), .c(\a[1] ), .d(\b[0] ), .o1(new_n358));
  oaib12aa1n02x5               g263(.a(new_n358), .b(new_n103), .c(\a[2] ), .out0(new_n359));
  norb02aa1n02x5               g264(.a(new_n109), .b(new_n108), .out0(new_n360));
  aboi22aa1n03x5               g265(.a(new_n108), .b(new_n109), .c(new_n102), .d(new_n103), .out0(new_n361));
  aoi022aa1n02x5               g266(.a(new_n359), .b(new_n361), .c(new_n139), .d(new_n360), .o1(\s[3] ));
  obai22aa1n02x7               g267(.a(new_n107), .b(new_n106), .c(\a[3] ), .d(\b[2] ), .out0(new_n363));
  aoi012aa1n02x5               g268(.a(new_n363), .b(new_n139), .c(new_n360), .o1(new_n364));
  oaoi13aa1n02x5               g269(.a(new_n364), .b(new_n112), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  norb02aa1n02x5               g270(.a(new_n116), .b(new_n115), .out0(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n366), .b(new_n141), .c(new_n111), .out0(\s[5] ));
  norb02aa1n02x5               g272(.a(new_n113), .b(new_n114), .out0(new_n368));
  aoai13aa1n02x5               g273(.a(new_n368), .b(new_n115), .c(new_n112), .d(new_n116), .o1(new_n369));
  aoi112aa1n02x5               g274(.a(new_n115), .b(new_n368), .c(new_n112), .d(new_n366), .o1(new_n370));
  norb02aa1n02x5               g275(.a(new_n369), .b(new_n370), .out0(\s[6] ));
  nanb02aa1n02x5               g276(.a(new_n114), .b(new_n369), .out0(new_n372));
  nona22aa1n02x4               g277(.a(new_n369), .b(new_n119), .c(new_n114), .out0(new_n373));
  aob012aa1n02x5               g278(.a(new_n373), .b(new_n372), .c(new_n119), .out0(\s[7] ));
  and002aa1n02x5               g279(.a(\b[6] ), .b(\a[7] ), .o(new_n375));
  inv000aa1d42x5               g280(.a(new_n375), .o1(new_n376));
  xnbna2aa1n03x5               g281(.a(new_n118), .b(new_n373), .c(new_n376), .out0(\s[8] ));
  nanp02aa1n02x5               g282(.a(new_n112), .b(new_n120), .o1(new_n378));
  aoi122aa1n02x5               g283(.a(new_n132), .b(new_n122), .c(new_n121), .d(new_n144), .e(new_n128), .o1(new_n379));
  aoi022aa1n02x5               g284(.a(new_n146), .b(new_n132), .c(new_n378), .d(new_n379), .o1(\s[9] ));
endmodule


