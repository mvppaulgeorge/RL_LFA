// Benchmark "adder" written by ABC on Thu Jul 18 09:15:24 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n216, new_n217, new_n218, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n301, new_n304, new_n305,
    new_n307, new_n309;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  nor002aa1n08x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  xnrc02aa1n12x5               g003(.a(\b[7] ), .b(\a[8] ), .out0(new_n99));
  xnrc02aa1n06x5               g004(.a(\b[6] ), .b(\a[7] ), .out0(new_n100));
  nor042aa1n02x5               g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  nor022aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor022aa1n08x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n03x5               g010(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n106));
  nanp02aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nor002aa1n02x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nand22aa1n03x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  tech160nm_fioai012aa1n05x5   g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  oai012aa1n02x5               g015(.a(new_n103), .b(new_n104), .c(new_n102), .o1(new_n111));
  oai012aa1n04x7               g016(.a(new_n111), .b(new_n106), .c(new_n110), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[5] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\a[6] ), .o1(new_n114));
  xroi22aa1d04x5               g019(.a(new_n113), .b(\b[4] ), .c(new_n114), .d(\b[5] ), .out0(new_n115));
  nand23aa1n06x5               g020(.a(new_n112), .b(new_n101), .c(new_n115), .o1(new_n116));
  aoi112aa1n03x5               g021(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n117));
  aoib12aa1n02x5               g022(.a(new_n117), .b(new_n114), .c(\b[5] ), .out0(new_n118));
  orn002aa1n02x5               g023(.a(\a[7] ), .b(\b[6] ), .o(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  aoib12aa1n12x5               g025(.a(new_n120), .b(new_n101), .c(new_n118), .out0(new_n121));
  nanp02aa1n02x5               g026(.a(new_n116), .b(new_n121), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  nanp02aa1n02x5               g028(.a(new_n122), .b(new_n123), .o1(new_n124));
  nona22aa1n02x4               g029(.a(new_n124), .b(new_n98), .c(new_n97), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n97), .b(new_n98), .c(new_n122), .d(new_n123), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(new_n125), .b(new_n126), .o1(\s[10] ));
  aoi112aa1n02x5               g032(.a(new_n97), .b(new_n98), .c(new_n122), .d(new_n123), .o1(new_n128));
  xnrc02aa1n12x5               g033(.a(\b[10] ), .b(\a[11] ), .out0(new_n129));
  aoi112aa1n02x5               g034(.a(new_n128), .b(new_n129), .c(\a[10] ), .d(\b[9] ), .o1(new_n130));
  inv000aa1d42x5               g035(.a(\a[10] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(\b[9] ), .o1(new_n132));
  xorc02aa1n12x5               g037(.a(\a[11] ), .b(\b[10] ), .out0(new_n133));
  oaoi13aa1n02x5               g038(.a(new_n133), .b(new_n125), .c(new_n131), .d(new_n132), .o1(new_n134));
  norp02aa1n02x5               g039(.a(new_n134), .b(new_n130), .o1(\s[11] ));
  nor002aa1n12x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n136), .o1(new_n137));
  nor002aa1n12x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand22aa1n09x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanb02aa1d24x5               g044(.a(new_n138), .b(new_n139), .out0(new_n140));
  nano22aa1n02x4               g045(.a(new_n130), .b(new_n137), .c(new_n140), .out0(new_n141));
  oai112aa1n02x5               g046(.a(new_n125), .b(new_n133), .c(new_n132), .d(new_n131), .o1(new_n142));
  aoi012aa1n02x5               g047(.a(new_n140), .b(new_n142), .c(new_n137), .o1(new_n143));
  norp02aa1n02x5               g048(.a(new_n143), .b(new_n141), .o1(\s[12] ));
  nano23aa1d15x5               g049(.a(new_n140), .b(new_n97), .c(new_n123), .d(new_n133), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  oaoi03aa1n12x5               g051(.a(new_n131), .b(new_n132), .c(new_n98), .o1(new_n147));
  tech160nm_fiaoi012aa1n04x5   g052(.a(new_n138), .b(new_n136), .c(new_n139), .o1(new_n148));
  oai013aa1n09x5               g053(.a(new_n148), .b(new_n147), .c(new_n129), .d(new_n140), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n146), .c(new_n116), .d(new_n121), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g057(.a(\a[14] ), .o1(new_n153));
  nor022aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  xorc02aa1n02x5               g059(.a(\a[13] ), .b(\b[12] ), .out0(new_n155));
  aoi012aa1n02x5               g060(.a(new_n154), .b(new_n151), .c(new_n155), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(new_n153), .out0(\s[14] ));
  tech160nm_fixorc02aa1n04x5   g062(.a(\a[15] ), .b(\b[14] ), .out0(new_n158));
  xorc02aa1n02x5               g063(.a(\a[14] ), .b(\b[13] ), .out0(new_n159));
  and002aa1n02x5               g064(.a(new_n159), .b(new_n155), .o(new_n160));
  inv000aa1d42x5               g065(.a(\b[13] ), .o1(new_n161));
  oaoi03aa1n12x5               g066(.a(new_n153), .b(new_n161), .c(new_n154), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoai13aa1n03x5               g068(.a(new_n158), .b(new_n163), .c(new_n151), .d(new_n160), .o1(new_n164));
  aoi112aa1n02x5               g069(.a(new_n158), .b(new_n163), .c(new_n151), .d(new_n160), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(\s[15] ));
  xorc02aa1n12x5               g071(.a(\a[16] ), .b(\b[15] ), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  oai112aa1n02x5               g073(.a(new_n164), .b(new_n168), .c(\b[14] ), .d(\a[15] ), .o1(new_n169));
  oaoi13aa1n06x5               g074(.a(new_n168), .b(new_n164), .c(\a[15] ), .d(\b[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nand42aa1n08x5               g076(.a(new_n167), .b(new_n158), .o1(new_n172));
  nano22aa1n03x7               g077(.a(new_n172), .b(new_n155), .c(new_n159), .out0(new_n173));
  nand02aa1d04x5               g078(.a(new_n145), .b(new_n173), .o1(new_n174));
  oai022aa1n02x5               g079(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n175));
  aob012aa1n02x5               g080(.a(new_n175), .b(\b[15] ), .c(\a[16] ), .out0(new_n176));
  oai012aa1n03x5               g081(.a(new_n176), .b(new_n172), .c(new_n162), .o1(new_n177));
  aoi012aa1n06x5               g082(.a(new_n177), .b(new_n149), .c(new_n173), .o1(new_n178));
  aoai13aa1n12x5               g083(.a(new_n178), .b(new_n174), .c(new_n116), .d(new_n121), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g085(.a(\a[18] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  tech160nm_fioaoi03aa1n03p5x5 g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  xroi22aa1d04x5               g090(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n186));
  nanp02aa1n02x5               g091(.a(\b[17] ), .b(\a[18] ), .o1(new_n187));
  nona22aa1n02x4               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(new_n188));
  oaib12aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n181), .out0(new_n189));
  nor002aa1n02x5               g094(.a(\b[18] ), .b(\a[19] ), .o1(new_n190));
  nand42aa1n10x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  norb02aa1n02x5               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n189), .c(new_n179), .d(new_n186), .o1(new_n193));
  aoi112aa1n02x5               g098(.a(new_n192), .b(new_n189), .c(new_n179), .d(new_n186), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g101(.a(\b[19] ), .b(\a[20] ), .o1(new_n197));
  nand42aa1n06x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  nona22aa1n03x5               g104(.a(new_n193), .b(new_n199), .c(new_n190), .out0(new_n200));
  orn002aa1n24x5               g105(.a(\a[19] ), .b(\b[18] ), .o(new_n201));
  aobi12aa1n02x7               g106(.a(new_n199), .b(new_n193), .c(new_n201), .out0(new_n202));
  norb02aa1n03x4               g107(.a(new_n200), .b(new_n202), .out0(\s[20] ));
  nona23aa1n02x4               g108(.a(new_n198), .b(new_n191), .c(new_n190), .d(new_n197), .out0(new_n204));
  norb02aa1n02x5               g109(.a(new_n186), .b(new_n204), .out0(new_n205));
  norp02aa1n02x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  aoi013aa1n02x4               g111(.a(new_n206), .b(new_n187), .c(new_n182), .d(new_n183), .o1(new_n207));
  oaoi03aa1n12x5               g112(.a(\a[20] ), .b(\b[19] ), .c(new_n201), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  tech160nm_fioai012aa1n05x5   g114(.a(new_n209), .b(new_n204), .c(new_n207), .o1(new_n210));
  xnrc02aa1n12x5               g115(.a(\b[20] ), .b(\a[21] ), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n04x5               g117(.a(new_n212), .b(new_n210), .c(new_n179), .d(new_n205), .o1(new_n213));
  aoi112aa1n02x5               g118(.a(new_n212), .b(new_n210), .c(new_n179), .d(new_n205), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(\s[21] ));
  xnrc02aa1n02x5               g120(.a(\b[21] ), .b(\a[22] ), .out0(new_n216));
  oai112aa1n03x5               g121(.a(new_n213), .b(new_n216), .c(\b[20] ), .d(\a[21] ), .o1(new_n217));
  oaoi13aa1n03x5               g122(.a(new_n216), .b(new_n213), .c(\a[21] ), .d(\b[20] ), .o1(new_n218));
  norb02aa1n02x7               g123(.a(new_n217), .b(new_n218), .out0(\s[22] ));
  nano23aa1n03x5               g124(.a(new_n190), .b(new_n197), .c(new_n198), .d(new_n191), .out0(new_n220));
  nor002aa1n03x5               g125(.a(new_n216), .b(new_n211), .o1(new_n221));
  and003aa1n06x5               g126(.a(new_n186), .b(new_n221), .c(new_n220), .o(new_n222));
  aoai13aa1n06x5               g127(.a(new_n221), .b(new_n208), .c(new_n220), .d(new_n189), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\a[22] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\b[21] ), .o1(new_n225));
  norp02aa1n02x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  oao003aa1n02x5               g131(.a(new_n224), .b(new_n225), .c(new_n226), .carry(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(new_n223), .b(new_n228), .o1(new_n229));
  xorc02aa1n12x5               g134(.a(\a[23] ), .b(\b[22] ), .out0(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n229), .c(new_n179), .d(new_n222), .o1(new_n231));
  aoi112aa1n02x5               g136(.a(new_n230), .b(new_n229), .c(new_n179), .d(new_n222), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n231), .b(new_n232), .out0(\s[23] ));
  norp02aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  xorc02aa1n02x5               g139(.a(\a[24] ), .b(\b[23] ), .out0(new_n235));
  nona22aa1n02x4               g140(.a(new_n231), .b(new_n235), .c(new_n234), .out0(new_n236));
  inv000aa1n02x5               g141(.a(new_n234), .o1(new_n237));
  aobi12aa1n03x5               g142(.a(new_n235), .b(new_n231), .c(new_n237), .out0(new_n238));
  norb02aa1n03x4               g143(.a(new_n236), .b(new_n238), .out0(\s[24] ));
  and002aa1n02x5               g144(.a(new_n235), .b(new_n230), .o(new_n240));
  inv000aa1n02x5               g145(.a(new_n240), .o1(new_n241));
  nano32aa1n02x4               g146(.a(new_n241), .b(new_n186), .c(new_n221), .d(new_n220), .out0(new_n242));
  oao003aa1n02x5               g147(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .carry(new_n243));
  aoai13aa1n04x5               g148(.a(new_n243), .b(new_n241), .c(new_n223), .d(new_n228), .o1(new_n244));
  xorc02aa1n02x5               g149(.a(\a[25] ), .b(\b[24] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n244), .c(new_n179), .d(new_n242), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n245), .b(new_n244), .c(new_n179), .d(new_n242), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[26] ), .b(\b[25] ), .out0(new_n250));
  nona22aa1n03x5               g155(.a(new_n246), .b(new_n250), .c(new_n249), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n249), .o1(new_n252));
  aobi12aa1n03x5               g157(.a(new_n250), .b(new_n246), .c(new_n252), .out0(new_n253));
  norb02aa1n03x4               g158(.a(new_n251), .b(new_n253), .out0(\s[26] ));
  inv000aa1d42x5               g159(.a(\a[25] ), .o1(new_n255));
  inv040aa1d32x5               g160(.a(\a[26] ), .o1(new_n256));
  xroi22aa1d06x4               g161(.a(new_n255), .b(\b[24] ), .c(new_n256), .d(\b[25] ), .out0(new_n257));
  and003aa1n12x5               g162(.a(new_n222), .b(new_n257), .c(new_n240), .o(new_n258));
  nand02aa1d08x5               g163(.a(new_n179), .b(new_n258), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .c(new_n252), .carry(new_n260));
  aobi12aa1n06x5               g165(.a(new_n260), .b(new_n244), .c(new_n257), .out0(new_n261));
  xorc02aa1n02x5               g166(.a(\a[27] ), .b(\b[26] ), .out0(new_n262));
  xnbna2aa1n03x5               g167(.a(new_n262), .b(new_n259), .c(new_n261), .out0(\s[27] ));
  norp02aa1n02x5               g168(.a(\b[26] ), .b(\a[27] ), .o1(new_n264));
  inv040aa1n03x5               g169(.a(new_n264), .o1(new_n265));
  aobi12aa1n03x5               g170(.a(new_n262), .b(new_n259), .c(new_n261), .out0(new_n266));
  xnrc02aa1n02x5               g171(.a(\b[27] ), .b(\a[28] ), .out0(new_n267));
  nano22aa1n03x5               g172(.a(new_n266), .b(new_n265), .c(new_n267), .out0(new_n268));
  aoai13aa1n02x5               g173(.a(new_n240), .b(new_n227), .c(new_n210), .d(new_n221), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n257), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n260), .b(new_n270), .c(new_n269), .d(new_n243), .o1(new_n271));
  aoai13aa1n02x7               g176(.a(new_n262), .b(new_n271), .c(new_n179), .d(new_n258), .o1(new_n272));
  tech160nm_fiaoi012aa1n02p5x5 g177(.a(new_n267), .b(new_n272), .c(new_n265), .o1(new_n273));
  norp02aa1n03x5               g178(.a(new_n273), .b(new_n268), .o1(\s[28] ));
  norb02aa1n02x5               g179(.a(new_n262), .b(new_n267), .out0(new_n275));
  aobi12aa1n03x5               g180(.a(new_n275), .b(new_n259), .c(new_n261), .out0(new_n276));
  oao003aa1n02x5               g181(.a(\a[28] ), .b(\b[27] ), .c(new_n265), .carry(new_n277));
  xnrc02aa1n02x5               g182(.a(\b[28] ), .b(\a[29] ), .out0(new_n278));
  nano22aa1n03x5               g183(.a(new_n276), .b(new_n277), .c(new_n278), .out0(new_n279));
  aoai13aa1n02x5               g184(.a(new_n275), .b(new_n271), .c(new_n179), .d(new_n258), .o1(new_n280));
  aoi012aa1n02x5               g185(.a(new_n278), .b(new_n280), .c(new_n277), .o1(new_n281));
  norp02aa1n03x5               g186(.a(new_n281), .b(new_n279), .o1(\s[29] ));
  xorb03aa1n02x5               g187(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g188(.a(new_n262), .b(new_n278), .c(new_n267), .out0(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n259), .c(new_n261), .out0(new_n285));
  oao003aa1n02x5               g190(.a(\a[29] ), .b(\b[28] ), .c(new_n277), .carry(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[29] ), .b(\a[30] ), .out0(new_n287));
  nano22aa1n03x7               g192(.a(new_n285), .b(new_n286), .c(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n284), .b(new_n271), .c(new_n179), .d(new_n258), .o1(new_n289));
  tech160nm_fiaoi012aa1n02p5x5 g194(.a(new_n287), .b(new_n289), .c(new_n286), .o1(new_n290));
  nor002aa1n02x5               g195(.a(new_n290), .b(new_n288), .o1(\s[30] ));
  norb02aa1n02x5               g196(.a(new_n284), .b(new_n287), .out0(new_n292));
  aobi12aa1n03x5               g197(.a(new_n292), .b(new_n259), .c(new_n261), .out0(new_n293));
  oao003aa1n02x5               g198(.a(\a[30] ), .b(\b[29] ), .c(new_n286), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[30] ), .b(\a[31] ), .out0(new_n295));
  nano22aa1n03x5               g200(.a(new_n293), .b(new_n294), .c(new_n295), .out0(new_n296));
  aoai13aa1n02x5               g201(.a(new_n292), .b(new_n271), .c(new_n179), .d(new_n258), .o1(new_n297));
  aoi012aa1n02x5               g202(.a(new_n295), .b(new_n297), .c(new_n294), .o1(new_n298));
  norp02aa1n03x5               g203(.a(new_n298), .b(new_n296), .o1(\s[31] ));
  xnrb03aa1n02x5               g204(.a(new_n110), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g205(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n301));
  xorb03aa1n02x5               g206(.a(new_n301), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g207(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g208(.a(\b[4] ), .o1(new_n304));
  oaoi03aa1n02x5               g209(.a(new_n113), .b(new_n304), .c(new_n112), .o1(new_n305));
  xorb03aa1n02x5               g210(.a(new_n305), .b(\b[5] ), .c(new_n114), .out0(\s[6] ));
  aob012aa1n02x5               g211(.a(new_n118), .b(new_n112), .c(new_n115), .out0(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g213(.a(new_n100), .b(new_n307), .out0(new_n309));
  xobna2aa1n03x5               g214(.a(new_n99), .b(new_n309), .c(new_n119), .out0(\s[8] ));
  xnbna2aa1n03x5               g215(.a(new_n123), .b(new_n116), .c(new_n121), .out0(\s[9] ));
endmodule


