// Benchmark "adder" written by ABC on Wed Jul 17 16:56:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n322, new_n323, new_n326,
    new_n328, new_n330, new_n331, new_n332, new_n334, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n02p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\a[9] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\b[8] ), .b(new_n98), .out0(new_n99));
  nor042aa1n06x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand02aa1d16x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand02aa1d24x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  aoi012aa1d18x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand02aa1n08x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n06x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  xorc02aa1n12x5               g011(.a(\a[3] ), .b(\b[2] ), .out0(new_n107));
  nanb03aa1n12x5               g012(.a(new_n103), .b(new_n107), .c(new_n106), .out0(new_n108));
  nor002aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  aoi012aa1n09x5               g014(.a(new_n104), .b(new_n109), .c(new_n105), .o1(new_n110));
  xorc02aa1n06x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  inv000aa1d42x5               g016(.a(\b[6] ), .o1(new_n112));
  nanb02aa1d36x5               g017(.a(\a[7] ), .b(new_n112), .out0(new_n113));
  nand02aa1d24x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(new_n113), .b(new_n114), .o1(new_n115));
  nand02aa1d08x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor002aa1d32x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nanb02aa1n03x5               g022(.a(new_n117), .b(new_n116), .out0(new_n118));
  xorc02aa1n12x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nona23aa1n09x5               g024(.a(new_n111), .b(new_n119), .c(new_n118), .d(new_n115), .out0(new_n120));
  norp02aa1n02x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nor042aa1d18x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  tech160nm_fioai012aa1n03p5x5 g027(.a(new_n116), .b(new_n122), .c(new_n117), .o1(new_n123));
  nanp02aa1n03x5               g028(.a(new_n123), .b(new_n113), .o1(new_n124));
  aoi022aa1n02x7               g029(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n125));
  aoi012aa1n06x5               g030(.a(new_n121), .b(new_n124), .c(new_n125), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n126), .b(new_n120), .c(new_n108), .d(new_n110), .o1(new_n127));
  tech160nm_fixorc02aa1n03p5x5 g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  nanp02aa1n02x5               g033(.a(new_n127), .b(new_n128), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  nand42aa1n08x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor042aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nanb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  oa0022aa1n06x5               g038(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n134));
  nand22aa1n03x5               g039(.a(new_n129), .b(new_n134), .o1(new_n135));
  aob012aa1n02x5               g040(.a(new_n135), .b(\b[9] ), .c(\a[10] ), .out0(new_n136));
  nand42aa1n03x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nano22aa1n09x5               g042(.a(new_n132), .b(new_n137), .c(new_n131), .out0(new_n138));
  aoi022aa1n02x5               g043(.a(new_n136), .b(new_n133), .c(new_n135), .d(new_n138), .o1(\s[11] ));
  nor042aa1n06x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1n06x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanb02aa1n03x5               g046(.a(new_n140), .b(new_n141), .out0(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n132), .c(new_n135), .d(new_n138), .o1(new_n143));
  aoi112aa1n03x5               g048(.a(new_n142), .b(new_n132), .c(new_n135), .d(new_n138), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(\s[12] ));
  nano23aa1n02x5               g050(.a(new_n140), .b(new_n132), .c(new_n141), .d(new_n131), .out0(new_n146));
  and003aa1n02x5               g051(.a(new_n146), .b(new_n128), .c(new_n97), .o(new_n147));
  nanp02aa1n02x5               g052(.a(new_n127), .b(new_n147), .o1(new_n148));
  nona22aa1n09x5               g053(.a(new_n138), .b(new_n142), .c(new_n134), .out0(new_n149));
  tech160nm_fiaoi012aa1n05x5   g054(.a(new_n140), .b(new_n132), .c(new_n141), .o1(new_n150));
  nand02aa1d06x5               g055(.a(new_n149), .b(new_n150), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(new_n148), .b(new_n152), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g059(.a(\a[14] ), .o1(new_n155));
  inv000aa1d42x5               g060(.a(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(\b[12] ), .o1(new_n157));
  oaoi03aa1n02x5               g062(.a(new_n156), .b(new_n157), .c(new_n153), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(new_n155), .out0(\s[14] ));
  nor002aa1n02x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand02aa1n03x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nor002aa1d32x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand42aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nano23aa1n03x7               g068(.a(new_n160), .b(new_n162), .c(new_n163), .d(new_n161), .out0(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n151), .c(new_n127), .d(new_n147), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n163), .b(new_n162), .c(new_n156), .d(new_n157), .o1(new_n166));
  nor042aa1n02x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nand42aa1n06x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n165), .c(new_n166), .out0(\s[15] ));
  nand22aa1n03x5               g075(.a(new_n165), .b(new_n166), .o1(new_n171));
  nor042aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand42aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  aoai13aa1n03x5               g079(.a(new_n174), .b(new_n167), .c(new_n171), .d(new_n168), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n171), .b(new_n169), .o1(new_n176));
  nona22aa1n02x4               g081(.a(new_n176), .b(new_n174), .c(new_n167), .out0(new_n177));
  nanp02aa1n02x5               g082(.a(new_n177), .b(new_n175), .o1(\s[16] ));
  nano23aa1n02x5               g083(.a(new_n167), .b(new_n172), .c(new_n173), .d(new_n168), .out0(new_n179));
  nand02aa1n03x5               g084(.a(new_n179), .b(new_n164), .o1(new_n180));
  nano32aa1n03x7               g085(.a(new_n180), .b(new_n146), .c(new_n128), .d(new_n97), .out0(new_n181));
  nand02aa1d06x5               g086(.a(new_n127), .b(new_n181), .o1(new_n182));
  nanb02aa1n02x5               g087(.a(new_n167), .b(new_n166), .out0(new_n183));
  aoi022aa1n02x5               g088(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n184));
  tech160nm_fiaoi012aa1n03p5x5 g089(.a(new_n172), .b(new_n183), .c(new_n184), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n185), .b(new_n180), .c(new_n149), .d(new_n150), .o1(new_n186));
  inv000aa1n06x5               g091(.a(new_n186), .o1(new_n187));
  nor042aa1d18x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  nand42aa1d28x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  norb02aa1n02x5               g094(.a(new_n189), .b(new_n188), .out0(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n190), .b(new_n182), .c(new_n187), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[18] ), .o1(new_n192));
  nand22aa1n09x5               g097(.a(new_n182), .b(new_n187), .o1(new_n193));
  tech160nm_fiaoi012aa1n05x5   g098(.a(new_n188), .b(new_n193), .c(new_n190), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  nor002aa1d32x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nand42aa1d28x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nano23aa1d15x5               g102(.a(new_n188), .b(new_n196), .c(new_n197), .d(new_n189), .out0(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n186), .c(new_n127), .d(new_n181), .o1(new_n199));
  oa0012aa1n02x5               g104(.a(new_n197), .b(new_n196), .c(new_n188), .o(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  nor042aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1d08x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n15x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n199), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n05x5   g111(.a(new_n199), .b(new_n201), .o1(new_n207));
  nor042aa1n12x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1n20x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n12x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n202), .c(new_n207), .d(new_n203), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(new_n207), .b(new_n204), .o1(new_n212));
  nona22aa1n02x4               g117(.a(new_n212), .b(new_n210), .c(new_n202), .out0(new_n213));
  nanp02aa1n02x5               g118(.a(new_n213), .b(new_n211), .o1(\s[20] ));
  nanb03aa1d24x5               g119(.a(new_n210), .b(new_n198), .c(new_n204), .out0(new_n215));
  nanb03aa1d24x5               g120(.a(new_n208), .b(new_n209), .c(new_n203), .out0(new_n216));
  orn002aa1n03x5               g121(.a(\a[19] ), .b(\b[18] ), .o(new_n217));
  oai112aa1n06x5               g122(.a(new_n217), .b(new_n197), .c(new_n196), .d(new_n188), .o1(new_n218));
  aoi012aa1d24x5               g123(.a(new_n208), .b(new_n202), .c(new_n209), .o1(new_n219));
  oai012aa1d24x5               g124(.a(new_n219), .b(new_n218), .c(new_n216), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n215), .c(new_n182), .d(new_n187), .o1(new_n222));
  nor042aa1n04x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n215), .o1(new_n226));
  aoi112aa1n02x5               g131(.a(new_n225), .b(new_n220), .c(new_n193), .d(new_n226), .o1(new_n227));
  aoi012aa1n02x5               g132(.a(new_n227), .b(new_n222), .c(new_n225), .o1(\s[21] ));
  nor042aa1n03x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  nand02aa1n06x5               g134(.a(\b[21] ), .b(\a[22] ), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(new_n229), .b(new_n230), .out0(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n223), .c(new_n222), .d(new_n225), .o1(new_n232));
  nand42aa1n02x5               g137(.a(new_n222), .b(new_n225), .o1(new_n233));
  nona22aa1n02x4               g138(.a(new_n233), .b(new_n231), .c(new_n223), .out0(new_n234));
  nanp02aa1n03x5               g139(.a(new_n234), .b(new_n232), .o1(\s[22] ));
  nano23aa1n09x5               g140(.a(new_n223), .b(new_n229), .c(new_n230), .d(new_n224), .out0(new_n236));
  nanb02aa1n02x5               g141(.a(new_n215), .b(new_n236), .out0(new_n237));
  aoi012aa1d18x5               g142(.a(new_n229), .b(new_n223), .c(new_n230), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n220), .c(new_n236), .o1(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n237), .c(new_n182), .d(new_n187), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  xnrc02aa1n12x5               g149(.a(\b[23] ), .b(\a[24] ), .out0(new_n245));
  aoai13aa1n03x5               g150(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n246));
  nand42aa1n02x5               g151(.a(new_n241), .b(new_n244), .o1(new_n247));
  nona22aa1n03x5               g152(.a(new_n247), .b(new_n245), .c(new_n243), .out0(new_n248));
  nanp02aa1n03x5               g153(.a(new_n248), .b(new_n246), .o1(\s[24] ));
  norb02aa1n06x4               g154(.a(new_n244), .b(new_n245), .out0(new_n250));
  nano22aa1n03x7               g155(.a(new_n215), .b(new_n250), .c(new_n236), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n186), .c(new_n127), .d(new_n181), .o1(new_n252));
  nano22aa1n03x5               g157(.a(new_n208), .b(new_n203), .c(new_n209), .out0(new_n253));
  oai012aa1n02x5               g158(.a(new_n197), .b(\b[18] ), .c(\a[19] ), .o1(new_n254));
  oab012aa1n02x4               g159(.a(new_n254), .b(new_n188), .c(new_n196), .out0(new_n255));
  inv040aa1n03x5               g160(.a(new_n219), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n236), .b(new_n256), .c(new_n255), .d(new_n253), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n250), .o1(new_n258));
  aoi112aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n259));
  oab012aa1n02x4               g164(.a(new_n259), .b(\a[24] ), .c(\b[23] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n258), .c(new_n257), .d(new_n238), .o1(new_n261));
  nanb02aa1n03x5               g166(.a(new_n261), .b(new_n252), .out0(new_n262));
  xorb03aa1n02x5               g167(.a(new_n262), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[25] ), .b(\b[24] ), .out0(new_n265));
  xnrc02aa1n12x5               g170(.a(\b[25] ), .b(\a[26] ), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n266), .b(new_n264), .c(new_n262), .d(new_n265), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n265), .b(new_n261), .c(new_n193), .d(new_n251), .o1(new_n268));
  nona22aa1n03x5               g173(.a(new_n268), .b(new_n266), .c(new_n264), .out0(new_n269));
  nanp02aa1n03x5               g174(.a(new_n267), .b(new_n269), .o1(\s[26] ));
  norb02aa1n12x5               g175(.a(new_n265), .b(new_n266), .out0(new_n271));
  inv030aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  nano23aa1d12x5               g177(.a(new_n272), .b(new_n215), .c(new_n250), .d(new_n236), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n186), .c(new_n127), .d(new_n181), .o1(new_n274));
  inv000aa1d42x5               g179(.a(\a[26] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(\b[25] ), .o1(new_n276));
  oaoi03aa1n02x5               g181(.a(new_n275), .b(new_n276), .c(new_n264), .o1(new_n277));
  inv000aa1n02x5               g182(.a(new_n277), .o1(new_n278));
  aoi012aa1n09x5               g183(.a(new_n278), .b(new_n261), .c(new_n271), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[27] ), .b(\b[26] ), .out0(new_n280));
  xnbna2aa1n03x5               g185(.a(new_n280), .b(new_n279), .c(new_n274), .out0(\s[27] ));
  tech160nm_finand02aa1n03p5x5 g186(.a(new_n279), .b(new_n274), .o1(new_n282));
  norp02aa1n02x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  nor002aa1n02x5               g188(.a(\b[27] ), .b(\a[28] ), .o1(new_n284));
  nand42aa1n06x5               g189(.a(\b[27] ), .b(\a[28] ), .o1(new_n285));
  nanb02aa1n12x5               g190(.a(new_n284), .b(new_n285), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n282), .d(new_n280), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n250), .b(new_n239), .c(new_n220), .d(new_n236), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n277), .b(new_n272), .c(new_n288), .d(new_n260), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n280), .b(new_n289), .c(new_n193), .d(new_n273), .o1(new_n290));
  nona22aa1n02x4               g195(.a(new_n290), .b(new_n286), .c(new_n283), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n287), .b(new_n291), .o1(\s[28] ));
  norb02aa1n03x5               g197(.a(new_n280), .b(new_n286), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n193), .d(new_n273), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n293), .o1(new_n295));
  oai012aa1n02x5               g200(.a(new_n285), .b(new_n284), .c(new_n283), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n295), .c(new_n279), .d(new_n274), .o1(new_n297));
  norp02aa1n02x5               g202(.a(\b[28] ), .b(\a[29] ), .o1(new_n298));
  nand42aa1n03x5               g203(.a(\b[28] ), .b(\a[29] ), .o1(new_n299));
  norb02aa1n02x5               g204(.a(new_n299), .b(new_n298), .out0(new_n300));
  oai022aa1n02x5               g205(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n301));
  aboi22aa1n03x5               g206(.a(new_n298), .b(new_n299), .c(new_n301), .d(new_n285), .out0(new_n302));
  aoi022aa1n03x5               g207(.a(new_n297), .b(new_n300), .c(new_n294), .d(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d21x5               g209(.a(new_n286), .b(new_n280), .c(new_n300), .out0(new_n305));
  aoai13aa1n06x5               g210(.a(new_n305), .b(new_n289), .c(new_n193), .d(new_n273), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n305), .o1(new_n307));
  aoi013aa1n02x4               g212(.a(new_n298), .b(new_n301), .c(new_n285), .d(new_n299), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n307), .c(new_n279), .d(new_n274), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .out0(new_n310));
  aoi113aa1n02x5               g215(.a(new_n310), .b(new_n298), .c(new_n301), .d(new_n299), .e(new_n285), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n306), .d(new_n311), .o1(\s[30] ));
  nand23aa1n04x5               g217(.a(new_n293), .b(new_n300), .c(new_n310), .o1(new_n313));
  nanb02aa1n03x5               g218(.a(new_n313), .b(new_n282), .out0(new_n314));
  xorc02aa1n02x5               g219(.a(\a[31] ), .b(\b[30] ), .out0(new_n315));
  oao003aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n316));
  norb02aa1n02x5               g221(.a(new_n316), .b(new_n315), .out0(new_n317));
  aoai13aa1n02x7               g222(.a(new_n316), .b(new_n313), .c(new_n279), .d(new_n274), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n314), .b(new_n317), .c(new_n318), .d(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n06x5               g225(.a(new_n108), .b(new_n110), .o1(new_n321));
  obai22aa1n02x7               g226(.a(new_n105), .b(new_n104), .c(\a[3] ), .d(\b[2] ), .out0(new_n322));
  aoib12aa1n02x5               g227(.a(new_n322), .b(new_n107), .c(new_n103), .out0(new_n323));
  oaoi13aa1n02x5               g228(.a(new_n323), .b(new_n321), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g229(.a(new_n119), .b(new_n108), .c(new_n110), .out0(\s[5] ));
  tech160nm_fiao0012aa1n03p5x5 g230(.a(new_n122), .b(new_n321), .c(new_n119), .o(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiaoi012aa1n04x5   g232(.a(new_n117), .b(new_n326), .c(new_n116), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n113), .c(new_n114), .out0(\s[7] ));
  inv000aa1d42x5               g234(.a(new_n114), .o1(new_n330));
  aoi112aa1n02x5               g235(.a(new_n330), .b(new_n111), .c(new_n328), .d(new_n113), .o1(new_n331));
  aoai13aa1n02x5               g236(.a(new_n111), .b(new_n330), .c(new_n328), .d(new_n113), .o1(new_n332));
  nanb02aa1n02x5               g237(.a(new_n331), .b(new_n332), .out0(\s[8] ));
  aoi112aa1n02x5               g238(.a(new_n128), .b(new_n121), .c(new_n124), .d(new_n125), .o1(new_n334));
  aoai13aa1n02x5               g239(.a(new_n334), .b(new_n120), .c(new_n108), .d(new_n110), .o1(new_n335));
  aobi12aa1n02x5               g240(.a(new_n335), .b(new_n128), .c(new_n127), .out0(\s[9] ));
endmodule


