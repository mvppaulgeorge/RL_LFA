// Benchmark "adder" written by ABC on Wed Jul 17 14:02:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n316, new_n318, new_n319, new_n321;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[8] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[4] ), .o1(new_n100));
  inv040aa1d32x5               g005(.a(\a[3] ), .o1(new_n101));
  inv040aa1d28x5               g006(.a(\b[2] ), .o1(new_n102));
  nanp02aa1n09x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand22aa1n04x5               g009(.a(new_n103), .b(new_n104), .o1(new_n105));
  nor042aa1n06x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nand42aa1n20x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nand42aa1d28x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  aoi012aa1n12x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  aboi22aa1d24x5               g014(.a(\b[3] ), .b(new_n100), .c(new_n101), .d(new_n102), .out0(new_n110));
  tech160nm_fioai012aa1n05x5   g015(.a(new_n110), .b(new_n109), .c(new_n105), .o1(new_n111));
  oaib12aa1n09x5               g016(.a(new_n111), .b(new_n100), .c(\b[3] ), .out0(new_n112));
  norp02aa1n12x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand22aa1n12x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor022aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand02aa1n06x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1d18x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  tech160nm_fixnrc02aa1n02p5x5 g022(.a(\b[5] ), .b(\a[6] ), .out0(new_n118));
  tech160nm_fixorc02aa1n05x5   g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nona22aa1n03x5               g024(.a(new_n119), .b(new_n117), .c(new_n118), .out0(new_n120));
  inv000aa1d42x5               g025(.a(\b[5] ), .o1(new_n121));
  oaih22aa1n06x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  oaib12aa1n12x5               g027(.a(new_n122), .b(new_n121), .c(\a[6] ), .out0(new_n123));
  ao0012aa1n03x7               g028(.a(new_n113), .b(new_n115), .c(new_n114), .o(new_n124));
  oabi12aa1n18x5               g029(.a(new_n124), .b(new_n117), .c(new_n123), .out0(new_n125));
  oabi12aa1n18x5               g030(.a(new_n125), .b(new_n120), .c(new_n112), .out0(new_n126));
  oaib12aa1n06x5               g031(.a(new_n126), .b(new_n99), .c(\a[9] ), .out0(new_n127));
  norb02aa1n03x5               g032(.a(new_n127), .b(new_n98), .out0(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  and002aa1n12x5               g034(.a(\b[9] ), .b(\a[10] ), .o(new_n130));
  nor042aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  and002aa1n02x5               g036(.a(\b[10] ), .b(\a[11] ), .o(new_n132));
  oai122aa1n06x5               g037(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .d(\b[8] ), .e(\a[9] ), .o1(new_n133));
  nona32aa1n03x5               g038(.a(new_n133), .b(new_n132), .c(new_n131), .d(new_n130), .out0(new_n134));
  inv030aa1n06x5               g039(.a(new_n131), .o1(new_n135));
  nand42aa1d28x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  aboi22aa1n03x5               g041(.a(new_n130), .b(new_n133), .c(new_n135), .d(new_n136), .out0(new_n137));
  norb02aa1n03x4               g042(.a(new_n134), .b(new_n137), .out0(\s[11] ));
  nor042aa1n12x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand42aa1d28x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  nona22aa1n03x5               g046(.a(new_n134), .b(new_n141), .c(new_n131), .out0(new_n142));
  aobi12aa1n06x5               g047(.a(new_n141), .b(new_n134), .c(new_n135), .out0(new_n143));
  norb02aa1n03x4               g048(.a(new_n142), .b(new_n143), .out0(\s[12] ));
  xnrc02aa1n12x5               g049(.a(\b[12] ), .b(\a[13] ), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  nona23aa1n09x5               g051(.a(new_n140), .b(new_n136), .c(new_n131), .d(new_n139), .out0(new_n147));
  oai022aa1n04x7               g052(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n148));
  nanb02aa1n09x5               g053(.a(new_n130), .b(new_n148), .out0(new_n149));
  oaoi03aa1n09x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n135), .o1(new_n150));
  oabi12aa1n18x5               g055(.a(new_n150), .b(new_n147), .c(new_n149), .out0(new_n151));
  inv040aa1n03x5               g056(.a(new_n151), .o1(new_n152));
  and002aa1n02x5               g057(.a(\b[3] ), .b(\a[4] ), .o(new_n153));
  oaoi13aa1n12x5               g058(.a(new_n153), .b(new_n110), .c(new_n109), .d(new_n105), .o1(new_n154));
  norb03aa1n03x5               g059(.a(new_n119), .b(new_n117), .c(new_n118), .out0(new_n155));
  xorc02aa1n12x5               g060(.a(\a[10] ), .b(\b[9] ), .out0(new_n156));
  nano23aa1n06x5               g061(.a(new_n131), .b(new_n139), .c(new_n140), .d(new_n136), .out0(new_n157));
  xorc02aa1n12x5               g062(.a(\a[9] ), .b(\b[8] ), .out0(new_n158));
  nand23aa1d12x5               g063(.a(new_n157), .b(new_n156), .c(new_n158), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  aoai13aa1n06x5               g065(.a(new_n160), .b(new_n125), .c(new_n154), .d(new_n155), .o1(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n146), .b(new_n161), .c(new_n152), .out0(\s[13] ));
  orn002aa1n03x5               g067(.a(\a[13] ), .b(\b[12] ), .o(new_n163));
  aoai13aa1n03x5               g068(.a(new_n163), .b(new_n145), .c(new_n161), .d(new_n152), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  tech160nm_fixnrc02aa1n02p5x5 g070(.a(\b[13] ), .b(\a[14] ), .out0(new_n166));
  nor042aa1n06x5               g071(.a(new_n166), .b(new_n145), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  oao003aa1n03x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .carry(new_n169));
  aoai13aa1n04x5               g074(.a(new_n169), .b(new_n168), .c(new_n161), .d(new_n152), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1d28x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nor042aa1n06x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand42aa1n20x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  aoi112aa1n02x5               g081(.a(new_n176), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n176), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n178), .b(new_n177), .out0(\s[16] ));
  nano23aa1d15x5               g084(.a(new_n172), .b(new_n174), .c(new_n175), .d(new_n173), .out0(new_n180));
  nona22aa1n09x5               g085(.a(new_n180), .b(new_n166), .c(new_n145), .out0(new_n181));
  nor042aa1n06x5               g086(.a(new_n181), .b(new_n159), .o1(new_n182));
  aoai13aa1n06x5               g087(.a(new_n182), .b(new_n125), .c(new_n154), .d(new_n155), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n174), .b(new_n172), .c(new_n175), .o1(new_n184));
  oaib12aa1n09x5               g089(.a(new_n184), .b(new_n169), .c(new_n180), .out0(new_n185));
  aoi013aa1n09x5               g090(.a(new_n185), .b(new_n151), .c(new_n167), .d(new_n180), .o1(new_n186));
  nand02aa1d08x5               g091(.a(new_n183), .b(new_n186), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[16] ), .o1(new_n191));
  oaoi03aa1n03x5               g096(.a(new_n190), .b(new_n191), .c(new_n187), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(new_n189), .out0(\s[18] ));
  xroi22aa1d06x4               g098(.a(new_n190), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n194));
  nand22aa1n09x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nona22aa1n02x4               g100(.a(new_n195), .b(\b[16] ), .c(\a[17] ), .out0(new_n196));
  oaib12aa1n06x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n189), .out0(new_n197));
  nor002aa1d32x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand22aa1n06x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n201));
  aoi112aa1n02x5               g106(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n202));
  norb02aa1n03x4               g107(.a(new_n201), .b(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand22aa1n09x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  nona22aa1n02x5               g112(.a(new_n201), .b(new_n207), .c(new_n198), .out0(new_n208));
  orn002aa1n02x5               g113(.a(\a[19] ), .b(\b[18] ), .o(new_n209));
  aobi12aa1n06x5               g114(.a(new_n207), .b(new_n201), .c(new_n209), .out0(new_n210));
  norb02aa1n03x4               g115(.a(new_n208), .b(new_n210), .out0(\s[20] ));
  nano23aa1n06x5               g116(.a(new_n198), .b(new_n205), .c(new_n206), .d(new_n199), .out0(new_n212));
  nanp02aa1n02x5               g117(.a(new_n194), .b(new_n212), .o1(new_n213));
  norp02aa1n04x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  aoi013aa1n06x4               g119(.a(new_n214), .b(new_n195), .c(new_n190), .d(new_n191), .o1(new_n215));
  nona23aa1d18x5               g120(.a(new_n206), .b(new_n199), .c(new_n198), .d(new_n205), .out0(new_n216));
  aoi012aa1n12x5               g121(.a(new_n205), .b(new_n198), .c(new_n206), .o1(new_n217));
  oai012aa1n18x5               g122(.a(new_n217), .b(new_n216), .c(new_n215), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n06x5               g124(.a(new_n219), .b(new_n213), .c(new_n183), .d(new_n186), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[21] ), .b(\b[20] ), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[22] ), .b(\b[21] ), .out0(new_n224));
  aoi112aa1n02x5               g129(.a(new_n222), .b(new_n224), .c(new_n220), .d(new_n223), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n224), .b(new_n222), .c(new_n220), .d(new_n223), .o1(new_n226));
  norb02aa1n02x7               g131(.a(new_n226), .b(new_n225), .out0(\s[22] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(\b[21] ), .o1(new_n231));
  oaoi03aa1n12x5               g136(.a(new_n229), .b(new_n231), .c(new_n222), .o1(new_n232));
  inv000aa1n02x5               g137(.a(new_n232), .o1(new_n233));
  aoi012aa1n02x5               g138(.a(new_n233), .b(new_n218), .c(new_n230), .o1(new_n234));
  nanp03aa1n02x5               g139(.a(new_n230), .b(new_n194), .c(new_n212), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n234), .b(new_n235), .c(new_n183), .d(new_n186), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  xorc02aa1n02x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xorc02aa1n02x5               g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  aoi112aa1n02x5               g145(.a(new_n238), .b(new_n240), .c(new_n236), .d(new_n239), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n238), .c(new_n236), .d(new_n239), .o1(new_n242));
  norb02aa1n02x7               g147(.a(new_n242), .b(new_n241), .out0(\s[24] ));
  inv000aa1d42x5               g148(.a(\a[23] ), .o1(new_n244));
  inv040aa1d32x5               g149(.a(\a[24] ), .o1(new_n245));
  xroi22aa1d06x4               g150(.a(new_n244), .b(\b[22] ), .c(new_n245), .d(\b[23] ), .out0(new_n246));
  nano22aa1n02x4               g151(.a(new_n213), .b(new_n230), .c(new_n246), .out0(new_n247));
  inv000aa1n02x5               g152(.a(new_n217), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n230), .b(new_n248), .c(new_n212), .d(new_n197), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n246), .o1(new_n250));
  aoi112aa1n02x5               g155(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n251));
  aoib12aa1n02x5               g156(.a(new_n251), .b(new_n245), .c(\b[23] ), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n250), .c(new_n249), .d(new_n232), .o1(new_n253));
  xorc02aa1n02x5               g158(.a(\a[25] ), .b(\b[24] ), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n253), .c(new_n187), .d(new_n247), .o1(new_n255));
  aoi112aa1n02x5               g160(.a(new_n254), .b(new_n253), .c(new_n187), .d(new_n247), .o1(new_n256));
  norb02aa1n03x4               g161(.a(new_n255), .b(new_n256), .out0(\s[25] ));
  norp02aa1n02x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  xorc02aa1n02x5               g163(.a(\a[26] ), .b(\b[25] ), .out0(new_n259));
  nona22aa1n02x5               g164(.a(new_n255), .b(new_n259), .c(new_n258), .out0(new_n260));
  inv000aa1n02x5               g165(.a(new_n258), .o1(new_n261));
  aobi12aa1n06x5               g166(.a(new_n259), .b(new_n255), .c(new_n261), .out0(new_n262));
  norb02aa1n03x4               g167(.a(new_n260), .b(new_n262), .out0(\s[26] ));
  oabi12aa1n03x5               g168(.a(new_n185), .b(new_n152), .c(new_n181), .out0(new_n264));
  inv000aa1d42x5               g169(.a(\a[25] ), .o1(new_n265));
  inv020aa1n04x5               g170(.a(\a[26] ), .o1(new_n266));
  xroi22aa1d06x4               g171(.a(new_n265), .b(\b[24] ), .c(new_n266), .d(\b[25] ), .out0(new_n267));
  nano32aa1n03x7               g172(.a(new_n213), .b(new_n267), .c(new_n230), .d(new_n246), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n264), .c(new_n126), .d(new_n182), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .c(new_n261), .carry(new_n270));
  aobi12aa1n06x5               g175(.a(new_n270), .b(new_n253), .c(new_n267), .out0(new_n271));
  nor042aa1n03x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  norb02aa1n02x5               g178(.a(new_n273), .b(new_n272), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n271), .c(new_n269), .out0(\s[27] ));
  inv000aa1n06x5               g180(.a(new_n272), .o1(new_n276));
  xnrc02aa1n02x5               g181(.a(\b[27] ), .b(\a[28] ), .out0(new_n277));
  aobi12aa1n06x5               g182(.a(new_n268), .b(new_n183), .c(new_n186), .out0(new_n278));
  aoai13aa1n02x5               g183(.a(new_n246), .b(new_n233), .c(new_n218), .d(new_n230), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n267), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n270), .b(new_n280), .c(new_n279), .d(new_n252), .o1(new_n281));
  oaih12aa1n02x5               g186(.a(new_n273), .b(new_n281), .c(new_n278), .o1(new_n282));
  tech160nm_fiaoi012aa1n02p5x5 g187(.a(new_n277), .b(new_n282), .c(new_n276), .o1(new_n283));
  aobi12aa1n02x7               g188(.a(new_n273), .b(new_n271), .c(new_n269), .out0(new_n284));
  nano22aa1n02x4               g189(.a(new_n284), .b(new_n276), .c(new_n277), .out0(new_n285));
  norp02aa1n03x5               g190(.a(new_n283), .b(new_n285), .o1(\s[28] ));
  nano22aa1n02x4               g191(.a(new_n277), .b(new_n276), .c(new_n273), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n281), .c(new_n278), .o1(new_n288));
  oao003aa1n03x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n276), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[28] ), .b(\a[29] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  aobi12aa1n02x7               g196(.a(new_n287), .b(new_n271), .c(new_n269), .out0(new_n292));
  nano22aa1n02x4               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g200(.a(new_n274), .b(new_n290), .c(new_n277), .out0(new_n296));
  oaih12aa1n02x5               g201(.a(new_n296), .b(new_n281), .c(new_n278), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[29] ), .b(\a[30] ), .out0(new_n299));
  tech160nm_fiaoi012aa1n02p5x5 g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n296), .b(new_n271), .c(new_n269), .out0(new_n301));
  nano22aa1n02x4               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[30] ));
  norb03aa1n02x5               g208(.a(new_n287), .b(new_n299), .c(new_n290), .out0(new_n304));
  aobi12aa1n02x7               g209(.a(new_n304), .b(new_n271), .c(new_n269), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  nano22aa1n02x4               g212(.a(new_n305), .b(new_n306), .c(new_n307), .out0(new_n308));
  oaih12aa1n02x5               g213(.a(new_n304), .b(new_n281), .c(new_n278), .o1(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n307), .b(new_n309), .c(new_n306), .o1(new_n310));
  norp02aa1n03x5               g215(.a(new_n310), .b(new_n308), .o1(\s[31] ));
  xnbna2aa1n03x5               g216(.a(new_n109), .b(new_n103), .c(new_n104), .out0(\s[3] ));
  oaoi03aa1n02x5               g217(.a(\a[3] ), .b(\b[2] ), .c(new_n109), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g219(.a(new_n154), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g220(.a(\a[5] ), .b(\b[4] ), .c(new_n112), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g222(.a(\a[6] ), .o1(new_n318));
  oaoi03aa1n03x5               g223(.a(new_n318), .b(new_n121), .c(new_n316), .o1(new_n319));
  xnrb03aa1n02x5               g224(.a(new_n319), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g225(.a(\a[7] ), .b(\b[6] ), .c(new_n319), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g227(.a(new_n126), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


