// Benchmark "adder" written by ABC on Wed Jul 17 23:00:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n328, new_n330, new_n331,
    new_n333, new_n335, new_n337, new_n338, new_n339, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1n06x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  nor042aa1n03x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nanp02aa1n06x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  tech160nm_fiaoi012aa1n03p5x5 g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  norb02aa1n06x4               g008(.a(new_n101), .b(new_n100), .out0(new_n104));
  nanp02aa1n12x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano22aa1n02x4               g011(.a(new_n102), .b(new_n105), .c(new_n106), .out0(new_n107));
  nand02aa1n03x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  nona22aa1n02x4               g014(.a(new_n105), .b(new_n109), .c(new_n108), .out0(new_n110));
  nanp03aa1n06x5               g015(.a(new_n107), .b(new_n110), .c(new_n104), .o1(new_n111));
  nor042aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor002aa1n03x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nanp02aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  xorc02aa1n02x5               g021(.a(\a[6] ), .b(\b[5] ), .out0(new_n117));
  xorc02aa1n02x5               g022(.a(\a[5] ), .b(\b[4] ), .out0(new_n118));
  nand03aa1n02x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .o1(new_n119));
  nor042aa1n03x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  inv000aa1n02x5               g025(.a(new_n120), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  oa0012aa1n06x5               g027(.a(new_n113), .b(new_n114), .c(new_n112), .o(new_n123));
  tech160nm_fiaoi012aa1n03p5x5 g028(.a(new_n123), .b(new_n116), .c(new_n122), .o1(new_n124));
  aoai13aa1n12x5               g029(.a(new_n124), .b(new_n119), .c(new_n111), .d(new_n103), .o1(new_n125));
  aob012aa1n06x5               g030(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  and002aa1n24x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  inv000aa1d42x5               g033(.a(new_n97), .o1(new_n129));
  nona22aa1n06x5               g034(.a(new_n126), .b(new_n98), .c(new_n129), .out0(new_n130));
  nand02aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor002aa1n20x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nona23aa1n06x5               g037(.a(new_n130), .b(new_n131), .c(new_n132), .d(new_n128), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n128), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n132), .o1(new_n135));
  aoi022aa1n02x5               g040(.a(new_n130), .b(new_n134), .c(new_n135), .d(new_n131), .o1(new_n136));
  norb02aa1n02x7               g041(.a(new_n133), .b(new_n136), .out0(\s[11] ));
  nor042aa1n06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1n16x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoi113aa1n02x5               g045(.a(new_n140), .b(new_n132), .c(new_n130), .d(new_n131), .e(new_n134), .o1(new_n141));
  aobi12aa1n06x5               g046(.a(new_n140), .b(new_n133), .c(new_n135), .out0(new_n142));
  nor002aa1n02x5               g047(.a(new_n142), .b(new_n141), .o1(\s[12] ));
  nano23aa1d15x5               g048(.a(new_n138), .b(new_n132), .c(new_n139), .d(new_n131), .out0(new_n144));
  tech160nm_fixorc02aa1n04x5   g049(.a(\a[9] ), .b(\b[8] ), .out0(new_n145));
  nand23aa1d12x5               g050(.a(new_n144), .b(new_n97), .c(new_n145), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  nona23aa1n09x5               g052(.a(new_n131), .b(new_n139), .c(new_n138), .d(new_n132), .out0(new_n148));
  oai022aa1n02x5               g053(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n149));
  nanb02aa1n06x5               g054(.a(new_n128), .b(new_n149), .out0(new_n150));
  aoi012aa1d18x5               g055(.a(new_n138), .b(new_n132), .c(new_n139), .o1(new_n151));
  oai012aa1n09x5               g056(.a(new_n151), .b(new_n148), .c(new_n150), .o1(new_n152));
  xnrc02aa1n12x5               g057(.a(\b[12] ), .b(\a[13] ), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n152), .c(new_n125), .d(new_n147), .o1(new_n155));
  oai112aa1n02x5               g060(.a(new_n151), .b(new_n153), .c(new_n148), .d(new_n150), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n156), .b(new_n125), .c(new_n147), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n155), .b(new_n157), .out0(\s[13] ));
  nor002aa1n16x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nor042aa1n02x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nanb02aa1n06x5               g067(.a(new_n161), .b(new_n162), .out0(new_n163));
  nona32aa1n03x5               g068(.a(new_n125), .b(new_n163), .c(new_n153), .d(new_n146), .out0(new_n164));
  nor042aa1n06x5               g069(.a(new_n153), .b(new_n163), .o1(new_n165));
  aoi012aa1n02x5               g070(.a(new_n161), .b(new_n159), .c(new_n162), .o1(new_n166));
  inv020aa1n02x5               g071(.a(new_n166), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n152), .c(new_n165), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n161), .b(new_n164), .c(new_n168), .o1(new_n169));
  aoi013aa1n02x4               g074(.a(new_n169), .b(new_n155), .c(new_n163), .d(new_n160), .o1(\s[14] ));
  nor042aa1n04x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand42aa1n03x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n164), .c(new_n168), .out0(\s[15] ));
  nor042aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  aob012aa1n03x5               g080(.a(new_n173), .b(new_n164), .c(new_n168), .out0(new_n176));
  nand02aa1n08x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  oaib12aa1n03x5               g082(.a(new_n176), .b(new_n175), .c(new_n177), .out0(new_n178));
  nano23aa1d15x5               g083(.a(new_n171), .b(new_n175), .c(new_n177), .d(new_n172), .out0(new_n179));
  nano22aa1d15x5               g084(.a(new_n146), .b(new_n165), .c(new_n179), .out0(new_n180));
  oaoi03aa1n02x5               g085(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n181));
  inv000aa1n02x5               g086(.a(new_n151), .o1(new_n182));
  aoai13aa1n02x7               g087(.a(new_n165), .b(new_n182), .c(new_n144), .d(new_n181), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n179), .o1(new_n184));
  aoi012aa1n02x7               g089(.a(new_n184), .b(new_n183), .c(new_n166), .o1(new_n185));
  aoi012aa1d24x5               g090(.a(new_n175), .b(new_n171), .c(new_n177), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  aoi112aa1n06x5               g092(.a(new_n185), .b(new_n187), .c(new_n125), .d(new_n180), .o1(new_n188));
  oa0022aa1n03x5               g093(.a(new_n178), .b(new_n171), .c(new_n175), .d(new_n188), .o(\s[16] ));
  nanb02aa1n02x5               g094(.a(new_n100), .b(new_n101), .out0(new_n190));
  nanb03aa1n02x5               g095(.a(new_n102), .b(new_n106), .c(new_n105), .out0(new_n191));
  norb03aa1n03x5               g096(.a(new_n105), .b(new_n109), .c(new_n108), .out0(new_n192));
  oai013aa1n06x5               g097(.a(new_n103), .b(new_n192), .c(new_n191), .d(new_n190), .o1(new_n193));
  nona23aa1n02x4               g098(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n194));
  xnrc02aa1n02x5               g099(.a(\b[5] ), .b(\a[6] ), .out0(new_n195));
  norb03aa1n06x5               g100(.a(new_n118), .b(new_n194), .c(new_n195), .out0(new_n196));
  tech160nm_fiao0012aa1n02p5x5 g101(.a(new_n123), .b(new_n116), .c(new_n122), .o(new_n197));
  aoai13aa1n12x5               g102(.a(new_n180), .b(new_n197), .c(new_n193), .d(new_n196), .o1(new_n198));
  aoai13aa1n09x5               g103(.a(new_n179), .b(new_n167), .c(new_n152), .d(new_n165), .o1(new_n199));
  nanp03aa1d24x5               g104(.a(new_n198), .b(new_n199), .c(new_n186), .o1(new_n200));
  tech160nm_fixorc02aa1n04x5   g105(.a(\a[17] ), .b(\b[16] ), .out0(new_n201));
  norp03aa1n02x5               g106(.a(new_n185), .b(new_n187), .c(new_n201), .o1(new_n202));
  aoi022aa1n02x5               g107(.a(new_n200), .b(new_n201), .c(new_n202), .d(new_n198), .o1(\s[17] ));
  nor042aa1n02x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nor042aa1n02x5               g109(.a(\b[16] ), .b(\a[17] ), .o1(new_n205));
  nand22aa1n04x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  norb02aa1n03x5               g111(.a(new_n206), .b(new_n204), .out0(new_n207));
  aoi112aa1n02x5               g112(.a(new_n205), .b(new_n207), .c(new_n200), .d(new_n201), .o1(new_n208));
  and002aa1n02x5               g113(.a(new_n201), .b(new_n207), .o(new_n209));
  tech160nm_fiaoi012aa1n04x5   g114(.a(new_n204), .b(new_n205), .c(new_n206), .o1(new_n210));
  oaib12aa1n02x7               g115(.a(new_n210), .b(new_n188), .c(new_n209), .out0(new_n211));
  aoib12aa1n02x5               g116(.a(new_n208), .b(new_n211), .c(new_n204), .out0(\s[18] ));
  nor042aa1n09x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  inv000aa1n03x5               g120(.a(new_n210), .o1(new_n216));
  aoi112aa1n02x5               g121(.a(new_n215), .b(new_n216), .c(new_n200), .d(new_n209), .o1(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(new_n211), .c(new_n215), .o1(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g124(.a(new_n213), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n215), .b(new_n216), .c(new_n200), .d(new_n209), .o1(new_n221));
  nor002aa1n03x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand02aa1n08x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n223), .o1(new_n225));
  oai022aa1n02x5               g130(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n226));
  nona22aa1n02x5               g131(.a(new_n221), .b(new_n225), .c(new_n226), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n224), .c(new_n220), .d(new_n221), .o1(\s[20] ));
  nona23aa1n09x5               g133(.a(new_n223), .b(new_n214), .c(new_n213), .d(new_n222), .out0(new_n229));
  nano22aa1n12x5               g134(.a(new_n229), .b(new_n201), .c(new_n207), .out0(new_n230));
  oab012aa1n06x5               g135(.a(new_n225), .b(new_n213), .c(new_n222), .out0(new_n231));
  oabi12aa1n06x5               g136(.a(new_n231), .b(new_n229), .c(new_n210), .out0(new_n232));
  nor002aa1d32x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  nanp02aa1n02x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n232), .c(new_n200), .d(new_n230), .o1(new_n236));
  nano23aa1n06x5               g141(.a(new_n213), .b(new_n222), .c(new_n223), .d(new_n214), .out0(new_n237));
  aoi112aa1n02x5               g142(.a(new_n231), .b(new_n235), .c(new_n237), .d(new_n216), .o1(new_n238));
  aobi12aa1n02x5               g143(.a(new_n238), .b(new_n200), .c(new_n230), .out0(new_n239));
  norb02aa1n02x7               g144(.a(new_n236), .b(new_n239), .out0(\s[21] ));
  inv000aa1d42x5               g145(.a(new_n233), .o1(new_n241));
  xnrc02aa1n12x5               g146(.a(\b[21] ), .b(\a[22] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  and002aa1n02x5               g148(.a(\b[21] ), .b(\a[22] ), .o(new_n244));
  oai022aa1n02x5               g149(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n245));
  nona22aa1n02x5               g150(.a(new_n236), .b(new_n244), .c(new_n245), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n243), .c(new_n241), .d(new_n236), .o1(\s[22] ));
  nano22aa1n06x5               g152(.a(new_n242), .b(new_n241), .c(new_n234), .out0(new_n248));
  nand22aa1n09x5               g153(.a(new_n230), .b(new_n248), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n248), .b(new_n231), .c(new_n237), .d(new_n216), .o1(new_n251));
  oaoi03aa1n09x5               g156(.a(\a[22] ), .b(\b[21] ), .c(new_n241), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n251), .b(new_n253), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[22] ), .b(\a[23] ), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n254), .c(new_n200), .d(new_n250), .o1(new_n257));
  aoi112aa1n02x5               g162(.a(new_n256), .b(new_n254), .c(new_n200), .d(new_n250), .o1(new_n258));
  norb02aa1n03x4               g163(.a(new_n257), .b(new_n258), .out0(\s[23] ));
  norp02aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  and002aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .o(new_n263));
  oai022aa1n02x5               g168(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n264));
  nona22aa1n02x5               g169(.a(new_n257), .b(new_n263), .c(new_n264), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n262), .c(new_n261), .d(new_n257), .o1(\s[24] ));
  norb02aa1n09x5               g171(.a(new_n262), .b(new_n255), .out0(new_n267));
  and003aa1n02x5               g172(.a(new_n230), .b(new_n267), .c(new_n248), .o(new_n268));
  inv000aa1n02x5               g173(.a(new_n267), .o1(new_n269));
  aob012aa1n02x5               g174(.a(new_n264), .b(\b[23] ), .c(\a[24] ), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n251), .d(new_n253), .o1(new_n271));
  tech160nm_fixorc02aa1n03p5x5 g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n271), .c(new_n200), .d(new_n268), .o1(new_n273));
  aoi112aa1n02x5               g178(.a(new_n272), .b(new_n271), .c(new_n200), .d(new_n268), .o1(new_n274));
  norb02aa1n02x7               g179(.a(new_n273), .b(new_n274), .out0(\s[25] ));
  norp02aa1n02x5               g180(.a(\b[24] ), .b(\a[25] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[26] ), .b(\b[25] ), .out0(new_n278));
  and002aa1n02x5               g183(.a(\b[25] ), .b(\a[26] ), .o(new_n279));
  oai022aa1n02x5               g184(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n280));
  nona22aa1n02x5               g185(.a(new_n273), .b(new_n279), .c(new_n280), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n278), .c(new_n277), .d(new_n273), .o1(\s[26] ));
  and002aa1n06x5               g187(.a(new_n278), .b(new_n272), .o(new_n283));
  nano22aa1n09x5               g188(.a(new_n249), .b(new_n283), .c(new_n267), .out0(new_n284));
  inv020aa1n04x5               g189(.a(new_n284), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n279), .o1(new_n286));
  aoi022aa1n06x5               g191(.a(new_n271), .b(new_n283), .c(new_n286), .d(new_n280), .o1(new_n287));
  oaih12aa1n06x5               g192(.a(new_n287), .b(new_n188), .c(new_n285), .o1(new_n288));
  xorb03aa1n02x5               g193(.a(new_n288), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .out0(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n290), .c(new_n288), .d(new_n291), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n267), .b(new_n252), .c(new_n232), .d(new_n248), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n283), .o1(new_n295));
  aob012aa1n02x5               g200(.a(new_n280), .b(\b[25] ), .c(\a[26] ), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n295), .c(new_n294), .d(new_n270), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n291), .b(new_n297), .c(new_n200), .d(new_n284), .o1(new_n298));
  and002aa1n02x5               g203(.a(\b[27] ), .b(\a[28] ), .o(new_n299));
  oai022aa1n02x5               g204(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n300));
  nona22aa1n02x5               g205(.a(new_n298), .b(new_n299), .c(new_n300), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n293), .b(new_n301), .o1(\s[28] ));
  norb02aa1n02x5               g207(.a(new_n291), .b(new_n292), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n297), .c(new_n200), .d(new_n284), .o1(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[28] ), .b(\a[29] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n300), .b(new_n299), .out0(new_n306));
  nona22aa1n02x5               g211(.a(new_n304), .b(new_n305), .c(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n288), .d(new_n303), .o1(new_n308));
  nanp02aa1n03x5               g213(.a(new_n308), .b(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g215(.a(new_n291), .b(new_n305), .c(new_n292), .out0(new_n311));
  aob012aa1n02x5               g216(.a(new_n306), .b(\b[28] ), .c(\a[29] ), .out0(new_n312));
  oai012aa1n02x5               g217(.a(new_n312), .b(\b[28] ), .c(\a[29] ), .o1(new_n313));
  tech160nm_fixorc02aa1n02p5x5 g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n288), .d(new_n311), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n311), .b(new_n297), .c(new_n200), .d(new_n284), .o1(new_n317));
  nona22aa1n02x5               g222(.a(new_n317), .b(new_n313), .c(new_n315), .out0(new_n318));
  nanp02aa1n03x5               g223(.a(new_n316), .b(new_n318), .o1(\s[30] ));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nano23aa1n02x4               g225(.a(new_n305), .b(new_n292), .c(new_n314), .d(new_n291), .out0(new_n321));
  and002aa1n02x5               g226(.a(\b[29] ), .b(\a[30] ), .o(new_n322));
  oab012aa1n02x4               g227(.a(new_n322), .b(new_n313), .c(new_n315), .out0(new_n323));
  aoai13aa1n03x5               g228(.a(new_n320), .b(new_n323), .c(new_n288), .d(new_n321), .o1(new_n324));
  aoai13aa1n03x5               g229(.a(new_n321), .b(new_n297), .c(new_n200), .d(new_n284), .o1(new_n325));
  nona22aa1n02x5               g230(.a(new_n325), .b(new_n323), .c(new_n320), .out0(new_n326));
  nanp02aa1n03x5               g231(.a(new_n324), .b(new_n326), .o1(\s[31] ));
  norb02aa1n02x5               g232(.a(new_n106), .b(new_n102), .out0(new_n328));
  xobna2aa1n03x5               g233(.a(new_n328), .b(new_n110), .c(new_n105), .out0(\s[3] ));
  inv000aa1d42x5               g234(.a(new_n102), .o1(new_n330));
  oai112aa1n02x5               g235(.a(new_n328), .b(new_n105), .c(new_n108), .d(new_n109), .o1(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n104), .b(new_n331), .c(new_n330), .out0(\s[4] ));
  aoi112aa1n02x5               g237(.a(new_n118), .b(new_n100), .c(new_n101), .d(new_n102), .o1(new_n333));
  aoi022aa1n02x5               g238(.a(new_n193), .b(new_n118), .c(new_n111), .d(new_n333), .o1(\s[5] ));
  nanp02aa1n02x5               g239(.a(new_n193), .b(new_n118), .o1(new_n335));
  xnbna2aa1n03x5               g240(.a(new_n117), .b(new_n335), .c(new_n121), .out0(\s[6] ));
  nanb02aa1n02x5               g241(.a(new_n114), .b(new_n115), .out0(new_n337));
  nanp02aa1n02x5               g242(.a(\b[5] ), .b(\a[6] ), .o1(new_n338));
  nona22aa1n02x4               g243(.a(new_n335), .b(new_n120), .c(new_n195), .out0(new_n339));
  xnbna2aa1n03x5               g244(.a(new_n337), .b(new_n339), .c(new_n338), .out0(\s[7] ));
  aoi013aa1n02x4               g245(.a(new_n114), .b(new_n339), .c(new_n338), .d(new_n115), .o1(new_n341));
  xnrb03aa1n02x5               g246(.a(new_n341), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g247(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


