// Benchmark "adder" written by ABC on Wed Jul 17 19:07:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n326, new_n328, new_n330, new_n332, new_n333, new_n335,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n16x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor002aa1n10x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nona23aa1n09x5               g007(.a(new_n102), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n103));
  xorc02aa1n02x5               g008(.a(\a[5] ), .b(\b[4] ), .out0(new_n104));
  tech160nm_fixorc02aa1n02p5x5 g009(.a(\a[6] ), .b(\b[5] ), .out0(new_n105));
  nano22aa1n03x7               g010(.a(new_n103), .b(new_n104), .c(new_n105), .out0(new_n106));
  and002aa1n24x5               g011(.a(\b[3] ), .b(\a[4] ), .o(new_n107));
  norp02aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor002aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nor043aa1n02x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nanb02aa1n06x5               g016(.a(new_n109), .b(new_n111), .out0(new_n112));
  nor042aa1n02x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  tech160nm_fioai012aa1n05x5   g020(.a(new_n115), .b(new_n113), .c(new_n114), .o1(new_n116));
  oaoi13aa1n06x5               g021(.a(new_n107), .b(new_n110), .c(new_n116), .d(new_n112), .o1(new_n117));
  nor042aa1n03x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  inv000aa1n02x5               g023(.a(new_n118), .o1(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[6] ), .b(\b[5] ), .c(new_n119), .o1(new_n120));
  oai012aa1n02x5               g025(.a(new_n100), .b(new_n101), .c(new_n99), .o1(new_n121));
  oaib12aa1n02x5               g026(.a(new_n121), .b(new_n103), .c(new_n120), .out0(new_n122));
  xorc02aa1n12x5               g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  aoai13aa1n02x5               g028(.a(new_n123), .b(new_n122), .c(new_n117), .d(new_n106), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[10] ), .b(\b[9] ), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n125), .b(new_n124), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g031(.a(\a[5] ), .o1(new_n127));
  inv000aa1d42x5               g032(.a(\a[6] ), .o1(new_n128));
  xroi22aa1d04x5               g033(.a(new_n127), .b(\b[4] ), .c(new_n128), .d(\b[5] ), .out0(new_n129));
  tech160nm_fioai012aa1n03p5x5 g034(.a(new_n110), .b(new_n116), .c(new_n112), .o1(new_n130));
  nona23aa1n06x5               g035(.a(new_n130), .b(new_n129), .c(new_n103), .d(new_n107), .out0(new_n131));
  nona22aa1n02x4               g036(.a(new_n100), .b(new_n101), .c(new_n99), .out0(new_n132));
  aboi22aa1n03x5               g037(.a(new_n103), .b(new_n120), .c(new_n132), .d(new_n100), .out0(new_n133));
  nanp02aa1n02x5               g038(.a(new_n125), .b(new_n123), .o1(new_n134));
  norp02aa1n02x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  tech160nm_fioai012aa1n04x5   g041(.a(new_n136), .b(new_n135), .c(new_n97), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n137), .b(new_n134), .c(new_n131), .d(new_n133), .o1(new_n138));
  xorb03aa1n02x5               g043(.a(new_n138), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  orn002aa1n02x5               g044(.a(\a[11] ), .b(\b[10] ), .o(new_n140));
  nor022aa1n08x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nanp02aa1n09x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  nanp02aa1n02x5               g048(.a(new_n138), .b(new_n143), .o1(new_n144));
  norp02aa1n12x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand02aa1n06x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n140), .out0(\s[12] ));
  nanp02aa1n03x5               g053(.a(new_n131), .b(new_n133), .o1(new_n149));
  nano23aa1n06x5               g054(.a(new_n141), .b(new_n145), .c(new_n146), .d(new_n142), .out0(new_n150));
  nand23aa1d12x5               g055(.a(new_n150), .b(new_n123), .c(new_n125), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nona23aa1n03x5               g057(.a(new_n146), .b(new_n142), .c(new_n141), .d(new_n145), .out0(new_n153));
  oai012aa1n02x5               g058(.a(new_n146), .b(new_n145), .c(new_n141), .o1(new_n154));
  tech160nm_fioai012aa1n05x5   g059(.a(new_n154), .b(new_n153), .c(new_n137), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n155), .b(new_n149), .c(new_n152), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n02x5               g062(.a(\a[13] ), .b(\b[12] ), .c(new_n156), .o1(new_n158));
  nor002aa1n04x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nanp02aa1n04x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(new_n161));
  norp02aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand42aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  norb03aa1n02x5               g069(.a(new_n160), .b(new_n162), .c(new_n159), .out0(new_n165));
  oai012aa1n02x5               g070(.a(new_n165), .b(new_n156), .c(new_n164), .o1(new_n166));
  aob012aa1n02x5               g071(.a(new_n166), .b(new_n158), .c(new_n161), .out0(\s[14] ));
  nano23aa1n02x5               g072(.a(new_n162), .b(new_n159), .c(new_n160), .d(new_n163), .out0(new_n168));
  oaih12aa1n02x5               g073(.a(new_n160), .b(new_n159), .c(new_n162), .o1(new_n169));
  aobi12aa1n02x5               g074(.a(new_n169), .b(new_n155), .c(new_n168), .out0(new_n170));
  nona32aa1n02x4               g075(.a(new_n149), .b(new_n161), .c(new_n164), .d(new_n151), .out0(new_n171));
  nor042aa1n09x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand02aa1n06x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanb02aa1d24x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n171), .c(new_n170), .out0(\s[15] ));
  nanp02aa1n03x5               g081(.a(new_n171), .b(new_n170), .o1(new_n177));
  nor042aa1n02x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand42aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n03x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n172), .c(new_n177), .d(new_n175), .o1(new_n181));
  nona22aa1n02x4               g086(.a(new_n179), .b(new_n178), .c(new_n172), .out0(new_n182));
  aoai13aa1n02x5               g087(.a(new_n181), .b(new_n182), .c(new_n175), .d(new_n177), .o1(\s[16] ));
  nano23aa1n02x4               g088(.a(new_n172), .b(new_n178), .c(new_n179), .d(new_n173), .out0(new_n184));
  nano22aa1n03x7               g089(.a(new_n151), .b(new_n168), .c(new_n184), .out0(new_n185));
  aoai13aa1n06x5               g090(.a(new_n185), .b(new_n122), .c(new_n117), .d(new_n106), .o1(new_n186));
  nona23aa1n03x5               g091(.a(new_n160), .b(new_n163), .c(new_n162), .d(new_n159), .out0(new_n187));
  nor003aa1n03x5               g092(.a(new_n187), .b(new_n174), .c(new_n180), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n179), .b(new_n178), .c(new_n172), .o1(new_n189));
  oai013aa1n03x4               g094(.a(new_n189), .b(new_n169), .c(new_n174), .d(new_n180), .o1(new_n190));
  aoi012aa1n09x5               g095(.a(new_n190), .b(new_n155), .c(new_n188), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n192), .b(new_n186), .c(new_n191), .out0(\s[17] ));
  nor042aa1d18x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  inv040aa1n09x5               g099(.a(new_n194), .o1(new_n195));
  nona22aa1n02x4               g100(.a(new_n188), .b(new_n134), .c(new_n153), .out0(new_n196));
  aoai13aa1n09x5               g101(.a(new_n191), .b(new_n196), .c(new_n131), .d(new_n133), .o1(new_n197));
  nand22aa1n03x5               g102(.a(new_n197), .b(new_n192), .o1(new_n198));
  xnrc02aa1n02x5               g103(.a(\b[17] ), .b(\a[18] ), .out0(new_n199));
  xobna2aa1n03x5               g104(.a(new_n199), .b(new_n198), .c(new_n195), .out0(\s[18] ));
  inv000aa1d42x5               g105(.a(\a[17] ), .o1(new_n201));
  inv020aa1n04x5               g106(.a(\a[18] ), .o1(new_n202));
  xroi22aa1d06x4               g107(.a(new_n201), .b(\b[16] ), .c(new_n202), .d(\b[17] ), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  oaoi03aa1n12x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n195), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n204), .c(new_n186), .d(new_n191), .o1(new_n207));
  xorb03aa1n02x5               g112(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nand42aa1d28x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nor042aa1n04x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand42aa1n16x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanb02aa1n02x5               g118(.a(new_n212), .b(new_n213), .out0(new_n214));
  aoai13aa1n03x5               g119(.a(new_n214), .b(new_n210), .c(new_n207), .d(new_n211), .o1(new_n215));
  nand22aa1n03x5               g120(.a(new_n197), .b(new_n203), .o1(new_n216));
  nanb02aa1n02x5               g121(.a(new_n210), .b(new_n211), .out0(new_n217));
  norb03aa1n02x5               g122(.a(new_n213), .b(new_n210), .c(new_n212), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n217), .c(new_n216), .d(new_n206), .o1(new_n219));
  nanp02aa1n03x5               g124(.a(new_n215), .b(new_n219), .o1(\s[20] ));
  nano23aa1d15x5               g125(.a(new_n210), .b(new_n212), .c(new_n213), .d(new_n211), .out0(new_n221));
  nano22aa1n03x7               g126(.a(new_n199), .b(new_n221), .c(new_n192), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  nand02aa1d08x5               g128(.a(new_n221), .b(new_n205), .o1(new_n224));
  tech160nm_fioai012aa1n03p5x5 g129(.a(new_n213), .b(new_n212), .c(new_n210), .o1(new_n225));
  nand22aa1n03x5               g130(.a(new_n224), .b(new_n225), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n223), .c(new_n186), .d(new_n191), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand02aa1n08x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  nor042aa1n09x5               g137(.a(\b[21] ), .b(\a[22] ), .o1(new_n233));
  nand02aa1d28x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n230), .c(new_n228), .d(new_n232), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n232), .b(new_n226), .c(new_n197), .d(new_n222), .o1(new_n238));
  nona22aa1n03x5               g143(.a(new_n238), .b(new_n236), .c(new_n230), .out0(new_n239));
  nanp02aa1n03x5               g144(.a(new_n237), .b(new_n239), .o1(\s[22] ));
  nano23aa1d15x5               g145(.a(new_n230), .b(new_n233), .c(new_n234), .d(new_n231), .out0(new_n241));
  nanp03aa1n02x5               g146(.a(new_n203), .b(new_n221), .c(new_n241), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n234), .o1(new_n243));
  oab012aa1d18x5               g148(.a(new_n243), .b(new_n230), .c(new_n233), .out0(new_n244));
  aoi012aa1n03x5               g149(.a(new_n244), .b(new_n226), .c(new_n241), .o1(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n242), .c(new_n186), .d(new_n191), .o1(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1d32x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  nand02aa1n06x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  nor002aa1d32x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nand02aa1d28x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n248), .c(new_n246), .d(new_n250), .o1(new_n255));
  nanp02aa1n03x5               g160(.a(new_n246), .b(new_n250), .o1(new_n256));
  nona22aa1d36x5               g161(.a(new_n252), .b(new_n251), .c(new_n248), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  tech160nm_finand02aa1n03p5x5 g163(.a(new_n256), .b(new_n258), .o1(new_n259));
  nanp02aa1n03x5               g164(.a(new_n255), .b(new_n259), .o1(\s[24] ));
  nano23aa1d15x5               g165(.a(new_n248), .b(new_n251), .c(new_n252), .d(new_n249), .out0(new_n261));
  nand22aa1n12x5               g166(.a(new_n261), .b(new_n241), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(new_n222), .b(new_n263), .o1(new_n264));
  aoi022aa1d24x5               g169(.a(new_n261), .b(new_n244), .c(new_n252), .d(new_n257), .o1(new_n265));
  aoai13aa1n12x5               g170(.a(new_n265), .b(new_n262), .c(new_n224), .d(new_n225), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n264), .c(new_n186), .d(new_n191), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  inv000aa1d42x5               g174(.a(new_n221), .o1(new_n270));
  nona32aa1n03x5               g175(.a(new_n197), .b(new_n262), .c(new_n270), .d(new_n204), .out0(new_n271));
  xnrc02aa1n12x5               g176(.a(\b[24] ), .b(\a[25] ), .out0(new_n272));
  aoi012aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n267), .o1(new_n273));
  norp02aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n272), .o1(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n274), .c(new_n268), .d(new_n275), .o1(new_n277));
  oabi12aa1n02x5               g182(.a(new_n276), .b(\a[25] ), .c(\b[24] ), .out0(new_n278));
  oai012aa1n03x5               g183(.a(new_n277), .b(new_n273), .c(new_n278), .o1(\s[26] ));
  nor042aa1n02x5               g184(.a(new_n276), .b(new_n272), .o1(new_n280));
  nano32aa1n03x7               g185(.a(new_n262), .b(new_n203), .c(new_n280), .d(new_n221), .out0(new_n281));
  inv020aa1n03x5               g186(.a(new_n281), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(\b[25] ), .b(\a[26] ), .o1(new_n283));
  aoi022aa1n06x5               g188(.a(new_n266), .b(new_n280), .c(new_n283), .d(new_n278), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n282), .c(new_n186), .d(new_n191), .o1(new_n285));
  xorb03aa1n03x5               g190(.a(new_n285), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[27] ), .b(\b[26] ), .out0(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[27] ), .b(\a[28] ), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n287), .c(new_n285), .d(new_n288), .o1(new_n290));
  nanp02aa1n03x5               g195(.a(new_n266), .b(new_n280), .o1(new_n291));
  oai012aa1n02x5               g196(.a(new_n283), .b(new_n276), .c(new_n274), .o1(new_n292));
  nanp02aa1n06x5               g197(.a(new_n291), .b(new_n292), .o1(new_n293));
  aoai13aa1n02x7               g198(.a(new_n288), .b(new_n293), .c(new_n197), .d(new_n281), .o1(new_n294));
  nona22aa1n03x5               g199(.a(new_n294), .b(new_n289), .c(new_n287), .out0(new_n295));
  nanp02aa1n03x5               g200(.a(new_n290), .b(new_n295), .o1(\s[28] ));
  norb02aa1n02x5               g201(.a(new_n288), .b(new_n289), .out0(new_n297));
  aoai13aa1n02x7               g202(.a(new_n297), .b(new_n293), .c(new_n197), .d(new_n281), .o1(new_n298));
  tech160nm_fixorc02aa1n03p5x5 g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(\a[28] ), .o1(new_n301));
  inv000aa1d42x5               g206(.a(\b[27] ), .o1(new_n302));
  oao003aa1n02x5               g207(.a(new_n301), .b(new_n302), .c(new_n287), .carry(new_n303));
  nona22aa1n03x5               g208(.a(new_n298), .b(new_n300), .c(new_n303), .out0(new_n304));
  aoai13aa1n02x7               g209(.a(new_n300), .b(new_n303), .c(new_n285), .d(new_n297), .o1(new_n305));
  nanp02aa1n03x5               g210(.a(new_n305), .b(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g211(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g212(.a(new_n289), .b(new_n288), .c(new_n299), .out0(new_n308));
  inv000aa1n03x5               g213(.a(new_n303), .o1(new_n309));
  oaoi03aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .o1(new_n310));
  xnrc02aa1n02x5               g215(.a(\b[29] ), .b(\a[30] ), .out0(new_n311));
  aoai13aa1n02x7               g216(.a(new_n311), .b(new_n310), .c(new_n285), .d(new_n308), .o1(new_n312));
  aoai13aa1n02x7               g217(.a(new_n308), .b(new_n293), .c(new_n197), .d(new_n281), .o1(new_n313));
  nona22aa1n03x5               g218(.a(new_n313), .b(new_n310), .c(new_n311), .out0(new_n314));
  nanp02aa1n03x5               g219(.a(new_n312), .b(new_n314), .o1(\s[30] ));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  nano23aa1n02x4               g221(.a(new_n311), .b(new_n289), .c(new_n288), .d(new_n299), .out0(new_n317));
  and002aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .o(new_n318));
  oab012aa1n02x4               g223(.a(new_n318), .b(new_n310), .c(new_n311), .out0(new_n319));
  aoai13aa1n02x7               g224(.a(new_n316), .b(new_n319), .c(new_n285), .d(new_n317), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n317), .b(new_n293), .c(new_n197), .d(new_n281), .o1(new_n321));
  nona22aa1n03x5               g226(.a(new_n321), .b(new_n319), .c(new_n316), .out0(new_n322));
  nanp02aa1n03x5               g227(.a(new_n320), .b(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  xnrc02aa1n02x5               g229(.a(\b[3] ), .b(\a[4] ), .out0(new_n325));
  oaoi03aa1n02x5               g230(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n326));
  aob012aa1n02x5               g231(.a(new_n130), .b(new_n326), .c(new_n325), .out0(\s[4] ));
  inv000aa1d42x5               g232(.a(new_n107), .o1(new_n328));
  xobna2aa1n03x5               g233(.a(new_n104), .b(new_n130), .c(new_n328), .out0(\s[5] ));
  nanp03aa1n02x5               g234(.a(new_n130), .b(new_n104), .c(new_n328), .o1(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n105), .b(new_n330), .c(new_n119), .out0(\s[6] ));
  norb02aa1n02x5               g236(.a(new_n105), .b(new_n118), .out0(new_n332));
  aoi022aa1n02x5               g237(.a(new_n330), .b(new_n332), .c(\a[6] ), .d(\b[5] ), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nano22aa1n02x4               g239(.a(new_n101), .b(new_n333), .c(new_n102), .out0(new_n335));
  obai22aa1n02x7               g240(.a(new_n100), .b(new_n99), .c(new_n335), .d(new_n101), .out0(new_n336));
  oai012aa1n02x5               g241(.a(new_n336), .b(new_n335), .c(new_n132), .o1(\s[8] ));
  xnbna2aa1n03x5               g242(.a(new_n123), .b(new_n131), .c(new_n133), .out0(\s[9] ));
endmodule


