// Benchmark "adder" written by ABC on Thu Jul 18 08:25:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n300, new_n303, new_n305, new_n306,
    new_n308, new_n309, new_n310;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  tech160nm_finand02aa1n03p5x5 g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n06x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1n12x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  norp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n02x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  aoi012aa1n02x7               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor022aa1n02x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n03x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  aoi012aa1n02x5               g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1n06x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  nor022aa1n08x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n03x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .out0(new_n118));
  xnrc02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .out0(new_n119));
  nor043aa1n03x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  tech160nm_fioai012aa1n03p5x5 g025(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n121));
  orn002aa1n03x5               g026(.a(\a[5] ), .b(\b[4] ), .o(new_n122));
  tech160nm_fioaoi03aa1n03p5x5 g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  oaib12aa1n18x5               g028(.a(new_n121), .b(new_n117), .c(new_n123), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n112), .d(new_n120), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n99), .b(new_n126), .c(new_n101), .out0(\s[10] ));
  nanp02aa1n03x5               g032(.a(new_n126), .b(new_n101), .o1(new_n128));
  nor002aa1n06x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nand42aa1n06x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  aoai13aa1n06x5               g036(.a(new_n131), .b(new_n97), .c(new_n128), .d(new_n99), .o1(new_n132));
  aoi112aa1n02x5               g037(.a(new_n131), .b(new_n97), .c(new_n128), .d(new_n99), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n132), .b(new_n133), .out0(\s[11] ));
  orn002aa1n02x5               g039(.a(\a[11] ), .b(\b[10] ), .o(new_n135));
  nor042aa1n06x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanp02aa1n09x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aobi12aa1n06x5               g043(.a(new_n138), .b(new_n132), .c(new_n135), .out0(new_n139));
  nona22aa1n02x4               g044(.a(new_n132), .b(new_n138), .c(new_n129), .out0(new_n140));
  norb02aa1n03x4               g045(.a(new_n140), .b(new_n139), .out0(\s[12] ));
  nanp02aa1n02x5               g046(.a(new_n112), .b(new_n120), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n124), .o1(new_n143));
  nano23aa1n03x5               g048(.a(new_n129), .b(new_n136), .c(new_n137), .d(new_n130), .out0(new_n144));
  nand03aa1n02x5               g049(.a(new_n144), .b(new_n99), .c(new_n125), .o1(new_n145));
  nona23aa1n09x5               g050(.a(new_n137), .b(new_n130), .c(new_n129), .d(new_n136), .out0(new_n146));
  tech160nm_fioai012aa1n03p5x5 g051(.a(new_n137), .b(new_n136), .c(new_n129), .o1(new_n147));
  tech160nm_fioai012aa1n05x5   g052(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n148));
  oai012aa1n12x5               g053(.a(new_n147), .b(new_n146), .c(new_n148), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n145), .c(new_n143), .d(new_n142), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n09x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand42aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nano23aa1n03x7               g063(.a(new_n153), .b(new_n157), .c(new_n158), .d(new_n154), .out0(new_n159));
  oai012aa1n12x5               g064(.a(new_n158), .b(new_n157), .c(new_n153), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  xorc02aa1n02x5               g066(.a(\a[15] ), .b(\b[14] ), .out0(new_n162));
  aoai13aa1n04x5               g067(.a(new_n162), .b(new_n161), .c(new_n151), .d(new_n159), .o1(new_n163));
  aoi112aa1n02x5               g068(.a(new_n162), .b(new_n161), .c(new_n151), .d(new_n159), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(\s[15] ));
  xnrc02aa1n12x5               g070(.a(\b[15] ), .b(\a[16] ), .out0(new_n166));
  oaoi13aa1n03x5               g071(.a(new_n166), .b(new_n163), .c(\a[15] ), .d(\b[14] ), .o1(new_n167));
  oai112aa1n03x5               g072(.a(new_n163), .b(new_n166), .c(\b[14] ), .d(\a[15] ), .o1(new_n168));
  norb02aa1n02x7               g073(.a(new_n168), .b(new_n167), .out0(\s[16] ));
  inv000aa1d42x5               g074(.a(new_n166), .o1(new_n170));
  nano32aa1n03x7               g075(.a(new_n145), .b(new_n170), .c(new_n159), .d(new_n162), .out0(new_n171));
  aoai13aa1n12x5               g076(.a(new_n171), .b(new_n124), .c(new_n112), .d(new_n120), .o1(new_n172));
  nona23aa1n02x4               g077(.a(new_n158), .b(new_n154), .c(new_n153), .d(new_n157), .out0(new_n173));
  xnrc02aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .out0(new_n174));
  nor043aa1n02x5               g079(.a(new_n173), .b(new_n174), .c(new_n166), .o1(new_n175));
  aoi112aa1n02x5               g080(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n176));
  orn002aa1n02x5               g081(.a(\a[16] ), .b(\b[15] ), .o(new_n177));
  oai013aa1n03x4               g082(.a(new_n177), .b(new_n174), .c(new_n166), .d(new_n160), .o1(new_n178));
  aoi112aa1n09x5               g083(.a(new_n178), .b(new_n176), .c(new_n149), .d(new_n175), .o1(new_n179));
  nand02aa1d08x5               g084(.a(new_n172), .b(new_n179), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g086(.a(\a[18] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  oaoi03aa1n03x5               g089(.a(new_n183), .b(new_n184), .c(new_n180), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n182), .out0(\s[18] ));
  xroi22aa1d04x5               g091(.a(new_n183), .b(\b[16] ), .c(new_n182), .d(\b[17] ), .out0(new_n187));
  nanp02aa1n02x5               g092(.a(new_n184), .b(new_n183), .o1(new_n188));
  oaoi03aa1n02x5               g093(.a(\a[18] ), .b(\b[17] ), .c(new_n188), .o1(new_n189));
  tech160nm_fiaoi012aa1n05x5   g094(.a(new_n189), .b(new_n180), .c(new_n187), .o1(new_n190));
  nor042aa1n09x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  nand42aa1n03x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n190), .b(new_n193), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g100(.a(new_n191), .b(new_n193), .out0(new_n196));
  nor002aa1n04x5               g101(.a(\b[19] ), .b(\a[20] ), .o1(new_n197));
  nand22aa1n03x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nanb02aa1n02x5               g103(.a(new_n197), .b(new_n198), .out0(new_n199));
  oaoi13aa1n02x7               g104(.a(new_n199), .b(new_n192), .c(new_n190), .d(new_n196), .o1(new_n200));
  nor042aa1n02x5               g105(.a(new_n190), .b(new_n196), .o1(new_n201));
  nano22aa1n03x7               g106(.a(new_n201), .b(new_n192), .c(new_n199), .out0(new_n202));
  norp02aa1n03x5               g107(.a(new_n200), .b(new_n202), .o1(\s[20] ));
  nano23aa1n09x5               g108(.a(new_n191), .b(new_n197), .c(new_n198), .d(new_n193), .out0(new_n204));
  nanp02aa1n02x5               g109(.a(new_n187), .b(new_n204), .o1(new_n205));
  oai022aa1n02x5               g110(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n206));
  oaib12aa1n02x5               g111(.a(new_n206), .b(new_n182), .c(\b[17] ), .out0(new_n207));
  nona23aa1n09x5               g112(.a(new_n198), .b(new_n193), .c(new_n191), .d(new_n197), .out0(new_n208));
  tech160nm_fiaoi012aa1n04x5   g113(.a(new_n197), .b(new_n191), .c(new_n198), .o1(new_n209));
  oai012aa1n12x5               g114(.a(new_n209), .b(new_n208), .c(new_n207), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n205), .c(new_n172), .d(new_n179), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g118(.a(\b[20] ), .b(\a[21] ), .o1(new_n214));
  xorc02aa1n02x5               g119(.a(\a[21] ), .b(\b[20] ), .out0(new_n215));
  xorc02aa1n02x5               g120(.a(\a[22] ), .b(\b[21] ), .out0(new_n216));
  aoai13aa1n02x7               g121(.a(new_n216), .b(new_n214), .c(new_n212), .d(new_n215), .o1(new_n217));
  aoi112aa1n02x5               g122(.a(new_n214), .b(new_n216), .c(new_n212), .d(new_n215), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(\s[22] ));
  inv000aa1d42x5               g124(.a(\a[21] ), .o1(new_n220));
  inv000aa1d42x5               g125(.a(\a[22] ), .o1(new_n221));
  xroi22aa1d04x5               g126(.a(new_n220), .b(\b[20] ), .c(new_n221), .d(\b[21] ), .out0(new_n222));
  nanp03aa1n02x5               g127(.a(new_n222), .b(new_n187), .c(new_n204), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[21] ), .o1(new_n224));
  oaoi03aa1n12x5               g129(.a(new_n221), .b(new_n224), .c(new_n214), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoi012aa1n02x5               g131(.a(new_n226), .b(new_n210), .c(new_n222), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n223), .c(new_n172), .d(new_n179), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g134(.a(\b[22] ), .b(\a[23] ), .o1(new_n230));
  tech160nm_fixorc02aa1n05x5   g135(.a(\a[23] ), .b(\b[22] ), .out0(new_n231));
  xorc02aa1n03x5               g136(.a(\a[24] ), .b(\b[23] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n233));
  aoi112aa1n02x5               g138(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n233), .b(new_n234), .out0(\s[24] ));
  and002aa1n06x5               g140(.a(new_n232), .b(new_n231), .o(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nano32aa1n02x4               g142(.a(new_n237), .b(new_n222), .c(new_n187), .d(new_n204), .out0(new_n238));
  inv020aa1n02x5               g143(.a(new_n209), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n222), .b(new_n239), .c(new_n204), .d(new_n189), .o1(new_n240));
  norp02aa1n02x5               g145(.a(\b[23] ), .b(\a[24] ), .o1(new_n241));
  nanp02aa1n02x5               g146(.a(\b[23] ), .b(\a[24] ), .o1(new_n242));
  aoi012aa1n02x5               g147(.a(new_n241), .b(new_n230), .c(new_n242), .o1(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n237), .c(new_n240), .d(new_n225), .o1(new_n244));
  tech160nm_fixorc02aa1n05x5   g149(.a(\a[25] ), .b(\b[24] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n244), .c(new_n180), .d(new_n238), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n245), .b(new_n244), .c(new_n180), .d(new_n238), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  tech160nm_fixorc02aa1n05x5   g155(.a(\a[26] ), .b(\b[25] ), .out0(new_n251));
  aobi12aa1n06x5               g156(.a(new_n251), .b(new_n246), .c(new_n250), .out0(new_n252));
  nona22aa1n02x5               g157(.a(new_n246), .b(new_n251), .c(new_n249), .out0(new_n253));
  norb02aa1n03x4               g158(.a(new_n253), .b(new_n252), .out0(\s[26] ));
  and002aa1n06x5               g159(.a(new_n251), .b(new_n245), .o(new_n255));
  nano22aa1n03x7               g160(.a(new_n223), .b(new_n236), .c(new_n255), .out0(new_n256));
  nand22aa1n09x5               g161(.a(new_n180), .b(new_n256), .o1(new_n257));
  oao003aa1n02x5               g162(.a(\a[26] ), .b(\b[25] ), .c(new_n250), .carry(new_n258));
  aobi12aa1n09x5               g163(.a(new_n258), .b(new_n244), .c(new_n255), .out0(new_n259));
  xorc02aa1n02x5               g164(.a(\a[27] ), .b(\b[26] ), .out0(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n259), .c(new_n257), .out0(\s[27] ));
  norp02aa1n02x5               g166(.a(\b[26] ), .b(\a[27] ), .o1(new_n262));
  inv040aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  aobi12aa1n06x5               g168(.a(new_n256), .b(new_n172), .c(new_n179), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n236), .b(new_n226), .c(new_n210), .d(new_n222), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n255), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n258), .b(new_n266), .c(new_n265), .d(new_n243), .o1(new_n267));
  oaih12aa1n02x5               g172(.a(new_n260), .b(new_n267), .c(new_n264), .o1(new_n268));
  xnrc02aa1n02x5               g173(.a(\b[27] ), .b(\a[28] ), .out0(new_n269));
  aoi012aa1n03x5               g174(.a(new_n269), .b(new_n268), .c(new_n263), .o1(new_n270));
  aobi12aa1n06x5               g175(.a(new_n260), .b(new_n259), .c(new_n257), .out0(new_n271));
  nano22aa1n03x5               g176(.a(new_n271), .b(new_n263), .c(new_n269), .out0(new_n272));
  nor002aa1n02x5               g177(.a(new_n270), .b(new_n272), .o1(\s[28] ));
  norb02aa1n02x5               g178(.a(new_n260), .b(new_n269), .out0(new_n274));
  oaih12aa1n02x5               g179(.a(new_n274), .b(new_n267), .c(new_n264), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[28] ), .b(\b[27] ), .c(new_n263), .carry(new_n276));
  xnrc02aa1n02x5               g181(.a(\b[28] ), .b(\a[29] ), .out0(new_n277));
  aoi012aa1n02x5               g182(.a(new_n277), .b(new_n275), .c(new_n276), .o1(new_n278));
  aobi12aa1n06x5               g183(.a(new_n274), .b(new_n259), .c(new_n257), .out0(new_n279));
  nano22aa1n03x7               g184(.a(new_n279), .b(new_n276), .c(new_n277), .out0(new_n280));
  norp02aa1n03x5               g185(.a(new_n278), .b(new_n280), .o1(\s[29] ));
  xorb03aa1n02x5               g186(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g187(.a(new_n260), .b(new_n277), .c(new_n269), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n283), .b(new_n267), .c(new_n264), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[29] ), .b(\b[28] ), .c(new_n276), .carry(new_n285));
  xnrc02aa1n02x5               g190(.a(\b[29] ), .b(\a[30] ), .out0(new_n286));
  aoi012aa1n02x5               g191(.a(new_n286), .b(new_n284), .c(new_n285), .o1(new_n287));
  aobi12aa1n06x5               g192(.a(new_n283), .b(new_n259), .c(new_n257), .out0(new_n288));
  nano22aa1n03x7               g193(.a(new_n288), .b(new_n285), .c(new_n286), .out0(new_n289));
  norp02aa1n03x5               g194(.a(new_n287), .b(new_n289), .o1(\s[30] ));
  norb02aa1n02x5               g195(.a(new_n283), .b(new_n286), .out0(new_n291));
  aobi12aa1n06x5               g196(.a(new_n291), .b(new_n259), .c(new_n257), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[30] ), .b(\b[29] ), .c(new_n285), .carry(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[30] ), .b(\a[31] ), .out0(new_n294));
  nano22aa1n03x7               g199(.a(new_n292), .b(new_n293), .c(new_n294), .out0(new_n295));
  oaih12aa1n02x5               g200(.a(new_n291), .b(new_n267), .c(new_n264), .o1(new_n296));
  aoi012aa1n03x5               g201(.a(new_n294), .b(new_n296), .c(new_n293), .o1(new_n297));
  nor002aa1n02x5               g202(.a(new_n297), .b(new_n295), .o1(\s[31] ));
  xnrb03aa1n02x5               g203(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g204(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n300));
  xorb03aa1n02x5               g205(.a(new_n300), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g206(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaib12aa1n02x5               g207(.a(new_n122), .b(new_n119), .c(new_n112), .out0(new_n303));
  xorb03aa1n02x5               g208(.a(new_n303), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g209(.a(new_n118), .b(new_n303), .out0(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(\b[5] ), .c(\a[6] ), .o1(new_n306));
  xorb03aa1n02x5               g211(.a(new_n306), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  norb02aa1n02x5               g212(.a(new_n114), .b(new_n113), .out0(new_n308));
  aoai13aa1n02x5               g213(.a(new_n308), .b(new_n115), .c(new_n306), .d(new_n116), .o1(new_n309));
  aoi112aa1n02x5               g214(.a(new_n308), .b(new_n115), .c(new_n306), .d(new_n116), .o1(new_n310));
  norb02aa1n02x5               g215(.a(new_n309), .b(new_n310), .out0(\s[8] ));
  xnbna2aa1n03x5               g216(.a(new_n125), .b(new_n143), .c(new_n142), .out0(\s[9] ));
endmodule


