// Benchmark "adder" written by ABC on Wed Jul 17 17:52:18 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n321, new_n322, new_n324,
    new_n325, new_n327, new_n328, new_n330, new_n331, new_n333, new_n334,
    new_n335, new_n337, new_n338, new_n339, new_n340, new_n342, new_n343,
    new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand22aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  oab012aa1d18x5               g004(.a(new_n99), .b(\a[2] ), .c(\b[1] ), .out0(new_n100));
  nand42aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanb03aa1n12x5               g008(.a(new_n102), .b(new_n103), .c(new_n101), .out0(new_n104));
  oab012aa1n06x5               g009(.a(new_n102), .b(\a[4] ), .c(\b[3] ), .out0(new_n105));
  oai012aa1n18x5               g010(.a(new_n105), .b(new_n104), .c(new_n100), .o1(new_n106));
  nanp02aa1n09x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nand02aa1d10x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  inv040aa1d32x5               g013(.a(\a[8] ), .o1(new_n109));
  inv020aa1d32x5               g014(.a(\b[7] ), .o1(new_n110));
  nand02aa1n08x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nand03aa1n02x5               g016(.a(new_n111), .b(new_n107), .c(new_n108), .o1(new_n112));
  oaih22aa1n04x5               g017(.a(\a[6] ), .b(\b[5] ), .c(\b[6] ), .d(\a[7] ), .o1(new_n113));
  aoi022aa1d24x5               g018(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  oai112aa1n06x5               g020(.a(new_n114), .b(new_n115), .c(\b[4] ), .d(\a[5] ), .o1(new_n116));
  nor043aa1n06x5               g021(.a(new_n116), .b(new_n112), .c(new_n113), .o1(new_n117));
  orn002aa1n24x5               g022(.a(\a[7] ), .b(\b[6] ), .o(new_n118));
  nor002aa1d32x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor042aa1n06x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  oai012aa1d24x5               g025(.a(new_n108), .b(new_n120), .c(new_n119), .o1(new_n121));
  aob012aa1n03x5               g026(.a(new_n107), .b(\b[6] ), .c(\a[7] ), .out0(new_n122));
  aoai13aa1n12x5               g027(.a(new_n111), .b(new_n122), .c(new_n121), .d(new_n118), .o1(new_n123));
  nanp02aa1n24x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  norb02aa1n06x4               g029(.a(new_n124), .b(new_n97), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n126));
  nor042aa1n04x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand22aa1n09x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n06x4               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nona23aa1n02x4               g034(.a(new_n126), .b(new_n128), .c(new_n127), .d(new_n97), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .d(new_n126), .o1(\s[10] ));
  nano23aa1n02x4               g036(.a(new_n97), .b(new_n127), .c(new_n128), .d(new_n124), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n133));
  aoi012aa1d18x5               g038(.a(new_n127), .b(new_n97), .c(new_n128), .o1(new_n134));
  nor002aa1d24x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanp02aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  aob012aa1n02x5               g044(.a(new_n138), .b(new_n133), .c(new_n134), .out0(new_n140));
  nor002aa1d32x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand02aa1n08x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  oaib12aa1n02x5               g048(.a(new_n143), .b(new_n135), .c(new_n140), .out0(new_n144));
  nona23aa1n02x4               g049(.a(new_n140), .b(new_n142), .c(new_n141), .d(new_n135), .out0(new_n145));
  nanp02aa1n02x5               g050(.a(new_n144), .b(new_n145), .o1(\s[12] ));
  nona23aa1d18x5               g051(.a(new_n142), .b(new_n136), .c(new_n135), .d(new_n141), .out0(new_n147));
  nano22aa1n03x7               g052(.a(new_n147), .b(new_n125), .c(new_n129), .out0(new_n148));
  aoai13aa1n06x5               g053(.a(new_n148), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n149));
  oaih12aa1n12x5               g054(.a(new_n142), .b(new_n141), .c(new_n135), .o1(new_n150));
  oai012aa1d24x5               g055(.a(new_n150), .b(new_n147), .c(new_n134), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand22aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  aob012aa1n02x5               g060(.a(new_n155), .b(new_n149), .c(new_n152), .out0(new_n156));
  oaib12aa1n02x5               g061(.a(new_n150), .b(new_n153), .c(new_n154), .out0(new_n157));
  oab012aa1n02x4               g062(.a(new_n157), .b(new_n147), .c(new_n134), .out0(new_n158));
  aobi12aa1n02x5               g063(.a(new_n156), .b(new_n158), .c(new_n149), .out0(\s[13] ));
  inv000aa1d42x5               g064(.a(new_n153), .o1(new_n160));
  nor022aa1n12x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand22aa1n12x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  nona23aa1n02x4               g068(.a(new_n156), .b(new_n162), .c(new_n161), .d(new_n153), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n163), .c(new_n160), .d(new_n156), .o1(\s[14] ));
  nona23aa1d16x5               g070(.a(new_n162), .b(new_n154), .c(new_n153), .d(new_n161), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aob012aa1n06x5               g072(.a(new_n167), .b(new_n149), .c(new_n152), .out0(new_n168));
  aoi012aa1n02x5               g073(.a(new_n161), .b(new_n153), .c(new_n162), .o1(new_n169));
  xnrc02aa1n12x5               g074(.a(\b[14] ), .b(\a[15] ), .out0(new_n170));
  xobna2aa1n03x5               g075(.a(new_n170), .b(new_n168), .c(new_n169), .out0(\s[15] ));
  nor042aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n06x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  inv000aa1d42x5               g079(.a(\a[15] ), .o1(new_n175));
  inv000aa1d42x5               g080(.a(\b[14] ), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(new_n176), .b(new_n175), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n170), .c(new_n168), .d(new_n169), .o1(new_n178));
  nano22aa1n02x4               g083(.a(new_n172), .b(new_n177), .c(new_n173), .out0(new_n179));
  aoai13aa1n02x5               g084(.a(new_n179), .b(new_n170), .c(new_n168), .d(new_n169), .o1(new_n180));
  aob012aa1n02x5               g085(.a(new_n180), .b(new_n178), .c(new_n174), .out0(\s[16] ));
  xnrc02aa1n02x5               g086(.a(\b[16] ), .b(\a[17] ), .out0(new_n182));
  aoi012aa1d18x5               g087(.a(new_n123), .b(new_n117), .c(new_n106), .o1(new_n183));
  nor043aa1d12x5               g088(.a(new_n166), .b(new_n170), .c(new_n174), .o1(new_n184));
  nand22aa1n09x5               g089(.a(new_n184), .b(new_n148), .o1(new_n185));
  oai022aa1n03x5               g090(.a(\a[14] ), .b(\b[13] ), .c(\b[14] ), .d(\a[15] ), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n187));
  aoai13aa1n02x7               g092(.a(new_n187), .b(new_n186), .c(new_n153), .d(new_n162), .o1(new_n188));
  tech160nm_fioai012aa1n04x5   g093(.a(new_n188), .b(\b[15] ), .c(\a[16] ), .o1(new_n189));
  aoi012aa1n12x5               g094(.a(new_n189), .b(new_n151), .c(new_n184), .o1(new_n190));
  oai012aa1d24x5               g095(.a(new_n190), .b(new_n183), .c(new_n185), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(new_n151), .b(new_n184), .o1(new_n192));
  nor042aa1n06x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  inv000aa1n06x5               g098(.a(new_n193), .o1(new_n194));
  and002aa1n02x5               g099(.a(\b[16] ), .b(\a[17] ), .o(new_n195));
  nona22aa1n02x4               g100(.a(new_n194), .b(new_n195), .c(new_n172), .out0(new_n196));
  norb02aa1n02x5               g101(.a(new_n188), .b(new_n196), .out0(new_n197));
  oai112aa1n02x5               g102(.a(new_n192), .b(new_n197), .c(new_n183), .d(new_n185), .o1(new_n198));
  aob012aa1n02x5               g103(.a(new_n198), .b(new_n191), .c(new_n182), .out0(\s[17] ));
  inv000aa1d42x5               g104(.a(\b[16] ), .o1(new_n200));
  oaib12aa1n02x5               g105(.a(new_n191), .b(new_n200), .c(\a[17] ), .out0(new_n201));
  xorc02aa1n12x5               g106(.a(\a[18] ), .b(\b[17] ), .out0(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n201), .c(new_n194), .out0(\s[18] ));
  norb02aa1n02x5               g108(.a(new_n202), .b(new_n182), .out0(new_n204));
  oaoi03aa1n09x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n194), .o1(new_n205));
  xorc02aa1n12x5               g110(.a(\a[19] ), .b(\b[18] ), .out0(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n205), .c(new_n191), .d(new_n204), .o1(new_n207));
  aoi112aa1n02x5               g112(.a(new_n206), .b(new_n205), .c(new_n191), .d(new_n204), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n207), .b(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  orn002aa1n02x5               g115(.a(\a[19] ), .b(\b[18] ), .o(new_n211));
  xorc02aa1n12x5               g116(.a(\a[20] ), .b(\b[19] ), .out0(new_n212));
  oai022aa1n02x7               g117(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n213));
  aoi012aa1n02x5               g118(.a(new_n213), .b(\a[20] ), .c(\b[19] ), .o1(new_n214));
  nanp02aa1n02x5               g119(.a(new_n207), .b(new_n214), .o1(new_n215));
  aoai13aa1n02x5               g120(.a(new_n215), .b(new_n212), .c(new_n207), .d(new_n211), .o1(\s[20] ));
  nano32aa1n03x7               g121(.a(new_n182), .b(new_n212), .c(new_n202), .d(new_n206), .out0(new_n217));
  nanp03aa1d12x5               g122(.a(new_n205), .b(new_n206), .c(new_n212), .o1(new_n218));
  aob012aa1n06x5               g123(.a(new_n213), .b(\b[19] ), .c(\a[20] ), .out0(new_n219));
  nanp02aa1n02x5               g124(.a(new_n218), .b(new_n219), .o1(new_n220));
  xorc02aa1n12x5               g125(.a(\a[21] ), .b(\b[20] ), .out0(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n220), .c(new_n191), .d(new_n217), .o1(new_n222));
  nano22aa1n02x4               g127(.a(new_n221), .b(new_n218), .c(new_n219), .out0(new_n223));
  aobi12aa1n02x5               g128(.a(new_n223), .b(new_n191), .c(new_n217), .out0(new_n224));
  norb02aa1n02x5               g129(.a(new_n222), .b(new_n224), .out0(\s[21] ));
  norp02aa1n02x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  inv000aa1n02x5               g131(.a(new_n226), .o1(new_n227));
  nor002aa1n03x5               g132(.a(\b[21] ), .b(\a[22] ), .o1(new_n228));
  and002aa1n12x5               g133(.a(\b[21] ), .b(\a[22] ), .o(new_n229));
  nor042aa1n04x5               g134(.a(new_n229), .b(new_n228), .o1(new_n230));
  norp03aa1n02x5               g135(.a(new_n229), .b(new_n228), .c(new_n226), .o1(new_n231));
  nand42aa1n03x5               g136(.a(new_n222), .b(new_n231), .o1(new_n232));
  aoai13aa1n02x5               g137(.a(new_n232), .b(new_n230), .c(new_n222), .d(new_n227), .o1(\s[22] ));
  nand02aa1d06x5               g138(.a(new_n221), .b(new_n230), .o1(new_n234));
  nano32aa1n02x4               g139(.a(new_n234), .b(new_n204), .c(new_n206), .d(new_n212), .out0(new_n235));
  oab012aa1n06x5               g140(.a(new_n228), .b(new_n227), .c(new_n229), .out0(new_n236));
  aoai13aa1n12x5               g141(.a(new_n236), .b(new_n234), .c(new_n218), .d(new_n219), .o1(new_n237));
  tech160nm_fixorc02aa1n03p5x5 g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n237), .c(new_n191), .d(new_n235), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n236), .b(new_n238), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n234), .c(new_n218), .d(new_n219), .o1(new_n241));
  aoi012aa1n02x5               g146(.a(new_n241), .b(new_n191), .c(new_n235), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n239), .b(new_n242), .out0(\s[23] ));
  nor042aa1n03x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  tech160nm_fixorc02aa1n02p5x5 g150(.a(\a[24] ), .b(\b[23] ), .out0(new_n246));
  and002aa1n02x5               g151(.a(\b[23] ), .b(\a[24] ), .o(new_n247));
  oai022aa1n02x5               g152(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n248));
  nona22aa1n06x5               g153(.a(new_n239), .b(new_n247), .c(new_n248), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n246), .c(new_n245), .d(new_n239), .o1(\s[24] ));
  nano22aa1n03x7               g155(.a(new_n234), .b(new_n238), .c(new_n246), .out0(new_n251));
  and002aa1n02x5               g156(.a(new_n217), .b(new_n251), .o(new_n252));
  and002aa1n02x5               g157(.a(new_n191), .b(new_n252), .o(new_n253));
  and002aa1n02x5               g158(.a(new_n246), .b(new_n238), .o(new_n254));
  nanp02aa1n02x5               g159(.a(new_n237), .b(new_n254), .o1(new_n255));
  oaib12aa1n02x5               g160(.a(new_n255), .b(new_n247), .c(new_n248), .out0(new_n256));
  tech160nm_fixorc02aa1n05x5   g161(.a(\a[25] ), .b(\b[24] ), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n256), .c(new_n191), .d(new_n252), .o1(new_n258));
  oaoi03aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n245), .o1(new_n259));
  nona22aa1n02x4               g164(.a(new_n255), .b(new_n259), .c(new_n257), .out0(new_n260));
  oa0012aa1n02x5               g165(.a(new_n258), .b(new_n260), .c(new_n253), .o(\s[25] ));
  norp02aa1n02x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[26] ), .b(\b[25] ), .out0(new_n264));
  and002aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .o(new_n265));
  oai022aa1n02x5               g170(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n266));
  nona22aa1n02x5               g171(.a(new_n258), .b(new_n265), .c(new_n266), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n264), .c(new_n263), .d(new_n258), .o1(\s[26] ));
  and002aa1n02x5               g173(.a(new_n264), .b(new_n257), .o(new_n269));
  aoai13aa1n12x5               g174(.a(new_n269), .b(new_n259), .c(new_n237), .d(new_n254), .o1(new_n270));
  nor042aa1d18x5               g175(.a(\b[26] ), .b(\a[27] ), .o1(new_n271));
  and002aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o(new_n272));
  norp02aa1n02x5               g177(.a(new_n272), .b(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n265), .o1(new_n274));
  and003aa1n06x5               g179(.a(new_n217), .b(new_n269), .c(new_n251), .o(new_n275));
  aoi122aa1n02x5               g180(.a(new_n273), .b(new_n274), .c(new_n266), .d(new_n191), .e(new_n275), .o1(new_n276));
  nand02aa1d04x5               g181(.a(new_n191), .b(new_n275), .o1(new_n277));
  aob012aa1n02x5               g182(.a(new_n266), .b(\b[25] ), .c(\a[26] ), .out0(new_n278));
  nanp03aa1n06x5               g183(.a(new_n277), .b(new_n270), .c(new_n278), .o1(new_n279));
  aoi022aa1n02x5               g184(.a(new_n276), .b(new_n270), .c(new_n279), .d(new_n273), .o1(\s[27] ));
  inv000aa1d42x5               g185(.a(\b[26] ), .o1(new_n281));
  oaib12aa1n03x5               g186(.a(new_n279), .b(new_n281), .c(\a[27] ), .out0(new_n282));
  inv040aa1n08x5               g187(.a(new_n271), .o1(new_n283));
  aoi022aa1n12x5               g188(.a(new_n191), .b(new_n275), .c(new_n274), .d(new_n266), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n283), .b(new_n272), .c(new_n284), .d(new_n270), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .out0(new_n286));
  norp02aa1n02x5               g191(.a(new_n286), .b(new_n271), .o1(new_n287));
  aoi022aa1n03x5               g192(.a(new_n285), .b(new_n286), .c(new_n282), .d(new_n287), .o1(\s[28] ));
  inv000aa1d42x5               g193(.a(\a[28] ), .o1(new_n289));
  xroi22aa1d04x5               g194(.a(\a[27] ), .b(new_n281), .c(new_n289), .d(\b[27] ), .out0(new_n290));
  nanp02aa1n03x5               g195(.a(new_n279), .b(new_n290), .o1(new_n291));
  inv000aa1n03x5               g196(.a(new_n290), .o1(new_n292));
  oao003aa1n03x5               g197(.a(\a[28] ), .b(\b[27] ), .c(new_n283), .carry(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n292), .c(new_n284), .d(new_n270), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[29] ), .b(\b[28] ), .out0(new_n295));
  norb02aa1n02x5               g200(.a(new_n293), .b(new_n295), .out0(new_n296));
  aoi022aa1n03x5               g201(.a(new_n294), .b(new_n295), .c(new_n291), .d(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g202(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g203(.a(new_n286), .b(new_n295), .c(new_n273), .o(new_n299));
  nanp02aa1n03x5               g204(.a(new_n279), .b(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n299), .o1(new_n301));
  tech160nm_fioaoi03aa1n03p5x5 g206(.a(\a[29] ), .b(\b[28] ), .c(new_n293), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n301), .c(new_n284), .d(new_n270), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .out0(new_n305));
  and002aa1n02x5               g210(.a(\b[28] ), .b(\a[29] ), .o(new_n306));
  oabi12aa1n02x5               g211(.a(new_n305), .b(\a[29] ), .c(\b[28] ), .out0(new_n307));
  oab012aa1n02x4               g212(.a(new_n307), .b(new_n293), .c(new_n306), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n304), .b(new_n305), .c(new_n300), .d(new_n308), .o1(\s[30] ));
  nano22aa1n02x4               g214(.a(new_n292), .b(new_n295), .c(new_n305), .out0(new_n310));
  nanp02aa1n03x5               g215(.a(new_n279), .b(new_n310), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[31] ), .b(\b[30] ), .out0(new_n312));
  inv000aa1d42x5               g217(.a(\a[30] ), .o1(new_n313));
  inv000aa1d42x5               g218(.a(\b[29] ), .o1(new_n314));
  oabi12aa1n02x5               g219(.a(new_n312), .b(\a[30] ), .c(\b[29] ), .out0(new_n315));
  oaoi13aa1n04x5               g220(.a(new_n315), .b(new_n302), .c(new_n313), .d(new_n314), .o1(new_n316));
  inv000aa1n02x5               g221(.a(new_n310), .o1(new_n317));
  oaoi03aa1n03x5               g222(.a(new_n313), .b(new_n314), .c(new_n302), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n284), .d(new_n270), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n319), .b(new_n312), .c(new_n311), .d(new_n316), .o1(\s[31] ));
  inv000aa1d42x5               g225(.a(new_n100), .o1(new_n321));
  nanb02aa1n02x5               g226(.a(new_n102), .b(new_n103), .out0(new_n322));
  xnbna2aa1n03x5               g227(.a(new_n322), .b(new_n321), .c(new_n101), .out0(\s[3] ));
  xorc02aa1n02x5               g228(.a(\a[4] ), .b(\b[3] ), .out0(new_n324));
  aoi113aa1n02x5               g229(.a(new_n324), .b(new_n102), .c(new_n321), .d(new_n103), .e(new_n101), .o1(new_n325));
  aoi012aa1n02x5               g230(.a(new_n325), .b(new_n106), .c(new_n324), .o1(\s[4] ));
  nanp02aa1n02x5               g231(.a(\b[4] ), .b(\a[5] ), .o1(new_n327));
  norb02aa1n02x5               g232(.a(new_n327), .b(new_n120), .out0(new_n328));
  xobna2aa1n03x5               g233(.a(new_n328), .b(new_n106), .c(new_n115), .out0(\s[5] ));
  aob012aa1n02x5               g234(.a(new_n328), .b(new_n106), .c(new_n115), .out0(new_n330));
  norb02aa1n02x5               g235(.a(new_n108), .b(new_n119), .out0(new_n331));
  xobna2aa1n03x5               g236(.a(new_n331), .b(new_n330), .c(new_n327), .out0(\s[6] ));
  inv000aa1d42x5               g237(.a(new_n119), .o1(new_n333));
  nanp03aa1n02x5               g238(.a(new_n330), .b(new_n327), .c(new_n331), .o1(new_n334));
  xorc02aa1n02x5               g239(.a(\a[7] ), .b(\b[6] ), .out0(new_n335));
  xnbna2aa1n03x5               g240(.a(new_n335), .b(new_n334), .c(new_n333), .out0(\s[7] ));
  aob012aa1n02x5               g241(.a(new_n335), .b(new_n334), .c(new_n333), .out0(new_n337));
  xorc02aa1n02x5               g242(.a(\a[8] ), .b(\b[7] ), .out0(new_n338));
  and003aa1n02x5               g243(.a(new_n118), .b(new_n111), .c(new_n107), .o(new_n339));
  nanp02aa1n02x5               g244(.a(new_n337), .b(new_n339), .o1(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n338), .c(new_n118), .d(new_n337), .o1(\s[8] ));
  nanp02aa1n02x5               g246(.a(new_n117), .b(new_n106), .o1(new_n342));
  aoi012aa1n02x5               g247(.a(new_n122), .b(new_n121), .c(new_n118), .o1(new_n343));
  aoi112aa1n02x5               g248(.a(new_n343), .b(new_n125), .c(new_n109), .d(new_n110), .o1(new_n344));
  aboi22aa1n03x5               g249(.a(new_n183), .b(new_n125), .c(new_n344), .d(new_n342), .out0(\s[9] ));
endmodule


