// Benchmark "adder" written by ABC on Thu Jul 18 05:01:18 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n330,
    new_n332, new_n333, new_n335, new_n337, new_n339, new_n340, new_n341,
    new_n342, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nand22aa1n09x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  oab012aa1d15x5               g003(.a(new_n98), .b(\a[2] ), .c(\b[1] ), .out0(new_n99));
  nand02aa1n03x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  inv040aa1d32x5               g005(.a(\a[3] ), .o1(new_n101));
  inv030aa1d32x5               g006(.a(\b[2] ), .o1(new_n102));
  nand22aa1n04x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nand02aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp03aa1d12x5               g009(.a(new_n103), .b(new_n100), .c(new_n104), .o1(new_n105));
  oa0022aa1n12x5               g010(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n105), .c(new_n99), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor042aa1d18x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  aoi012aa1n02x5               g014(.a(new_n109), .b(\a[8] ), .c(\b[7] ), .o1(new_n110));
  nand02aa1d06x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor042aa1n02x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  norb02aa1n06x4               g017(.a(new_n111), .b(new_n112), .out0(new_n113));
  nor042aa1d18x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1d28x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor042aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nona23aa1n02x4               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nano32aa1n03x7               g023(.a(new_n118), .b(new_n113), .c(new_n110), .d(new_n108), .out0(new_n119));
  nand02aa1d06x5               g024(.a(new_n119), .b(new_n107), .o1(new_n120));
  inv040aa1n03x5               g025(.a(new_n109), .o1(new_n121));
  oaoi03aa1n12x5               g026(.a(\a[8] ), .b(\b[7] ), .c(new_n121), .o1(new_n122));
  nor042aa1n04x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  inv040aa1n08x5               g028(.a(new_n114), .o1(new_n124));
  oaoi03aa1n09x5               g029(.a(\a[6] ), .b(\b[5] ), .c(new_n124), .o1(new_n125));
  tech160nm_fioai012aa1n04x5   g030(.a(new_n116), .b(\b[7] ), .c(\a[8] ), .o1(new_n126));
  aoi112aa1n03x5               g031(.a(new_n126), .b(new_n109), .c(\a[8] ), .d(\b[7] ), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(new_n127), .b(new_n125), .o1(new_n128));
  nona23aa1n02x4               g033(.a(new_n120), .b(new_n128), .c(new_n123), .d(new_n122), .out0(new_n129));
  xnrc02aa1n12x5               g034(.a(\b[9] ), .b(\a[10] ), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n97), .out0(\s[10] ));
  nanp02aa1n02x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n132), .b(new_n133), .out0(new_n134));
  nanp02aa1n02x5               g039(.a(new_n129), .b(new_n97), .o1(new_n135));
  oaoi03aa1n02x5               g040(.a(\a[10] ), .b(\b[9] ), .c(new_n135), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n133), .o1(new_n137));
  inv000aa1d42x5               g042(.a(\a[10] ), .o1(new_n138));
  oaib12aa1n02x5               g043(.a(new_n135), .b(\b[9] ), .c(new_n138), .out0(new_n139));
  aoi022aa1d24x5               g044(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n140));
  nanp03aa1n02x5               g045(.a(new_n139), .b(new_n137), .c(new_n140), .o1(new_n141));
  oa0012aa1n02x5               g046(.a(new_n141), .b(new_n136), .c(new_n134), .o(\s[11] ));
  aob012aa1n02x5               g047(.a(new_n137), .b(new_n139), .c(new_n140), .out0(new_n143));
  nor002aa1n04x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n02x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  aoib12aa1n02x5               g051(.a(new_n133), .b(new_n145), .c(new_n144), .out0(new_n147));
  aoi022aa1n02x5               g052(.a(new_n143), .b(new_n146), .c(new_n141), .d(new_n147), .o1(\s[12] ));
  aoi012aa1n09x5               g053(.a(new_n122), .b(new_n127), .c(new_n125), .o1(new_n149));
  nanb02aa1n06x5               g054(.a(new_n123), .b(new_n97), .out0(new_n150));
  nona23aa1n02x4               g055(.a(new_n134), .b(new_n146), .c(new_n130), .d(new_n150), .out0(new_n151));
  nor002aa1n02x5               g056(.a(\b[9] ), .b(\a[10] ), .o1(new_n152));
  tech160nm_fioai012aa1n03p5x5 g057(.a(new_n140), .b(new_n152), .c(new_n123), .o1(new_n153));
  nona22aa1n03x5               g058(.a(new_n153), .b(new_n144), .c(new_n133), .out0(new_n154));
  and002aa1n02x5               g059(.a(new_n154), .b(new_n145), .o(new_n155));
  inv000aa1n02x5               g060(.a(new_n155), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n151), .c(new_n120), .d(new_n149), .o1(new_n157));
  xnrc02aa1n12x5               g062(.a(\b[12] ), .b(\a[13] ), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(new_n120), .b(new_n149), .o1(new_n160));
  nona23aa1n03x5               g065(.a(new_n132), .b(new_n145), .c(new_n144), .d(new_n133), .out0(new_n161));
  nor043aa1n03x5               g066(.a(new_n161), .b(new_n150), .c(new_n130), .o1(new_n162));
  aoi112aa1n02x5               g067(.a(new_n159), .b(new_n155), .c(new_n160), .d(new_n162), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n163), .b(new_n157), .c(new_n159), .o1(\s[13] ));
  inv000aa1d42x5               g069(.a(\a[13] ), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[12] ), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(new_n166), .b(new_n165), .o1(new_n167));
  nanp02aa1n02x5               g072(.a(new_n157), .b(new_n159), .o1(new_n168));
  tech160nm_fixnrc02aa1n02p5x5 g073(.a(\b[13] ), .b(\a[14] ), .out0(new_n169));
  xobna2aa1n03x5               g074(.a(new_n169), .b(new_n168), .c(new_n167), .out0(\s[14] ));
  norp02aa1n02x5               g075(.a(new_n169), .b(new_n158), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(new_n157), .b(new_n171), .o1(new_n172));
  aoi112aa1n09x5               g077(.a(\b[12] ), .b(\a[13] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n173));
  oab012aa1n12x5               g078(.a(new_n173), .b(\a[14] ), .c(\b[13] ), .out0(new_n174));
  nor042aa1n09x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nanp02aa1n04x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n172), .c(new_n174), .out0(\s[15] ));
  aob012aa1n02x5               g083(.a(new_n177), .b(new_n172), .c(new_n174), .out0(new_n179));
  nor042aa1n06x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nand02aa1d06x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n181), .b(new_n180), .out0(new_n182));
  aoib12aa1n02x5               g087(.a(new_n175), .b(new_n181), .c(new_n180), .out0(new_n183));
  aobi12aa1n02x5               g088(.a(new_n174), .b(new_n157), .c(new_n171), .out0(new_n184));
  oaoi03aa1n02x5               g089(.a(\a[15] ), .b(\b[14] ), .c(new_n184), .o1(new_n185));
  aoi022aa1n03x5               g090(.a(new_n185), .b(new_n182), .c(new_n179), .d(new_n183), .o1(\s[16] ));
  nano32aa1n03x7               g091(.a(new_n151), .b(new_n182), .c(new_n171), .d(new_n177), .out0(new_n187));
  nanp02aa1n02x5               g092(.a(new_n160), .b(new_n187), .o1(new_n188));
  nona23aa1n09x5               g093(.a(new_n181), .b(new_n176), .c(new_n175), .d(new_n180), .out0(new_n189));
  nona32aa1n09x5               g094(.a(new_n162), .b(new_n189), .c(new_n169), .d(new_n158), .out0(new_n190));
  nanb03aa1n06x5               g095(.a(new_n180), .b(new_n181), .c(new_n176), .out0(new_n191));
  aoi022aa1n02x5               g096(.a(new_n166), .b(new_n165), .c(\a[12] ), .d(\b[11] ), .o1(new_n192));
  oai022aa1d24x5               g097(.a(new_n165), .b(new_n166), .c(\b[13] ), .d(\a[14] ), .o1(new_n193));
  aoi012aa1n02x5               g098(.a(new_n175), .b(\a[14] ), .c(\b[13] ), .o1(new_n194));
  nano23aa1n09x5               g099(.a(new_n191), .b(new_n193), .c(new_n192), .d(new_n194), .out0(new_n195));
  tech160nm_fiaoi012aa1n03p5x5 g100(.a(new_n180), .b(new_n175), .c(new_n181), .o1(new_n196));
  tech160nm_fioai012aa1n04x5   g101(.a(new_n196), .b(new_n189), .c(new_n174), .o1(new_n197));
  aoi012aa1n12x5               g102(.a(new_n197), .b(new_n195), .c(new_n154), .o1(new_n198));
  aoai13aa1n12x5               g103(.a(new_n198), .b(new_n190), .c(new_n120), .d(new_n149), .o1(new_n199));
  xorc02aa1n02x5               g104(.a(\a[17] ), .b(\b[16] ), .out0(new_n200));
  norp02aa1n02x5               g105(.a(new_n189), .b(new_n174), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(new_n200), .b(new_n196), .out0(new_n202));
  aoi112aa1n02x5               g107(.a(new_n201), .b(new_n202), .c(new_n195), .d(new_n154), .o1(new_n203));
  aoi022aa1n02x5               g108(.a(new_n199), .b(new_n200), .c(new_n188), .d(new_n203), .o1(\s[17] ));
  inv020aa1n12x5               g109(.a(\a[17] ), .o1(new_n205));
  nanb02aa1n12x5               g110(.a(\b[16] ), .b(new_n205), .out0(new_n206));
  nanp02aa1n02x5               g111(.a(new_n199), .b(new_n200), .o1(new_n207));
  xorc02aa1n02x5               g112(.a(\a[18] ), .b(\b[17] ), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n207), .c(new_n206), .out0(\s[18] ));
  inv020aa1n04x5               g114(.a(\a[18] ), .o1(new_n210));
  xroi22aa1d06x4               g115(.a(new_n205), .b(\b[16] ), .c(new_n210), .d(\b[17] ), .out0(new_n211));
  oaoi03aa1n12x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n206), .o1(new_n212));
  xorc02aa1n12x5               g117(.a(\a[19] ), .b(\b[18] ), .out0(new_n213));
  aoai13aa1n06x5               g118(.a(new_n213), .b(new_n212), .c(new_n199), .d(new_n211), .o1(new_n214));
  aoi112aa1n02x5               g119(.a(new_n213), .b(new_n212), .c(new_n199), .d(new_n211), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n214), .b(new_n215), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  xorc02aa1n12x5               g122(.a(\a[20] ), .b(\b[19] ), .out0(new_n218));
  orn002aa1n03x5               g123(.a(\a[19] ), .b(\b[18] ), .o(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  nanp02aa1n02x5               g125(.a(new_n214), .b(new_n219), .o1(new_n221));
  aoi022aa1n02x5               g126(.a(new_n221), .b(new_n218), .c(new_n214), .d(new_n220), .o1(\s[20] ));
  nand23aa1n06x5               g127(.a(new_n211), .b(new_n213), .c(new_n218), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  nand23aa1n06x5               g129(.a(new_n212), .b(new_n213), .c(new_n218), .o1(new_n225));
  oao003aa1n03x5               g130(.a(\a[20] ), .b(\b[19] ), .c(new_n219), .carry(new_n226));
  nanp02aa1n02x5               g131(.a(new_n225), .b(new_n226), .o1(new_n227));
  xorc02aa1n02x5               g132(.a(\a[21] ), .b(\b[20] ), .out0(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n227), .c(new_n199), .d(new_n224), .o1(new_n229));
  nano22aa1n02x4               g134(.a(new_n228), .b(new_n225), .c(new_n226), .out0(new_n230));
  aobi12aa1n02x5               g135(.a(new_n230), .b(new_n199), .c(new_n224), .out0(new_n231));
  norb02aa1n02x5               g136(.a(new_n229), .b(new_n231), .out0(\s[21] ));
  xorc02aa1n02x5               g137(.a(\a[22] ), .b(\b[21] ), .out0(new_n233));
  norp02aa1n02x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norp02aa1n02x5               g139(.a(new_n233), .b(new_n234), .o1(new_n235));
  inv040aa1d30x5               g140(.a(\a[21] ), .o1(new_n236));
  oaib12aa1n02x5               g141(.a(new_n229), .b(\b[20] ), .c(new_n236), .out0(new_n237));
  aoi022aa1n02x5               g142(.a(new_n237), .b(new_n233), .c(new_n229), .d(new_n235), .o1(\s[22] ));
  inv040aa1d32x5               g143(.a(\a[22] ), .o1(new_n239));
  xroi22aa1d06x4               g144(.a(new_n236), .b(\b[20] ), .c(new_n239), .d(\b[21] ), .out0(new_n240));
  inv020aa1n04x5               g145(.a(new_n240), .o1(new_n241));
  nona22aa1n06x5               g146(.a(new_n199), .b(new_n223), .c(new_n241), .out0(new_n242));
  oai022aa1n02x5               g147(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n243));
  oaib12aa1n06x5               g148(.a(new_n243), .b(new_n239), .c(\b[21] ), .out0(new_n244));
  aoai13aa1n12x5               g149(.a(new_n244), .b(new_n241), .c(new_n225), .d(new_n226), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xorc02aa1n12x5               g151(.a(\a[23] ), .b(\b[22] ), .out0(new_n247));
  aob012aa1n03x5               g152(.a(new_n247), .b(new_n242), .c(new_n246), .out0(new_n248));
  nanb02aa1n02x5               g153(.a(new_n247), .b(new_n244), .out0(new_n249));
  aoi012aa1n02x5               g154(.a(new_n249), .b(new_n227), .c(new_n240), .o1(new_n250));
  aobi12aa1n02x7               g155(.a(new_n248), .b(new_n250), .c(new_n242), .out0(\s[23] ));
  xorc02aa1n02x5               g156(.a(\a[24] ), .b(\b[23] ), .out0(new_n252));
  nor042aa1n06x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  norp02aa1n02x5               g158(.a(new_n252), .b(new_n253), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n253), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n247), .o1(new_n256));
  aoai13aa1n02x5               g161(.a(new_n255), .b(new_n256), .c(new_n242), .d(new_n246), .o1(new_n257));
  aoi022aa1n02x7               g162(.a(new_n257), .b(new_n252), .c(new_n248), .d(new_n254), .o1(\s[24] ));
  and002aa1n12x5               g163(.a(new_n252), .b(new_n247), .o(new_n259));
  nona23aa1n06x5               g164(.a(new_n199), .b(new_n259), .c(new_n241), .d(new_n223), .out0(new_n260));
  oaoi03aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .c(new_n255), .o1(new_n261));
  tech160nm_fiaoi012aa1n05x5   g166(.a(new_n261), .b(new_n245), .c(new_n259), .o1(new_n262));
  inv040aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  aobi12aa1n02x5               g168(.a(new_n198), .b(new_n160), .c(new_n187), .out0(new_n264));
  nano32aa1n03x7               g169(.a(new_n264), .b(new_n259), .c(new_n224), .d(new_n240), .out0(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  oai012aa1n06x5               g171(.a(new_n266), .b(new_n265), .c(new_n263), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n266), .b(new_n261), .c(new_n245), .d(new_n259), .o1(new_n268));
  aobi12aa1n02x7               g173(.a(new_n267), .b(new_n268), .c(new_n260), .out0(\s[25] ));
  xorc02aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .out0(new_n270));
  norp02aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  norp02aa1n02x5               g176(.a(new_n270), .b(new_n271), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n266), .o1(new_n274));
  aoai13aa1n04x5               g179(.a(new_n273), .b(new_n274), .c(new_n260), .d(new_n262), .o1(new_n275));
  aoi022aa1n03x5               g180(.a(new_n275), .b(new_n270), .c(new_n267), .d(new_n272), .o1(\s[26] ));
  and002aa1n02x5               g181(.a(new_n270), .b(new_n266), .o(new_n277));
  aoai13aa1n12x5               g182(.a(new_n277), .b(new_n261), .c(new_n245), .d(new_n259), .o1(new_n278));
  nano32aa1n06x5               g183(.a(new_n223), .b(new_n277), .c(new_n240), .d(new_n259), .out0(new_n279));
  nanp02aa1n02x5               g184(.a(new_n199), .b(new_n279), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(\b[25] ), .b(\a[26] ), .o1(new_n281));
  oai022aa1n02x5               g186(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(new_n282), .b(new_n281), .o1(new_n283));
  nand23aa1n06x5               g188(.a(new_n280), .b(new_n278), .c(new_n283), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  aoi122aa1n02x5               g190(.a(new_n285), .b(new_n281), .c(new_n282), .d(new_n199), .e(new_n279), .o1(new_n286));
  aoi022aa1n03x5               g191(.a(new_n286), .b(new_n278), .c(new_n284), .d(new_n285), .o1(\s[27] ));
  nanp02aa1n03x5               g192(.a(new_n284), .b(new_n285), .o1(new_n288));
  xorc02aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .out0(new_n289));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  norp02aa1n02x5               g195(.a(new_n289), .b(new_n290), .o1(new_n291));
  aoi022aa1n02x5               g196(.a(new_n199), .b(new_n279), .c(new_n281), .d(new_n282), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n290), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n285), .o1(new_n294));
  aoai13aa1n02x5               g199(.a(new_n293), .b(new_n294), .c(new_n292), .d(new_n278), .o1(new_n295));
  aoi022aa1n03x5               g200(.a(new_n295), .b(new_n289), .c(new_n288), .d(new_n291), .o1(\s[28] ));
  and002aa1n02x5               g201(.a(new_n289), .b(new_n285), .o(new_n297));
  nand22aa1n03x5               g202(.a(new_n284), .b(new_n297), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(\a[28] ), .o1(new_n300));
  inv000aa1d42x5               g205(.a(\b[27] ), .o1(new_n301));
  aoi112aa1n02x5               g206(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n302));
  aoi112aa1n02x5               g207(.a(new_n299), .b(new_n302), .c(new_n300), .d(new_n301), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n297), .o1(new_n304));
  aoi012aa1n02x5               g209(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n305));
  aoai13aa1n02x5               g210(.a(new_n305), .b(new_n304), .c(new_n292), .d(new_n278), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n299), .c(new_n298), .d(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g213(.a(new_n294), .b(new_n289), .c(new_n299), .out0(new_n309));
  nanp02aa1n03x5               g214(.a(new_n284), .b(new_n309), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .out0(new_n311));
  aoi012aa1n02x5               g216(.a(new_n305), .b(\a[29] ), .c(\b[28] ), .o1(new_n312));
  oabi12aa1n02x5               g217(.a(new_n311), .b(\a[29] ), .c(\b[28] ), .out0(new_n313));
  norp02aa1n02x5               g218(.a(new_n313), .b(new_n312), .o1(new_n314));
  inv000aa1n02x5               g219(.a(new_n309), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .carry(new_n316));
  aoai13aa1n02x5               g221(.a(new_n316), .b(new_n315), .c(new_n292), .d(new_n278), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n311), .c(new_n310), .d(new_n314), .o1(\s[30] ));
  nano32aa1n02x4               g223(.a(new_n294), .b(new_n311), .c(new_n289), .d(new_n299), .out0(new_n319));
  nanp02aa1n03x5               g224(.a(new_n284), .b(new_n319), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[31] ), .b(\b[30] ), .out0(new_n321));
  nanp02aa1n02x5               g226(.a(\b[29] ), .b(\a[30] ), .o1(new_n322));
  oai022aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(\b[29] ), .d(\a[30] ), .o1(new_n323));
  oaoi13aa1n02x5               g228(.a(new_n321), .b(new_n322), .c(new_n312), .d(new_n323), .o1(new_n324));
  inv000aa1n02x5               g229(.a(new_n319), .o1(new_n325));
  oai012aa1n02x5               g230(.a(new_n322), .b(new_n312), .c(new_n323), .o1(new_n326));
  aoai13aa1n02x5               g231(.a(new_n326), .b(new_n325), .c(new_n292), .d(new_n278), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n321), .c(new_n320), .d(new_n324), .o1(\s[31] ));
  norp02aa1n02x5               g233(.a(new_n105), .b(new_n99), .o1(new_n329));
  aboi22aa1n03x5               g234(.a(new_n99), .b(new_n100), .c(new_n103), .d(new_n104), .out0(new_n330));
  norp02aa1n02x5               g235(.a(new_n330), .b(new_n329), .o1(\s[3] ));
  inv000aa1n03x5               g236(.a(new_n329), .o1(new_n332));
  xorc02aa1n02x5               g237(.a(\a[4] ), .b(\b[3] ), .out0(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n332), .c(new_n103), .out0(\s[4] ));
  norb02aa1n02x5               g239(.a(new_n115), .b(new_n114), .out0(new_n335));
  xobna2aa1n03x5               g240(.a(new_n335), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  nanp03aa1n02x5               g241(.a(new_n107), .b(new_n108), .c(new_n335), .o1(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n113), .b(new_n337), .c(new_n124), .out0(\s[6] ));
  and003aa1n02x5               g243(.a(new_n113), .b(new_n335), .c(new_n108), .o(new_n339));
  norb02aa1n02x5               g244(.a(new_n116), .b(new_n109), .out0(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n125), .c(new_n339), .d(new_n107), .o1(new_n341));
  aoi112aa1n02x5               g246(.a(new_n340), .b(new_n125), .c(new_n339), .d(new_n107), .o1(new_n342));
  norb02aa1n02x5               g247(.a(new_n341), .b(new_n342), .out0(\s[7] ));
  xorc02aa1n02x5               g248(.a(\a[8] ), .b(\b[7] ), .out0(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n344), .b(new_n341), .c(new_n121), .out0(\s[8] ));
  nona23aa1n02x4               g250(.a(new_n120), .b(new_n128), .c(new_n150), .d(new_n122), .out0(new_n346));
  aob012aa1n02x5               g251(.a(new_n346), .b(new_n160), .c(new_n150), .out0(\s[9] ));
endmodule


