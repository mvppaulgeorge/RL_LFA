// Benchmark "adder" written by ABC on Wed Jul 17 19:22:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n314, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n334, new_n337, new_n338, new_n339, new_n340,
    new_n342, new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n12x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nanb02aa1n09x5               g005(.a(new_n99), .b(new_n100), .out0(new_n101));
  nand02aa1n03x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai112aa1n06x5               g007(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n103));
  nanp02aa1n09x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nand42aa1d28x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n04x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb03aa1n09x5               g011(.a(new_n105), .b(new_n99), .c(new_n106), .out0(new_n107));
  oai012aa1d24x5               g012(.a(new_n107), .b(new_n104), .c(new_n101), .o1(new_n108));
  nand02aa1d28x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  aoi022aa1d24x5               g014(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n110));
  oai112aa1n03x5               g015(.a(new_n110), .b(new_n109), .c(\b[7] ), .d(\a[8] ), .o1(new_n111));
  tech160nm_fixnrc02aa1n02p5x5 g016(.a(\b[4] ), .b(\a[5] ), .out0(new_n112));
  oai122aa1n12x5               g017(.a(new_n105), .b(\a[7] ), .c(\b[6] ), .d(\a[6] ), .e(\b[5] ), .o1(new_n113));
  nor043aa1n06x5               g018(.a(new_n111), .b(new_n112), .c(new_n113), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n08x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand23aa1n06x5               g021(.a(new_n115), .b(new_n109), .c(new_n116), .o1(new_n117));
  oai022aa1d18x5               g022(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n118));
  nanp02aa1n04x5               g023(.a(new_n118), .b(new_n116), .o1(new_n119));
  nor042aa1n03x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nor042aa1n03x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  norb03aa1d15x5               g026(.a(new_n109), .b(new_n121), .c(new_n120), .out0(new_n122));
  oai013aa1d12x5               g027(.a(new_n119), .b(new_n122), .c(new_n117), .d(new_n118), .o1(new_n123));
  nanp02aa1n04x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n97), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n123), .c(new_n114), .d(new_n108), .o1(new_n126));
  norp02aa1n12x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanb02aa1n02x5               g033(.a(new_n127), .b(new_n128), .out0(new_n129));
  xobna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  tech160nm_fioai012aa1n05x5   g035(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n131));
  aoai13aa1n04x5               g036(.a(new_n131), .b(new_n129), .c(new_n126), .d(new_n98), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d24x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand02aa1d06x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norp02aa1n12x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanp02aa1n06x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aoai13aa1n03x5               g043(.a(new_n138), .b(new_n134), .c(new_n132), .d(new_n135), .o1(new_n139));
  aoi112aa1n03x5               g044(.a(new_n134), .b(new_n138), .c(new_n132), .d(new_n135), .o1(new_n140));
  norb02aa1n02x7               g045(.a(new_n139), .b(new_n140), .out0(\s[12] ));
  nona23aa1n09x5               g046(.a(new_n137), .b(new_n135), .c(new_n134), .d(new_n136), .out0(new_n142));
  nona23aa1n09x5               g047(.a(new_n128), .b(new_n124), .c(new_n97), .d(new_n127), .out0(new_n143));
  nor042aa1n02x5               g048(.a(new_n143), .b(new_n142), .o1(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n123), .c(new_n114), .d(new_n108), .o1(new_n145));
  inv020aa1n02x5               g050(.a(new_n131), .o1(new_n146));
  nano23aa1n09x5               g051(.a(new_n134), .b(new_n136), .c(new_n137), .d(new_n135), .out0(new_n147));
  oa0012aa1n02x5               g052(.a(new_n137), .b(new_n136), .c(new_n134), .o(new_n148));
  aoi012aa1n06x5               g053(.a(new_n148), .b(new_n147), .c(new_n146), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n145), .b(new_n149), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1n20x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  tech160nm_fiaoi012aa1n05x5   g058(.a(new_n152), .b(new_n150), .c(new_n153), .o1(new_n154));
  xnrb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n06x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nand42aa1n08x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nona23aa1n09x5               g062(.a(new_n157), .b(new_n153), .c(new_n152), .d(new_n156), .out0(new_n158));
  tech160nm_fiaoi012aa1n03p5x5 g063(.a(new_n156), .b(new_n152), .c(new_n157), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n159), .b(new_n158), .c(new_n145), .d(new_n149), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nanp02aa1n04x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nor042aa1d18x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nand02aa1d12x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nanb02aa1d24x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n162), .c(new_n160), .d(new_n163), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n162), .b(new_n167), .c(new_n160), .d(new_n163), .o1(new_n169));
  norb02aa1n02x7               g074(.a(new_n168), .b(new_n169), .out0(\s[16] ));
  aoi012aa1d24x5               g075(.a(new_n123), .b(new_n114), .c(new_n108), .o1(new_n171));
  nona23aa1n09x5               g076(.a(new_n165), .b(new_n163), .c(new_n162), .d(new_n164), .out0(new_n172));
  nor042aa1n02x5               g077(.a(new_n172), .b(new_n158), .o1(new_n173));
  nand22aa1n03x5               g078(.a(new_n173), .b(new_n144), .o1(new_n174));
  oabi12aa1n03x5               g079(.a(new_n148), .b(new_n131), .c(new_n142), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n164), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(new_n162), .b(new_n165), .o1(new_n177));
  oai112aa1n03x5               g082(.a(new_n177), .b(new_n176), .c(new_n172), .d(new_n159), .o1(new_n178));
  aoi012aa1n06x5               g083(.a(new_n178), .b(new_n175), .c(new_n173), .o1(new_n179));
  oai012aa1d24x5               g084(.a(new_n179), .b(new_n171), .c(new_n174), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g086(.a(\a[18] ), .o1(new_n182));
  inv030aa1d32x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  oaoi03aa1n03x5               g089(.a(new_n183), .b(new_n184), .c(new_n180), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n182), .out0(\s[18] ));
  xroi22aa1d06x4               g091(.a(new_n183), .b(\b[16] ), .c(new_n182), .d(\b[17] ), .out0(new_n187));
  inv000aa1d42x5               g092(.a(\b[17] ), .o1(new_n188));
  norp02aa1n02x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  oao003aa1n02x5               g094(.a(new_n182), .b(new_n188), .c(new_n189), .carry(new_n190));
  tech160nm_fiaoi012aa1n05x5   g095(.a(new_n190), .b(new_n180), .c(new_n187), .o1(new_n191));
  nor042aa1d18x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  nand02aa1n06x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n191), .b(new_n194), .c(new_n193), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norb02aa1n12x5               g101(.a(new_n194), .b(new_n192), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n190), .c(new_n180), .d(new_n187), .o1(new_n198));
  nor002aa1d32x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1d28x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1d27x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  tech160nm_fiaoi012aa1n03p5x5 g107(.a(new_n202), .b(new_n198), .c(new_n193), .o1(new_n203));
  nona22aa1n02x5               g108(.a(new_n198), .b(new_n201), .c(new_n192), .out0(new_n204));
  norb02aa1n03x4               g109(.a(new_n204), .b(new_n203), .out0(\s[20] ));
  nanb02aa1n02x5               g110(.a(new_n106), .b(new_n105), .out0(new_n206));
  aoi113aa1n03x7               g111(.a(new_n206), .b(new_n99), .c(new_n103), .d(new_n100), .e(new_n102), .o1(new_n207));
  norp02aa1n02x5               g112(.a(\b[7] ), .b(\a[8] ), .o1(new_n208));
  inv040aa1n03x5               g113(.a(new_n117), .o1(new_n209));
  tech160nm_fixorc02aa1n03p5x5 g114(.a(\a[5] ), .b(\b[4] ), .out0(new_n210));
  nona23aa1n03x5               g115(.a(new_n209), .b(new_n210), .c(new_n113), .d(new_n208), .out0(new_n211));
  inv000aa1n02x5               g116(.a(new_n119), .o1(new_n212));
  nor003aa1n03x5               g117(.a(new_n122), .b(new_n118), .c(new_n117), .o1(new_n213));
  nor042aa1n02x5               g118(.a(new_n213), .b(new_n212), .o1(new_n214));
  oai012aa1n06x5               g119(.a(new_n214), .b(new_n211), .c(new_n207), .o1(new_n215));
  nano23aa1n02x5               g120(.a(new_n152), .b(new_n156), .c(new_n157), .d(new_n153), .out0(new_n216));
  nano23aa1n06x5               g121(.a(new_n172), .b(new_n143), .c(new_n147), .d(new_n216), .out0(new_n217));
  nanb02aa1n02x5               g122(.a(new_n162), .b(new_n163), .out0(new_n218));
  nona22aa1n03x5               g123(.a(new_n216), .b(new_n218), .c(new_n166), .out0(new_n219));
  nor043aa1n02x5               g124(.a(new_n159), .b(new_n218), .c(new_n166), .o1(new_n220));
  nano22aa1n03x7               g125(.a(new_n220), .b(new_n176), .c(new_n177), .out0(new_n221));
  oai012aa1n12x5               g126(.a(new_n221), .b(new_n149), .c(new_n219), .o1(new_n222));
  nano23aa1n09x5               g127(.a(new_n192), .b(new_n199), .c(new_n200), .d(new_n194), .out0(new_n223));
  nand22aa1n09x5               g128(.a(new_n187), .b(new_n223), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n222), .c(new_n215), .d(new_n217), .o1(new_n226));
  aoi112aa1n09x5               g131(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n227));
  nor042aa1n02x5               g132(.a(\b[17] ), .b(\a[18] ), .o1(new_n228));
  aoi112aa1n09x5               g133(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n229));
  oai112aa1n06x5               g134(.a(new_n197), .b(new_n201), .c(new_n229), .d(new_n228), .o1(new_n230));
  nona22aa1d18x5               g135(.a(new_n230), .b(new_n227), .c(new_n199), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  nor002aa1d32x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  nand42aa1n10x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n06x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n226), .c(new_n232), .out0(\s[21] ));
  inv000aa1d42x5               g141(.a(new_n233), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n235), .b(new_n231), .c(new_n180), .d(new_n225), .o1(new_n238));
  nor042aa1n04x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  tech160nm_finand02aa1n05x5   g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nanb02aa1n02x5               g145(.a(new_n239), .b(new_n240), .out0(new_n241));
  aoi012aa1n03x5               g146(.a(new_n241), .b(new_n238), .c(new_n237), .o1(new_n242));
  aobi12aa1n06x5               g147(.a(new_n235), .b(new_n226), .c(new_n232), .out0(new_n243));
  nano22aa1n02x4               g148(.a(new_n243), .b(new_n237), .c(new_n241), .out0(new_n244));
  norp02aa1n03x5               g149(.a(new_n242), .b(new_n244), .o1(\s[22] ));
  nano23aa1n06x5               g150(.a(new_n233), .b(new_n239), .c(new_n240), .d(new_n234), .out0(new_n246));
  and003aa1n02x5               g151(.a(new_n187), .b(new_n246), .c(new_n223), .o(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n222), .c(new_n215), .d(new_n217), .o1(new_n248));
  oaoi03aa1n02x5               g153(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .o1(new_n249));
  tech160nm_fiaoi012aa1n04x5   g154(.a(new_n249), .b(new_n231), .c(new_n246), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  xnbna2aa1n03x5               g156(.a(new_n251), .b(new_n248), .c(new_n250), .out0(\s[23] ));
  orn002aa1n02x5               g157(.a(\a[23] ), .b(\b[22] ), .o(new_n253));
  inv040aa1n02x5               g158(.a(new_n250), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n251), .b(new_n254), .c(new_n180), .d(new_n247), .o1(new_n255));
  norp02aa1n09x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nand42aa1n08x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  norb02aa1d21x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  aoi012aa1n03x5               g164(.a(new_n259), .b(new_n255), .c(new_n253), .o1(new_n260));
  xnrc02aa1n12x5               g165(.a(\b[22] ), .b(\a[23] ), .out0(new_n261));
  tech160nm_fiaoi012aa1n02p5x5 g166(.a(new_n261), .b(new_n248), .c(new_n250), .o1(new_n262));
  nano22aa1n02x4               g167(.a(new_n262), .b(new_n253), .c(new_n259), .out0(new_n263));
  norp02aa1n02x5               g168(.a(new_n260), .b(new_n263), .o1(\s[24] ));
  norb02aa1n03x5               g169(.a(new_n258), .b(new_n261), .out0(new_n265));
  nano22aa1n09x5               g170(.a(new_n224), .b(new_n246), .c(new_n265), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n222), .c(new_n215), .d(new_n217), .o1(new_n267));
  nano23aa1n06x5               g172(.a(new_n261), .b(new_n241), .c(new_n258), .d(new_n235), .out0(new_n268));
  aoi112aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n269));
  aoi112aa1n02x7               g174(.a(\b[20] ), .b(\a[21] ), .c(\a[22] ), .d(\b[21] ), .o1(new_n270));
  oai112aa1n02x7               g175(.a(new_n251), .b(new_n258), .c(new_n270), .d(new_n239), .o1(new_n271));
  nona22aa1n02x4               g176(.a(new_n271), .b(new_n269), .c(new_n256), .out0(new_n272));
  aoi012aa1n09x5               g177(.a(new_n272), .b(new_n231), .c(new_n268), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n267), .c(new_n273), .out0(\s[25] ));
  orn002aa1n02x5               g180(.a(\a[25] ), .b(\b[24] ), .o(new_n276));
  inv020aa1n08x5               g181(.a(new_n273), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n274), .b(new_n277), .c(new_n180), .d(new_n266), .o1(new_n278));
  tech160nm_fixnrc02aa1n05x5   g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  aoi012aa1n03x5               g184(.a(new_n279), .b(new_n278), .c(new_n276), .o1(new_n280));
  aobi12aa1n06x5               g185(.a(new_n274), .b(new_n267), .c(new_n273), .out0(new_n281));
  nano22aa1n03x7               g186(.a(new_n281), .b(new_n276), .c(new_n279), .out0(new_n282));
  nor002aa1n02x5               g187(.a(new_n280), .b(new_n282), .o1(\s[26] ));
  norb02aa1n09x5               g188(.a(new_n274), .b(new_n279), .out0(new_n284));
  nano32aa1d12x5               g189(.a(new_n224), .b(new_n284), .c(new_n246), .d(new_n265), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n222), .c(new_n215), .d(new_n217), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n199), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n227), .o1(new_n288));
  nanp03aa1n03x5               g193(.a(new_n246), .b(new_n251), .c(new_n258), .o1(new_n289));
  aoi013aa1n06x4               g194(.a(new_n289), .b(new_n230), .c(new_n288), .d(new_n287), .o1(new_n290));
  oaoi03aa1n12x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n276), .o1(new_n291));
  oaoi13aa1n09x5               g196(.a(new_n291), .b(new_n284), .c(new_n290), .d(new_n272), .o1(new_n292));
  xorc02aa1n12x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  xnbna2aa1n03x5               g198(.a(new_n293), .b(new_n292), .c(new_n286), .out0(\s[27] ));
  norp02aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  inv040aa1n03x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n284), .b(new_n272), .c(new_n231), .d(new_n268), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n291), .o1(new_n298));
  nand02aa1d06x5               g203(.a(new_n297), .b(new_n298), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n293), .b(new_n299), .c(new_n180), .d(new_n285), .o1(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[27] ), .b(\a[28] ), .out0(new_n301));
  aoi012aa1n03x5               g206(.a(new_n301), .b(new_n300), .c(new_n296), .o1(new_n302));
  aobi12aa1n02x7               g207(.a(new_n293), .b(new_n292), .c(new_n286), .out0(new_n303));
  nano22aa1n02x4               g208(.a(new_n303), .b(new_n296), .c(new_n301), .out0(new_n304));
  nor002aa1n02x5               g209(.a(new_n302), .b(new_n304), .o1(\s[28] ));
  norb02aa1n02x5               g210(.a(new_n293), .b(new_n301), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n299), .c(new_n180), .d(new_n285), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n296), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[28] ), .b(\a[29] ), .out0(new_n309));
  aoi012aa1n02x7               g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  aobi12aa1n02x7               g215(.a(new_n306), .b(new_n292), .c(new_n286), .out0(new_n311));
  nano22aa1n02x4               g216(.a(new_n311), .b(new_n308), .c(new_n309), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n310), .b(new_n312), .o1(\s[29] ));
  nanp02aa1n02x5               g218(.a(\b[0] ), .b(\a[1] ), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g220(.a(new_n293), .b(new_n309), .c(new_n301), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n299), .c(new_n180), .d(new_n285), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .carry(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .out0(new_n319));
  aoi012aa1n02x7               g224(.a(new_n319), .b(new_n317), .c(new_n318), .o1(new_n320));
  aobi12aa1n02x7               g225(.a(new_n316), .b(new_n292), .c(new_n286), .out0(new_n321));
  nano22aa1n02x4               g226(.a(new_n321), .b(new_n318), .c(new_n319), .out0(new_n322));
  norp02aa1n03x5               g227(.a(new_n320), .b(new_n322), .o1(\s[30] ));
  nona32aa1n02x4               g228(.a(new_n293), .b(new_n319), .c(new_n309), .d(new_n301), .out0(new_n324));
  aoi012aa1n02x7               g229(.a(new_n324), .b(new_n292), .c(new_n286), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .c(new_n318), .carry(new_n326));
  xnrc02aa1n02x5               g231(.a(\b[30] ), .b(\a[31] ), .out0(new_n327));
  nano22aa1n03x5               g232(.a(new_n325), .b(new_n326), .c(new_n327), .out0(new_n328));
  inv000aa1n02x5               g233(.a(new_n324), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n299), .c(new_n180), .d(new_n285), .o1(new_n330));
  aoi012aa1n02x7               g235(.a(new_n327), .b(new_n330), .c(new_n326), .o1(new_n331));
  nor002aa1n02x5               g236(.a(new_n331), .b(new_n328), .o1(\s[31] ));
  xnbna2aa1n03x5               g237(.a(new_n101), .b(new_n103), .c(new_n102), .out0(\s[3] ));
  aoi013aa1n02x4               g238(.a(new_n99), .b(new_n103), .c(new_n102), .d(new_n100), .o1(new_n334));
  oaib12aa1n02x5               g239(.a(new_n108), .b(new_n334), .c(new_n206), .out0(\s[4] ));
  xnbna2aa1n03x5               g240(.a(new_n112), .b(new_n108), .c(new_n105), .out0(\s[5] ));
  norb02aa1n02x5               g241(.a(new_n109), .b(new_n121), .out0(new_n337));
  aoi013aa1n02x4               g242(.a(new_n120), .b(new_n108), .c(new_n105), .d(new_n210), .o1(new_n338));
  nanp03aa1n02x5               g243(.a(new_n108), .b(new_n105), .c(new_n210), .o1(new_n339));
  nanp02aa1n02x5               g244(.a(new_n339), .b(new_n122), .o1(new_n340));
  oai012aa1n02x5               g245(.a(new_n340), .b(new_n338), .c(new_n337), .o1(\s[6] ));
  nanp02aa1n02x5               g246(.a(new_n340), .b(new_n109), .o1(new_n342));
  xnrb03aa1n02x5               g247(.a(new_n342), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g248(.a(\a[7] ), .b(\b[6] ), .c(new_n342), .o1(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g250(.a(new_n171), .b(new_n124), .c(new_n98), .out0(\s[9] ));
endmodule


