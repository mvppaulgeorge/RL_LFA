// Benchmark "adder" written by ABC on Thu Jul 18 11:20:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n330, new_n332, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n04x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n06x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  aoi012aa1n12x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor022aa1n08x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand42aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n03x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  tech160nm_fioai012aa1n03p5x5 g015(.a(new_n107), .b(new_n108), .c(new_n106), .o1(new_n111));
  tech160nm_fioai012aa1n03p5x5 g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[6] ), .o1(new_n113));
  nanb02aa1d36x5               g018(.a(\a[7] ), .b(new_n113), .out0(new_n114));
  nand42aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  tech160nm_fixorc02aa1n05x5   g020(.a(\a[5] ), .b(\b[4] ), .out0(new_n116));
  nand02aa1d16x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1n04x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[8] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[7] ), .o1(new_n120));
  nand42aa1n02x5               g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  and002aa1n12x5               g026(.a(\b[7] ), .b(\a[8] ), .o(new_n122));
  nona23aa1n02x4               g027(.a(new_n121), .b(new_n117), .c(new_n122), .d(new_n118), .out0(new_n123));
  nano32aa1n03x7               g028(.a(new_n123), .b(new_n116), .c(new_n115), .d(new_n114), .out0(new_n124));
  nor042aa1n03x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  aoai13aa1n06x5               g030(.a(new_n115), .b(new_n118), .c(new_n125), .d(new_n117), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n121), .b(new_n122), .c(new_n126), .d(new_n114), .o1(new_n127));
  nand42aa1n08x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n03x5               g034(.a(new_n129), .b(new_n127), .c(new_n124), .d(new_n112), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  xnrc02aa1n12x5               g036(.a(\b[10] ), .b(\a[11] ), .out0(new_n132));
  nona22aa1n02x4               g037(.a(new_n130), .b(new_n100), .c(new_n97), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n132), .b(new_n133), .c(new_n98), .out0(\s[11] ));
  inv000aa1d42x5               g039(.a(\a[12] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(\a[11] ), .o1(new_n136));
  inv000aa1d42x5               g041(.a(\b[10] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n98), .b(new_n132), .out0(new_n138));
  aoi022aa1n03x5               g043(.a(new_n133), .b(new_n138), .c(new_n137), .d(new_n136), .o1(new_n139));
  xorb03aa1n02x5               g044(.a(new_n139), .b(\b[11] ), .c(new_n135), .out0(\s[12] ));
  nanp02aa1n02x5               g045(.a(new_n124), .b(new_n112), .o1(new_n141));
  nanp02aa1n02x5               g046(.a(new_n126), .b(new_n114), .o1(new_n142));
  tech160nm_fioaoi03aa1n03p5x5 g047(.a(new_n119), .b(new_n120), .c(new_n142), .o1(new_n143));
  xnrc02aa1n12x5               g048(.a(\b[11] ), .b(\a[12] ), .out0(new_n144));
  nano23aa1d15x5               g049(.a(new_n97), .b(new_n100), .c(new_n128), .d(new_n98), .out0(new_n145));
  nona22aa1d30x5               g050(.a(new_n145), .b(new_n144), .c(new_n132), .out0(new_n146));
  tech160nm_finand02aa1n05x5   g051(.a(new_n100), .b(new_n98), .o1(new_n147));
  oai122aa1n06x5               g052(.a(new_n147), .b(\b[9] ), .c(\a[10] ), .d(\b[10] ), .e(\a[11] ), .o1(new_n148));
  aoi022aa1n02x5               g053(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n149));
  aboi22aa1n09x5               g054(.a(\b[11] ), .b(new_n135), .c(new_n148), .d(new_n149), .out0(new_n150));
  aoai13aa1n03x5               g055(.a(new_n150), .b(new_n146), .c(new_n141), .d(new_n143), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d28x5               g057(.a(\a[13] ), .o1(new_n153));
  inv040aa1d32x5               g058(.a(\b[12] ), .o1(new_n154));
  oaoi03aa1n02x5               g059(.a(new_n153), .b(new_n154), .c(new_n151), .o1(new_n155));
  xnrb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv020aa1n03x5               g061(.a(new_n105), .o1(new_n157));
  nano23aa1n03x5               g062(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n158));
  aobi12aa1n03x7               g063(.a(new_n111), .b(new_n158), .c(new_n157), .out0(new_n159));
  nanp02aa1n02x5               g064(.a(new_n114), .b(new_n115), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n118), .b(new_n117), .out0(new_n161));
  xorc02aa1n02x5               g066(.a(\a[8] ), .b(\b[7] ), .out0(new_n162));
  nona23aa1n02x4               g067(.a(new_n116), .b(new_n162), .c(new_n161), .d(new_n160), .out0(new_n163));
  oai012aa1n04x7               g068(.a(new_n143), .b(new_n159), .c(new_n163), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n146), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(new_n148), .b(new_n149), .o1(new_n166));
  oaib12aa1n02x5               g071(.a(new_n166), .b(\b[11] ), .c(new_n135), .out0(new_n167));
  norp02aa1n02x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  nand42aa1n02x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nor002aa1d32x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand42aa1n20x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nano23aa1n06x5               g076(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n167), .c(new_n164), .d(new_n165), .o1(new_n173));
  aoai13aa1n12x5               g078(.a(new_n171), .b(new_n170), .c(new_n153), .d(new_n154), .o1(new_n174));
  nor042aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nand42aa1n04x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n173), .c(new_n174), .out0(\s[15] ));
  nor002aa1d32x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanp02aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n03x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  inv000aa1n02x5               g086(.a(new_n175), .o1(new_n182));
  inv000aa1n02x5               g087(.a(new_n176), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n173), .d(new_n174), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n184), .b(new_n181), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n174), .o1(new_n186));
  aoai13aa1n02x5               g091(.a(new_n177), .b(new_n186), .c(new_n151), .d(new_n172), .o1(new_n187));
  nona22aa1n02x4               g092(.a(new_n187), .b(new_n181), .c(new_n175), .out0(new_n188));
  nanp02aa1n02x5               g093(.a(new_n185), .b(new_n188), .o1(\s[16] ));
  nona32aa1n09x5               g094(.a(new_n172), .b(new_n181), .c(new_n183), .d(new_n175), .out0(new_n190));
  nor042aa1n09x5               g095(.a(new_n190), .b(new_n146), .o1(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n127), .c(new_n124), .d(new_n112), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n179), .o1(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n183), .c(new_n174), .d(new_n182), .o1(new_n194));
  nanp02aa1n06x5               g099(.a(new_n194), .b(new_n180), .o1(new_n195));
  oai012aa1n12x5               g100(.a(new_n195), .b(new_n150), .c(new_n190), .o1(new_n196));
  inv040aa1n09x5               g101(.a(new_n196), .o1(new_n197));
  nor002aa1n16x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  nand42aa1d28x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n200), .b(new_n197), .c(new_n192), .out0(\s[17] ));
  nanp02aa1n12x5               g106(.a(new_n197), .b(new_n192), .o1(new_n202));
  tech160nm_fiaoi012aa1n05x5   g107(.a(new_n198), .b(new_n202), .c(new_n200), .o1(new_n203));
  xnrb03aa1n03x5               g108(.a(new_n203), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor042aa1n06x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nand42aa1d28x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nano23aa1d15x5               g111(.a(new_n198), .b(new_n205), .c(new_n206), .d(new_n199), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n196), .c(new_n164), .d(new_n191), .o1(new_n208));
  oa0012aa1n02x5               g113(.a(new_n206), .b(new_n205), .c(new_n198), .o(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor042aa1n06x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand02aa1n06x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n12x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n208), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g120(.a(new_n208), .b(new_n210), .o1(new_n216));
  nor042aa1n06x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1d06x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n06x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n211), .c(new_n216), .d(new_n212), .o1(new_n220));
  aoai13aa1n06x5               g125(.a(new_n213), .b(new_n209), .c(new_n202), .d(new_n207), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n219), .c(new_n211), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n220), .b(new_n222), .o1(\s[20] ));
  nanb03aa1d18x5               g128(.a(new_n219), .b(new_n207), .c(new_n213), .out0(new_n224));
  nanb03aa1n09x5               g129(.a(new_n217), .b(new_n218), .c(new_n212), .out0(new_n225));
  orn002aa1n02x5               g130(.a(\a[19] ), .b(\b[18] ), .o(new_n226));
  oai112aa1n06x5               g131(.a(new_n226), .b(new_n206), .c(new_n205), .d(new_n198), .o1(new_n227));
  aoi012aa1n06x5               g132(.a(new_n217), .b(new_n211), .c(new_n218), .o1(new_n228));
  oai012aa1d24x5               g133(.a(new_n228), .b(new_n227), .c(new_n225), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n04x5               g135(.a(new_n230), .b(new_n224), .c(new_n197), .d(new_n192), .o1(new_n231));
  nor042aa1n04x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n224), .o1(new_n235));
  aoi112aa1n03x4               g140(.a(new_n234), .b(new_n229), .c(new_n202), .d(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n231), .c(new_n234), .o1(\s[21] ));
  nor042aa1n02x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nand42aa1n02x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nanb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n232), .c(new_n231), .d(new_n234), .o1(new_n241));
  nand02aa1n02x5               g146(.a(new_n231), .b(new_n234), .o1(new_n242));
  nona22aa1n02x5               g147(.a(new_n242), .b(new_n240), .c(new_n232), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n243), .b(new_n241), .o1(\s[22] ));
  nano23aa1n06x5               g149(.a(new_n232), .b(new_n238), .c(new_n239), .d(new_n233), .out0(new_n245));
  nanb02aa1n03x5               g150(.a(new_n224), .b(new_n245), .out0(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(new_n197), .c(new_n192), .o1(new_n247));
  oa0012aa1n02x5               g152(.a(new_n239), .b(new_n238), .c(new_n232), .o(new_n248));
  aoi012aa1n02x5               g153(.a(new_n248), .b(new_n229), .c(new_n245), .o1(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n246), .c(new_n197), .d(new_n192), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  aoi112aa1n02x5               g156(.a(new_n251), .b(new_n248), .c(new_n229), .d(new_n245), .o1(new_n252));
  aboi22aa1n03x5               g157(.a(new_n247), .b(new_n252), .c(new_n250), .d(new_n251), .out0(\s[23] ));
  norp02aa1n02x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[23] ), .b(\a[24] ), .out0(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n254), .c(new_n250), .d(new_n251), .o1(new_n256));
  nand02aa1n02x5               g161(.a(new_n250), .b(new_n251), .o1(new_n257));
  nona22aa1n02x5               g162(.a(new_n257), .b(new_n255), .c(new_n254), .out0(new_n258));
  nanp02aa1n03x5               g163(.a(new_n258), .b(new_n256), .o1(\s[24] ));
  norb02aa1n03x5               g164(.a(new_n251), .b(new_n255), .out0(new_n260));
  nano22aa1n03x7               g165(.a(new_n224), .b(new_n260), .c(new_n245), .out0(new_n261));
  aoai13aa1n02x5               g166(.a(new_n261), .b(new_n196), .c(new_n164), .d(new_n191), .o1(new_n262));
  nano22aa1n02x4               g167(.a(new_n217), .b(new_n212), .c(new_n218), .out0(new_n263));
  oai012aa1n02x5               g168(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .o1(new_n264));
  oab012aa1n02x4               g169(.a(new_n264), .b(new_n198), .c(new_n205), .out0(new_n265));
  inv020aa1n04x5               g170(.a(new_n228), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n245), .b(new_n266), .c(new_n265), .d(new_n263), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n248), .o1(new_n268));
  inv040aa1n02x5               g173(.a(new_n260), .o1(new_n269));
  oai022aa1n02x5               g174(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n270));
  aob012aa1n02x5               g175(.a(new_n270), .b(\b[23] ), .c(\a[24] ), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n268), .o1(new_n272));
  nanb02aa1n03x5               g177(.a(new_n272), .b(new_n262), .out0(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  tech160nm_fixnrc02aa1n04x5   g181(.a(\b[25] ), .b(\a[26] ), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .d(new_n276), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n276), .b(new_n272), .c(new_n202), .d(new_n261), .o1(new_n279));
  nona22aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n278), .b(new_n280), .o1(\s[26] ));
  norb02aa1n06x5               g186(.a(new_n276), .b(new_n277), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  nano23aa1d15x5               g188(.a(new_n283), .b(new_n224), .c(new_n260), .d(new_n245), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n196), .c(new_n164), .d(new_n191), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(\b[25] ), .b(\a[26] ), .o1(new_n286));
  oai022aa1n02x5               g191(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n287));
  aoi022aa1n06x5               g192(.a(new_n272), .b(new_n282), .c(new_n286), .d(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  xnbna2aa1n03x5               g194(.a(new_n289), .b(new_n288), .c(new_n285), .out0(\s[27] ));
  nand42aa1n02x5               g195(.a(new_n288), .b(new_n285), .o1(new_n291));
  norp02aa1n02x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  norp02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .o1(new_n293));
  nand42aa1n03x5               g198(.a(\b[27] ), .b(\a[28] ), .o1(new_n294));
  nanb02aa1n06x5               g199(.a(new_n293), .b(new_n294), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n292), .c(new_n291), .d(new_n289), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n260), .b(new_n248), .c(new_n229), .d(new_n245), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(new_n287), .b(new_n286), .o1(new_n298));
  aoai13aa1n04x5               g203(.a(new_n298), .b(new_n283), .c(new_n297), .d(new_n271), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n289), .b(new_n299), .c(new_n202), .d(new_n284), .o1(new_n300));
  nona22aa1n02x5               g205(.a(new_n300), .b(new_n295), .c(new_n292), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n296), .b(new_n301), .o1(\s[28] ));
  norb02aa1n15x5               g207(.a(new_n289), .b(new_n295), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n299), .c(new_n202), .d(new_n284), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .out0(new_n305));
  aoi012aa1n02x5               g210(.a(new_n293), .b(new_n292), .c(new_n294), .o1(new_n306));
  norb02aa1n02x5               g211(.a(new_n306), .b(new_n305), .out0(new_n307));
  inv000aa1d42x5               g212(.a(new_n303), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n306), .b(new_n308), .c(new_n288), .d(new_n285), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n304), .d(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g215(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g216(.a(new_n295), .b(new_n289), .c(new_n305), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n299), .c(new_n202), .d(new_n284), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  oao003aa1n02x5               g219(.a(\a[29] ), .b(\b[28] ), .c(new_n306), .carry(new_n315));
  norb02aa1n02x5               g220(.a(new_n315), .b(new_n314), .out0(new_n316));
  inv000aa1d42x5               g221(.a(new_n312), .o1(new_n317));
  aoai13aa1n02x7               g222(.a(new_n315), .b(new_n317), .c(new_n288), .d(new_n285), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n313), .d(new_n316), .o1(\s[30] ));
  nanp03aa1n02x5               g224(.a(new_n303), .b(new_n305), .c(new_n314), .o1(new_n320));
  nanb02aa1n02x5               g225(.a(new_n320), .b(new_n291), .out0(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n323), .b(new_n320), .c(new_n288), .d(new_n285), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n321), .b(new_n324), .c(new_n325), .d(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g231(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g232(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  nanp02aa1n02x5               g234(.a(new_n158), .b(new_n157), .o1(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n116), .b(new_n330), .c(new_n111), .out0(\s[5] ));
  oaoi03aa1n02x5               g236(.a(\a[5] ), .b(\b[4] ), .c(new_n159), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fioai012aa1n05x5   g238(.a(new_n117), .b(new_n332), .c(new_n118), .o1(new_n334));
  xnbna2aa1n03x5               g239(.a(new_n334), .b(new_n114), .c(new_n115), .out0(\s[7] ));
  oaoi03aa1n03x5               g240(.a(\a[7] ), .b(\b[6] ), .c(new_n334), .o1(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g242(.a(new_n129), .b(new_n141), .c(new_n143), .out0(\s[9] ));
endmodule


