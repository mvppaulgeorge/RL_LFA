// Benchmark "adder" written by ABC on Thu Jul 18 09:35:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n305, new_n306, new_n308, new_n311, new_n313,
    new_n314, new_n316, new_n317, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n16x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand22aa1n09x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n06x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nand42aa1n04x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor022aa1n16x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  oa0022aa1n06x5               g008(.a(\a[8] ), .b(\b[7] ), .c(\a[7] ), .d(\b[6] ), .o(new_n104));
  nor042aa1n12x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  norp02aa1n12x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nand02aa1d28x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nona23aa1n02x5               g013(.a(new_n108), .b(new_n106), .c(new_n105), .d(new_n107), .out0(new_n109));
  nano32aa1n03x7               g014(.a(new_n109), .b(new_n104), .c(new_n103), .d(new_n102), .out0(new_n110));
  and002aa1n06x5               g015(.a(\b[3] ), .b(\a[4] ), .o(new_n111));
  inv000aa1d42x5               g016(.a(new_n111), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  oab012aa1n02x5               g018(.a(new_n113), .b(\a[4] ), .c(\b[3] ), .out0(new_n114));
  nand02aa1d12x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nand42aa1n06x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nanb03aa1d18x5               g021(.a(new_n113), .b(new_n116), .c(new_n115), .out0(new_n117));
  nand02aa1d06x5               g022(.a(\b[0] ), .b(\a[1] ), .o1(new_n118));
  nor042aa1n03x5               g023(.a(\b[1] ), .b(\a[2] ), .o1(new_n119));
  norb03aa1n12x5               g024(.a(new_n115), .b(new_n119), .c(new_n118), .out0(new_n120));
  oai012aa1n04x7               g025(.a(new_n114), .b(new_n120), .c(new_n117), .o1(new_n121));
  nanp03aa1d12x5               g026(.a(new_n110), .b(new_n121), .c(new_n112), .o1(new_n122));
  aoai13aa1n12x5               g027(.a(new_n102), .b(new_n107), .c(new_n105), .d(new_n108), .o1(new_n123));
  aoi022aa1d18x5               g028(.a(new_n123), .b(new_n104), .c(\a[8] ), .d(\b[7] ), .o1(new_n124));
  nona22aa1n09x5               g029(.a(new_n122), .b(new_n124), .c(new_n101), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n99), .b(new_n125), .c(new_n100), .out0(\s[10] ));
  nor002aa1d32x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  nand42aa1n08x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  aoai13aa1n06x5               g034(.a(new_n98), .b(new_n97), .c(new_n125), .d(new_n100), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n128), .c(new_n129), .out0(\s[11] ));
  nanb02aa1n02x5               g036(.a(new_n127), .b(new_n129), .out0(new_n132));
  nor022aa1n12x5               g037(.a(\b[11] ), .b(\a[12] ), .o1(new_n133));
  nand42aa1n10x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  oaoi13aa1n02x7               g040(.a(new_n135), .b(new_n128), .c(new_n130), .d(new_n132), .o1(new_n136));
  oai112aa1n02x7               g041(.a(new_n128), .b(new_n135), .c(new_n130), .d(new_n132), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(\s[12] ));
  inv000aa1d42x5               g043(.a(new_n124), .o1(new_n139));
  nano23aa1n06x5               g044(.a(new_n127), .b(new_n133), .c(new_n134), .d(new_n129), .out0(new_n140));
  nanb02aa1n03x5               g045(.a(new_n101), .b(new_n100), .out0(new_n141));
  nona22aa1n09x5               g046(.a(new_n140), .b(new_n141), .c(new_n99), .out0(new_n142));
  nona23aa1n12x5               g047(.a(new_n134), .b(new_n129), .c(new_n127), .d(new_n133), .out0(new_n143));
  aoi012aa1n06x5               g048(.a(new_n97), .b(new_n101), .c(new_n98), .o1(new_n144));
  aoi012aa1n06x5               g049(.a(new_n133), .b(new_n127), .c(new_n134), .o1(new_n145));
  oai012aa1d24x5               g050(.a(new_n145), .b(new_n143), .c(new_n144), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  aoai13aa1n06x5               g052(.a(new_n147), .b(new_n142), .c(new_n122), .d(new_n139), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g054(.a(\a[14] ), .o1(new_n150));
  nor002aa1n02x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[12] ), .b(\a[13] ), .out0(new_n152));
  inv040aa1n02x5               g057(.a(new_n152), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n151), .b(new_n148), .c(new_n153), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(new_n150), .out0(\s[14] ));
  tech160nm_fixorc02aa1n03p5x5 g060(.a(\a[14] ), .b(\b[13] ), .out0(new_n156));
  norb02aa1n06x4               g061(.a(new_n156), .b(new_n152), .out0(new_n157));
  inv000aa1d42x5               g062(.a(\b[13] ), .o1(new_n158));
  oao003aa1n02x5               g063(.a(new_n150), .b(new_n158), .c(new_n151), .carry(new_n159));
  nor042aa1n04x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nand42aa1d28x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n159), .c(new_n148), .d(new_n157), .o1(new_n163));
  aoi112aa1n02x5               g068(.a(new_n162), .b(new_n159), .c(new_n148), .d(new_n157), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(\s[15] ));
  nor042aa1n04x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand42aa1n16x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  nona22aa1n02x5               g073(.a(new_n163), .b(new_n168), .c(new_n160), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n168), .o1(new_n170));
  oaoi13aa1n06x5               g075(.a(new_n170), .b(new_n163), .c(\a[15] ), .d(\b[14] ), .o1(new_n171));
  norb02aa1n03x4               g076(.a(new_n169), .b(new_n171), .out0(\s[16] ));
  oaoi13aa1n09x5               g077(.a(new_n111), .b(new_n114), .c(new_n120), .d(new_n117), .o1(new_n173));
  nano23aa1d15x5               g078(.a(new_n160), .b(new_n166), .c(new_n167), .d(new_n161), .out0(new_n174));
  nano32aa1n03x7               g079(.a(new_n142), .b(new_n174), .c(new_n153), .d(new_n156), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n124), .c(new_n173), .d(new_n110), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n166), .b(new_n160), .c(new_n167), .o1(new_n177));
  aob012aa1n06x5               g082(.a(new_n177), .b(new_n174), .c(new_n159), .out0(new_n178));
  aoi013aa1n09x5               g083(.a(new_n178), .b(new_n146), .c(new_n157), .d(new_n174), .o1(new_n179));
  nanp02aa1n06x5               g084(.a(new_n176), .b(new_n179), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g086(.a(\a[18] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(new_n183), .b(new_n184), .c(new_n180), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n182), .out0(\s[18] ));
  xroi22aa1d06x4               g091(.a(new_n183), .b(\b[16] ), .c(new_n182), .d(\b[17] ), .out0(new_n187));
  nand02aa1d04x5               g092(.a(\b[17] ), .b(\a[18] ), .o1(new_n188));
  nona22aa1n02x4               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(new_n189));
  oaib12aa1n09x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n182), .out0(new_n190));
  nor022aa1n16x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nand42aa1n02x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  norb02aa1n02x5               g097(.a(new_n192), .b(new_n191), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n190), .c(new_n180), .d(new_n187), .o1(new_n194));
  aoi112aa1n02x5               g099(.a(new_n193), .b(new_n190), .c(new_n180), .d(new_n187), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n194), .b(new_n195), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n04x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nanp02aa1n04x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  nona22aa1n02x5               g105(.a(new_n194), .b(new_n200), .c(new_n191), .out0(new_n201));
  orn002aa1n02x5               g106(.a(\a[19] ), .b(\b[18] ), .o(new_n202));
  aobi12aa1n06x5               g107(.a(new_n200), .b(new_n194), .c(new_n202), .out0(new_n203));
  norb02aa1n03x4               g108(.a(new_n201), .b(new_n203), .out0(\s[20] ));
  nano23aa1n06x5               g109(.a(new_n191), .b(new_n198), .c(new_n199), .d(new_n192), .out0(new_n205));
  nanp02aa1n02x5               g110(.a(new_n187), .b(new_n205), .o1(new_n206));
  norp02aa1n02x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  aoi013aa1n06x4               g112(.a(new_n207), .b(new_n188), .c(new_n183), .d(new_n184), .o1(new_n208));
  nona23aa1n09x5               g113(.a(new_n199), .b(new_n192), .c(new_n191), .d(new_n198), .out0(new_n209));
  aoi012aa1n06x5               g114(.a(new_n198), .b(new_n191), .c(new_n199), .o1(new_n210));
  oai012aa1n18x5               g115(.a(new_n210), .b(new_n209), .c(new_n208), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n206), .c(new_n176), .d(new_n179), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n06x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  nanp02aa1n02x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  nor042aa1n02x5               g122(.a(\b[21] ), .b(\a[22] ), .o1(new_n218));
  nanp02aa1n04x5               g123(.a(\b[21] ), .b(\a[22] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  aoi112aa1n02x5               g125(.a(new_n215), .b(new_n220), .c(new_n213), .d(new_n217), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n220), .b(new_n215), .c(new_n213), .d(new_n217), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n222), .b(new_n221), .out0(\s[22] ));
  nano23aa1n06x5               g128(.a(new_n215), .b(new_n218), .c(new_n219), .d(new_n216), .out0(new_n224));
  nanp03aa1n02x5               g129(.a(new_n187), .b(new_n205), .c(new_n224), .o1(new_n225));
  aoi012aa1n12x5               g130(.a(new_n218), .b(new_n215), .c(new_n219), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoi012aa1n02x5               g132(.a(new_n227), .b(new_n211), .c(new_n224), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n225), .c(new_n176), .d(new_n179), .o1(new_n229));
  xorb03aa1n02x5               g134(.a(new_n229), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g135(.a(\b[22] ), .b(\a[23] ), .o1(new_n231));
  tech160nm_fixorc02aa1n02p5x5 g136(.a(\a[23] ), .b(\b[22] ), .out0(new_n232));
  tech160nm_fixorc02aa1n05x5   g137(.a(\a[24] ), .b(\b[23] ), .out0(new_n233));
  aoi112aa1n02x5               g138(.a(new_n231), .b(new_n233), .c(new_n229), .d(new_n232), .o1(new_n234));
  aoai13aa1n03x5               g139(.a(new_n233), .b(new_n231), .c(new_n229), .d(new_n232), .o1(new_n235));
  norb02aa1n02x7               g140(.a(new_n235), .b(new_n234), .out0(\s[24] ));
  inv000aa1n06x5               g141(.a(new_n210), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n224), .b(new_n237), .c(new_n205), .d(new_n190), .o1(new_n238));
  and002aa1n18x5               g143(.a(new_n233), .b(new_n232), .o(new_n239));
  inv000aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n241));
  oab012aa1n02x4               g146(.a(new_n241), .b(\a[24] ), .c(\b[23] ), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n240), .c(new_n238), .d(new_n226), .o1(new_n243));
  nano32aa1n02x4               g148(.a(new_n206), .b(new_n233), .c(new_n224), .d(new_n232), .out0(new_n244));
  xorc02aa1n02x5               g149(.a(\a[25] ), .b(\b[24] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n243), .c(new_n180), .d(new_n244), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n243), .b(new_n245), .c(new_n180), .d(new_n244), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[26] ), .b(\b[25] ), .out0(new_n250));
  nona22aa1n03x5               g155(.a(new_n246), .b(new_n250), .c(new_n249), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n249), .o1(new_n252));
  aobi12aa1n06x5               g157(.a(new_n250), .b(new_n246), .c(new_n252), .out0(new_n253));
  norb02aa1n03x4               g158(.a(new_n251), .b(new_n253), .out0(\s[26] ));
  nand42aa1n03x5               g159(.a(new_n122), .b(new_n139), .o1(new_n255));
  nanp03aa1n02x5               g160(.a(new_n153), .b(new_n174), .c(new_n156), .o1(new_n256));
  oabi12aa1n02x5               g161(.a(new_n178), .b(new_n147), .c(new_n256), .out0(new_n257));
  inv000aa1d42x5               g162(.a(\a[25] ), .o1(new_n258));
  inv020aa1n04x5               g163(.a(\a[26] ), .o1(new_n259));
  xroi22aa1d06x4               g164(.a(new_n258), .b(\b[24] ), .c(new_n259), .d(\b[25] ), .out0(new_n260));
  nano22aa1n03x7               g165(.a(new_n225), .b(new_n239), .c(new_n260), .out0(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n257), .c(new_n255), .d(new_n175), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[26] ), .b(\b[25] ), .c(new_n252), .carry(new_n263));
  aobi12aa1n06x5               g168(.a(new_n263), .b(new_n243), .c(new_n260), .out0(new_n264));
  xorc02aa1n02x5               g169(.a(\a[27] ), .b(\b[26] ), .out0(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n264), .c(new_n262), .out0(\s[27] ));
  norp02aa1n02x5               g171(.a(\b[26] ), .b(\a[27] ), .o1(new_n267));
  inv040aa1n03x5               g172(.a(new_n267), .o1(new_n268));
  aobi12aa1n06x5               g173(.a(new_n265), .b(new_n264), .c(new_n262), .out0(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[27] ), .b(\a[28] ), .out0(new_n270));
  nano22aa1n03x5               g175(.a(new_n269), .b(new_n268), .c(new_n270), .out0(new_n271));
  inv020aa1n02x5               g176(.a(new_n261), .o1(new_n272));
  aoi012aa1n06x5               g177(.a(new_n272), .b(new_n176), .c(new_n179), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n239), .b(new_n227), .c(new_n211), .d(new_n224), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n260), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n263), .b(new_n275), .c(new_n274), .d(new_n242), .o1(new_n276));
  oaih12aa1n02x5               g181(.a(new_n265), .b(new_n276), .c(new_n273), .o1(new_n277));
  tech160nm_fiaoi012aa1n02p5x5 g182(.a(new_n270), .b(new_n277), .c(new_n268), .o1(new_n278));
  norp02aa1n03x5               g183(.a(new_n278), .b(new_n271), .o1(\s[28] ));
  xnrc02aa1n02x5               g184(.a(\b[28] ), .b(\a[29] ), .out0(new_n280));
  norb02aa1n02x5               g185(.a(new_n265), .b(new_n270), .out0(new_n281));
  aobi12aa1n02x7               g186(.a(new_n281), .b(new_n264), .c(new_n262), .out0(new_n282));
  oao003aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n268), .carry(new_n283));
  nano22aa1n03x5               g188(.a(new_n282), .b(new_n280), .c(new_n283), .out0(new_n284));
  oaih12aa1n02x5               g189(.a(new_n281), .b(new_n276), .c(new_n273), .o1(new_n285));
  tech160nm_fiaoi012aa1n02p5x5 g190(.a(new_n280), .b(new_n285), .c(new_n283), .o1(new_n286));
  norp02aa1n03x5               g191(.a(new_n286), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n118), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g193(.a(new_n265), .b(new_n280), .c(new_n270), .out0(new_n289));
  aobi12aa1n02x7               g194(.a(new_n289), .b(new_n264), .c(new_n262), .out0(new_n290));
  oao003aa1n02x5               g195(.a(\a[29] ), .b(\b[28] ), .c(new_n283), .carry(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[29] ), .b(\a[30] ), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n290), .b(new_n291), .c(new_n292), .out0(new_n293));
  oaih12aa1n02x5               g198(.a(new_n289), .b(new_n276), .c(new_n273), .o1(new_n294));
  tech160nm_fiaoi012aa1n02p5x5 g199(.a(new_n292), .b(new_n294), .c(new_n291), .o1(new_n295));
  norp02aa1n03x5               g200(.a(new_n295), .b(new_n293), .o1(\s[30] ));
  norb02aa1n02x5               g201(.a(new_n289), .b(new_n292), .out0(new_n297));
  aobi12aa1n02x7               g202(.a(new_n297), .b(new_n264), .c(new_n262), .out0(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n291), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n300), .out0(new_n301));
  oaih12aa1n02x5               g206(.a(new_n297), .b(new_n276), .c(new_n273), .o1(new_n302));
  aoi012aa1n03x5               g207(.a(new_n300), .b(new_n302), .c(new_n299), .o1(new_n303));
  norp02aa1n03x5               g208(.a(new_n303), .b(new_n301), .o1(\s[31] ));
  norb02aa1n02x5               g209(.a(new_n116), .b(new_n113), .out0(new_n305));
  oaoi13aa1n02x5               g210(.a(new_n305), .b(new_n115), .c(new_n119), .d(new_n118), .o1(new_n306));
  oab012aa1n02x4               g211(.a(new_n306), .b(new_n117), .c(new_n120), .out0(\s[3] ));
  oabi12aa1n02x5               g212(.a(new_n113), .b(new_n120), .c(new_n117), .out0(new_n308));
  xorb03aa1n02x5               g213(.a(new_n308), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g214(.a(new_n173), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi013aa1n02x4               g215(.a(new_n105), .b(new_n121), .c(new_n112), .d(new_n106), .o1(new_n311));
  xnrb03aa1n02x5               g216(.a(new_n311), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb03aa1n02x5               g217(.a(new_n107), .b(new_n311), .c(new_n108), .out0(new_n313));
  xorc02aa1n02x5               g218(.a(\a[7] ), .b(\b[6] ), .out0(new_n314));
  xobna2aa1n03x5               g219(.a(new_n314), .b(new_n313), .c(new_n108), .out0(\s[7] ));
  orn002aa1n02x5               g220(.a(\a[7] ), .b(\b[6] ), .o(new_n316));
  nanp03aa1n02x5               g221(.a(new_n313), .b(new_n108), .c(new_n314), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[8] ), .b(\b[7] ), .out0(new_n318));
  xnbna2aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n316), .out0(\s[8] ));
  xobna2aa1n03x5               g224(.a(new_n141), .b(new_n122), .c(new_n139), .out0(\s[9] ));
endmodule


