// Benchmark "adder" written by ABC on Thu Jul 18 06:30:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n352, new_n354, new_n355, new_n357, new_n359, new_n360, new_n361,
    new_n363, new_n364, new_n366, new_n368;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  orn002aa1n03x5               g002(.a(\a[2] ), .b(\b[1] ), .o(new_n98));
  nand22aa1n04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nand42aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  aob012aa1n03x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .out0(new_n101));
  nor042aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand02aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n03x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor042aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n06x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nanp03aa1n06x5               g012(.a(new_n101), .b(new_n104), .c(new_n107), .o1(new_n108));
  oaih12aa1n06x5               g013(.a(new_n103), .b(new_n105), .c(new_n102), .o1(new_n109));
  tech160nm_fixorc02aa1n02p5x5 g014(.a(\a[8] ), .b(\b[7] ), .out0(new_n110));
  nor042aa1d18x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n16x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  norb02aa1n06x4               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nand02aa1d08x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor042aa1n04x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor042aa1n04x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanp02aa1n04x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nano23aa1n03x7               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nand23aa1n03x5               g023(.a(new_n118), .b(new_n110), .c(new_n113), .o1(new_n119));
  nand42aa1n04x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nano22aa1n03x5               g025(.a(new_n111), .b(new_n120), .c(new_n112), .out0(new_n121));
  oai022aa1n03x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  oa0012aa1n03x5               g027(.a(new_n114), .b(\b[7] ), .c(\a[8] ), .o(new_n123));
  inv040aa1n03x5               g028(.a(new_n111), .o1(new_n124));
  oaoi03aa1n09x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n121), .c(new_n123), .d(new_n122), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n126), .b(new_n119), .c(new_n108), .d(new_n109), .o1(new_n127));
  xnrc02aa1n12x5               g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(new_n127), .b(new_n129), .o1(new_n130));
  tech160nm_fixorc02aa1n03p5x5 g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  nanp02aa1n02x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  oai022aa1d18x5               g037(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  nanb03aa1n02x5               g038(.a(new_n133), .b(new_n130), .c(new_n132), .out0(new_n134));
  aoai13aa1n02x5               g039(.a(new_n134), .b(new_n131), .c(new_n97), .d(new_n130), .o1(\s[10] ));
  norb02aa1n02x5               g040(.a(new_n131), .b(new_n128), .out0(new_n136));
  nand22aa1n03x5               g041(.a(new_n127), .b(new_n136), .o1(new_n137));
  nanp02aa1n06x5               g042(.a(new_n133), .b(new_n132), .o1(new_n138));
  xorc02aa1n12x5               g043(.a(\a[11] ), .b(\b[10] ), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n137), .c(new_n138), .out0(\s[11] ));
  aobi12aa1n02x5               g045(.a(new_n139), .b(new_n137), .c(new_n138), .out0(new_n141));
  orn002aa1n02x5               g046(.a(\a[11] ), .b(\b[10] ), .o(new_n142));
  and002aa1n02x5               g047(.a(\b[10] ), .b(\a[11] ), .o(new_n143));
  aoai13aa1n02x5               g048(.a(new_n142), .b(new_n143), .c(new_n137), .d(new_n138), .o1(new_n144));
  orn002aa1n24x5               g049(.a(\a[12] ), .b(\b[11] ), .o(new_n145));
  nanp02aa1n09x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand02aa1d08x5               g051(.a(new_n145), .b(new_n146), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  oai112aa1n02x5               g053(.a(new_n145), .b(new_n146), .c(\b[10] ), .d(\a[11] ), .o1(new_n149));
  obai22aa1n03x5               g054(.a(new_n144), .b(new_n148), .c(new_n141), .d(new_n149), .out0(\s[12] ));
  nanp02aa1n02x5               g055(.a(new_n108), .b(new_n109), .o1(new_n151));
  nona23aa1n02x4               g056(.a(new_n114), .b(new_n117), .c(new_n116), .d(new_n115), .out0(new_n152));
  nano22aa1n02x4               g057(.a(new_n152), .b(new_n110), .c(new_n113), .out0(new_n153));
  nanp02aa1n02x5               g058(.a(new_n151), .b(new_n153), .o1(new_n154));
  nona23aa1d18x5               g059(.a(new_n131), .b(new_n139), .c(new_n128), .d(new_n147), .out0(new_n155));
  aoai13aa1n06x5               g060(.a(new_n145), .b(new_n143), .c(new_n138), .d(new_n142), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(new_n156), .b(new_n146), .o1(new_n157));
  aoai13aa1n04x5               g062(.a(new_n157), .b(new_n155), .c(new_n154), .d(new_n126), .o1(new_n158));
  xorc02aa1n02x5               g063(.a(\a[13] ), .b(\b[12] ), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n155), .o1(new_n160));
  inv000aa1n02x5               g065(.a(new_n157), .o1(new_n161));
  aoi112aa1n02x5               g066(.a(new_n159), .b(new_n161), .c(new_n127), .d(new_n160), .o1(new_n162));
  aoi012aa1n02x5               g067(.a(new_n162), .b(new_n158), .c(new_n159), .o1(\s[13] ));
  inv040aa1d32x5               g068(.a(\a[13] ), .o1(new_n164));
  inv040aa1d32x5               g069(.a(\b[12] ), .o1(new_n165));
  nand42aa1n02x5               g070(.a(new_n165), .b(new_n164), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n159), .b(new_n161), .c(new_n127), .d(new_n160), .o1(new_n167));
  nor002aa1d32x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand42aa1d28x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  nano22aa1n02x4               g075(.a(new_n168), .b(new_n166), .c(new_n169), .out0(new_n171));
  nanp02aa1n02x5               g076(.a(new_n167), .b(new_n171), .o1(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n170), .c(new_n166), .d(new_n167), .o1(\s[14] ));
  nand42aa1n03x5               g078(.a(\b[12] ), .b(\a[13] ), .o1(new_n174));
  nano32aa1n02x5               g079(.a(new_n168), .b(new_n166), .c(new_n169), .d(new_n174), .out0(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n161), .c(new_n127), .d(new_n160), .o1(new_n176));
  aoai13aa1n12x5               g081(.a(new_n169), .b(new_n168), .c(new_n164), .d(new_n165), .o1(new_n177));
  nor002aa1n12x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nand02aa1d24x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  norb02aa1n09x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n176), .c(new_n177), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(new_n178), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n177), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n180), .b(new_n183), .c(new_n158), .d(new_n175), .o1(new_n184));
  nor002aa1n10x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nand02aa1n06x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  norb02aa1n02x5               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n180), .o1(new_n188));
  norb03aa1n02x5               g093(.a(new_n186), .b(new_n178), .c(new_n185), .out0(new_n189));
  aoai13aa1n02x5               g094(.a(new_n189), .b(new_n188), .c(new_n176), .d(new_n177), .o1(new_n190));
  aoai13aa1n02x5               g095(.a(new_n190), .b(new_n187), .c(new_n184), .d(new_n182), .o1(\s[16] ));
  nano32aa1d12x5               g096(.a(new_n155), .b(new_n187), .c(new_n175), .d(new_n180), .out0(new_n192));
  nanp02aa1n06x5               g097(.a(new_n127), .b(new_n192), .o1(new_n193));
  aoi012aa1n02x5               g098(.a(new_n185), .b(\a[15] ), .c(\b[14] ), .o1(new_n194));
  aoi022aa1n02x5               g099(.a(new_n165), .b(new_n164), .c(\a[12] ), .d(\b[11] ), .o1(new_n195));
  nona23aa1n02x4               g100(.a(new_n169), .b(new_n174), .c(new_n178), .d(new_n168), .out0(new_n196));
  nano32aa1n03x7               g101(.a(new_n196), .b(new_n195), .c(new_n194), .d(new_n186), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n179), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n185), .o1(new_n199));
  aoai13aa1n02x5               g104(.a(new_n199), .b(new_n198), .c(new_n177), .d(new_n182), .o1(new_n200));
  aoi022aa1n06x5               g105(.a(new_n156), .b(new_n197), .c(new_n200), .d(new_n186), .o1(new_n201));
  nanp02aa1n09x5               g106(.a(new_n193), .b(new_n201), .o1(new_n202));
  xorc02aa1n12x5               g107(.a(\a[17] ), .b(\b[16] ), .out0(new_n203));
  aoi122aa1n02x5               g108(.a(new_n203), .b(new_n200), .c(new_n186), .d(new_n156), .e(new_n197), .o1(new_n204));
  aoi022aa1n02x5               g109(.a(new_n202), .b(new_n203), .c(new_n193), .d(new_n204), .o1(\s[17] ));
  nor042aa1n03x5               g110(.a(\b[16] ), .b(\a[17] ), .o1(new_n206));
  inv040aa1n03x5               g111(.a(new_n206), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n186), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(new_n156), .b(new_n197), .o1(new_n209));
  inv000aa1d42x5               g114(.a(\a[16] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(\b[15] ), .o1(new_n211));
  nand22aa1n03x5               g116(.a(new_n177), .b(new_n182), .o1(new_n212));
  aoi022aa1n06x5               g117(.a(new_n212), .b(new_n179), .c(new_n210), .d(new_n211), .o1(new_n213));
  oai012aa1n12x5               g118(.a(new_n209), .b(new_n213), .c(new_n208), .o1(new_n214));
  aoai13aa1n02x5               g119(.a(new_n203), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n215));
  xorc02aa1n12x5               g120(.a(\a[18] ), .b(\b[17] ), .out0(new_n216));
  oai022aa1d24x5               g121(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(\a[18] ), .c(\b[17] ), .o1(new_n218));
  nanp02aa1n02x5               g123(.a(new_n215), .b(new_n218), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n216), .c(new_n207), .d(new_n215), .o1(\s[18] ));
  and002aa1n02x5               g125(.a(new_n216), .b(new_n203), .o(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n222));
  oaoi03aa1n02x5               g127(.a(\a[18] ), .b(\b[17] ), .c(new_n207), .o1(new_n223));
  inv000aa1n02x5               g128(.a(new_n223), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[19] ), .b(\b[18] ), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n222), .c(new_n224), .out0(\s[19] ));
  xnrc02aa1n02x5               g131(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g132(.a(\a[19] ), .o1(new_n228));
  nanb02aa1n02x5               g133(.a(\b[18] ), .b(new_n228), .out0(new_n229));
  aoai13aa1n06x5               g134(.a(new_n225), .b(new_n223), .c(new_n202), .d(new_n221), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[20] ), .b(\b[19] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n225), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(\b[19] ), .b(\a[20] ), .o1(new_n233));
  oai022aa1d18x5               g138(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n233), .b(new_n234), .out0(new_n235));
  aoai13aa1n02x5               g140(.a(new_n235), .b(new_n232), .c(new_n222), .d(new_n224), .o1(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n231), .c(new_n230), .d(new_n229), .o1(\s[20] ));
  inv040aa1d32x5               g142(.a(\a[20] ), .o1(new_n238));
  xroi22aa1d06x4               g143(.a(new_n228), .b(\b[18] ), .c(new_n238), .d(\b[19] ), .out0(new_n239));
  nand23aa1n04x5               g144(.a(new_n239), .b(new_n203), .c(new_n216), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n242));
  aoi022aa1n12x5               g147(.a(\b[18] ), .b(\a[19] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n243));
  aoi012aa1n12x5               g148(.a(new_n234), .b(new_n217), .c(new_n243), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n233), .b(new_n244), .out0(new_n245));
  inv000aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  xorc02aa1n12x5               g151(.a(\a[21] ), .b(\b[20] ), .out0(new_n247));
  xnbna2aa1n03x5               g152(.a(new_n247), .b(new_n242), .c(new_n246), .out0(\s[21] ));
  nor002aa1d24x5               g153(.a(\b[20] ), .b(\a[21] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n03x5               g155(.a(new_n247), .b(new_n245), .c(new_n202), .d(new_n241), .o1(new_n251));
  nor022aa1n16x5               g156(.a(\b[21] ), .b(\a[22] ), .o1(new_n252));
  nanp02aa1n04x5               g157(.a(\b[21] ), .b(\a[22] ), .o1(new_n253));
  norb02aa1n03x5               g158(.a(new_n253), .b(new_n252), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n247), .o1(new_n255));
  norb03aa1n02x5               g160(.a(new_n253), .b(new_n249), .c(new_n252), .out0(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n255), .c(new_n242), .d(new_n246), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n254), .c(new_n251), .d(new_n250), .o1(\s[22] ));
  and002aa1n02x5               g163(.a(new_n247), .b(new_n254), .o(new_n259));
  norb02aa1n02x5               g164(.a(new_n259), .b(new_n240), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n261));
  tech160nm_fiaoi012aa1n04x5   g166(.a(new_n249), .b(\a[20] ), .c(\b[19] ), .o1(new_n262));
  tech160nm_fiaoi012aa1n04x5   g167(.a(new_n252), .b(\a[21] ), .c(\b[20] ), .o1(new_n263));
  nand23aa1n03x5               g168(.a(new_n262), .b(new_n263), .c(new_n253), .o1(new_n264));
  inv000aa1d42x5               g169(.a(\a[21] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(\b[20] ), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n253), .b(new_n252), .c(new_n265), .d(new_n266), .o1(new_n267));
  oai012aa1n12x5               g172(.a(new_n267), .b(new_n264), .c(new_n244), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[23] ), .b(\b[22] ), .out0(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoi012aa1n03x5               g176(.a(new_n271), .b(new_n261), .c(new_n269), .o1(new_n272));
  oai112aa1n02x5               g177(.a(new_n267), .b(new_n271), .c(new_n264), .d(new_n244), .o1(new_n273));
  aoib12aa1n02x7               g178(.a(new_n272), .b(new_n261), .c(new_n273), .out0(\s[23] ));
  nor042aa1n06x5               g179(.a(\b[22] ), .b(\a[23] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n270), .b(new_n268), .c(new_n202), .d(new_n260), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .out0(new_n278));
  oai022aa1n02x5               g183(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n279));
  aoi012aa1n02x5               g184(.a(new_n279), .b(\a[24] ), .c(\b[23] ), .o1(new_n280));
  aoai13aa1n02x7               g185(.a(new_n280), .b(new_n271), .c(new_n261), .d(new_n269), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n278), .c(new_n277), .d(new_n276), .o1(\s[24] ));
  nanp02aa1n02x5               g187(.a(\b[22] ), .b(\a[23] ), .o1(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[23] ), .b(\a[24] ), .out0(new_n284));
  nano22aa1n02x4               g189(.a(new_n284), .b(new_n276), .c(new_n283), .out0(new_n285));
  nano22aa1n02x5               g190(.a(new_n240), .b(new_n259), .c(new_n285), .out0(new_n286));
  oaoi03aa1n02x5               g191(.a(\a[24] ), .b(\b[23] ), .c(new_n276), .o1(new_n287));
  aoi012aa1n02x5               g192(.a(new_n287), .b(new_n268), .c(new_n285), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[25] ), .b(\b[24] ), .out0(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n289), .c(new_n202), .d(new_n286), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n286), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n292));
  nanp02aa1n02x5               g197(.a(new_n278), .b(new_n270), .o1(new_n293));
  oaoi13aa1n06x5               g198(.a(new_n293), .b(new_n267), .c(new_n264), .d(new_n244), .o1(new_n294));
  nona32aa1n02x4               g199(.a(new_n292), .b(new_n290), .c(new_n294), .d(new_n287), .out0(new_n295));
  and002aa1n03x5               g200(.a(new_n291), .b(new_n295), .o(\s[25] ));
  nor042aa1n03x5               g201(.a(\b[24] ), .b(\a[25] ), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n297), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[26] ), .b(\b[25] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n290), .o1(new_n300));
  oai022aa1n02x5               g205(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n301));
  aoi012aa1n02x5               g206(.a(new_n301), .b(\a[26] ), .c(\b[25] ), .o1(new_n302));
  aoai13aa1n04x5               g207(.a(new_n302), .b(new_n300), .c(new_n292), .d(new_n288), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n299), .c(new_n291), .d(new_n298), .o1(\s[26] ));
  and002aa1n02x5               g209(.a(new_n299), .b(new_n290), .o(new_n305));
  nano32aa1n03x7               g210(.a(new_n240), .b(new_n305), .c(new_n259), .d(new_n285), .out0(new_n306));
  aoai13aa1n12x5               g211(.a(new_n306), .b(new_n214), .c(new_n127), .d(new_n192), .o1(new_n307));
  oaoi03aa1n02x5               g212(.a(\a[26] ), .b(\b[25] ), .c(new_n298), .o1(new_n308));
  oaoi13aa1n04x5               g213(.a(new_n308), .b(new_n305), .c(new_n294), .d(new_n287), .o1(new_n309));
  nanp02aa1n09x5               g214(.a(new_n307), .b(new_n309), .o1(new_n310));
  xorc02aa1n12x5               g215(.a(\a[27] ), .b(\b[26] ), .out0(new_n311));
  aoi112aa1n02x5               g216(.a(new_n311), .b(new_n308), .c(new_n289), .d(new_n305), .o1(new_n312));
  aoi022aa1n02x5               g217(.a(new_n312), .b(new_n307), .c(new_n310), .d(new_n311), .o1(\s[27] ));
  norp02aa1n02x5               g218(.a(\b[26] ), .b(\a[27] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  nanp02aa1n03x5               g220(.a(new_n310), .b(new_n311), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[28] ), .b(\b[27] ), .out0(new_n317));
  inv000aa1d42x5               g222(.a(new_n311), .o1(new_n318));
  oai022aa1n02x5               g223(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n319), .b(\a[28] ), .c(\b[27] ), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n318), .c(new_n307), .d(new_n309), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n316), .d(new_n315), .o1(\s[28] ));
  xnrc02aa1n02x5               g227(.a(\b[28] ), .b(\a[29] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(new_n317), .b(new_n311), .o(new_n324));
  inv000aa1d42x5               g229(.a(new_n324), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[27] ), .o1(new_n326));
  oaib12aa1n02x5               g231(.a(new_n319), .b(new_n326), .c(\a[28] ), .out0(new_n327));
  aoai13aa1n02x7               g232(.a(new_n327), .b(new_n325), .c(new_n307), .d(new_n309), .o1(new_n328));
  nand02aa1n02x5               g233(.a(new_n328), .b(new_n323), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n327), .b(new_n323), .out0(new_n330));
  aoai13aa1n02x7               g235(.a(new_n330), .b(new_n325), .c(new_n307), .d(new_n309), .o1(new_n331));
  nanp02aa1n03x5               g236(.a(new_n329), .b(new_n331), .o1(\s[29] ));
  xorb03aa1n02x5               g237(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n09x5               g238(.a(new_n323), .b(new_n311), .c(new_n317), .out0(new_n334));
  oaoi03aa1n02x5               g239(.a(\a[29] ), .b(\b[28] ), .c(new_n327), .o1(new_n335));
  xnrc02aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n335), .c(new_n310), .d(new_n334), .o1(new_n337));
  inv000aa1d42x5               g242(.a(new_n334), .o1(new_n338));
  norp02aa1n02x5               g243(.a(new_n335), .b(new_n336), .o1(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n338), .c(new_n307), .d(new_n309), .o1(new_n340));
  nanp02aa1n03x5               g245(.a(new_n337), .b(new_n340), .o1(\s[30] ));
  nano23aa1n02x4               g246(.a(new_n336), .b(new_n323), .c(new_n317), .d(new_n311), .out0(new_n342));
  nanp02aa1n03x5               g247(.a(new_n310), .b(new_n342), .o1(new_n343));
  norb02aa1n02x5               g248(.a(new_n335), .b(new_n336), .out0(new_n344));
  oab012aa1n02x4               g249(.a(new_n344), .b(\a[30] ), .c(\b[29] ), .out0(new_n345));
  xorc02aa1n02x5               g250(.a(\a[31] ), .b(\b[30] ), .out0(new_n346));
  inv000aa1n02x5               g251(.a(new_n342), .o1(new_n347));
  oai022aa1n02x5               g252(.a(\a[30] ), .b(\b[29] ), .c(\b[30] ), .d(\a[31] ), .o1(new_n348));
  aoi112aa1n02x5               g253(.a(new_n344), .b(new_n348), .c(\a[31] ), .d(\b[30] ), .o1(new_n349));
  aoai13aa1n02x7               g254(.a(new_n349), .b(new_n347), .c(new_n307), .d(new_n309), .o1(new_n350));
  aoai13aa1n03x5               g255(.a(new_n350), .b(new_n346), .c(new_n343), .d(new_n345), .o1(\s[31] ));
  nanp03aa1n02x5               g256(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n107), .b(new_n352), .c(new_n98), .out0(\s[3] ));
  inv000aa1d42x5               g258(.a(new_n105), .o1(new_n354));
  nanp02aa1n02x5               g259(.a(new_n101), .b(new_n107), .o1(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n104), .b(new_n355), .c(new_n354), .out0(\s[4] ));
  norb02aa1n02x5               g261(.a(new_n117), .b(new_n116), .out0(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n357), .b(new_n108), .c(new_n109), .out0(\s[5] ));
  aobi12aa1n02x5               g263(.a(new_n357), .b(new_n108), .c(new_n109), .out0(new_n359));
  obai22aa1n02x7               g264(.a(new_n114), .b(new_n115), .c(new_n359), .d(new_n116), .out0(new_n360));
  norb03aa1n02x5               g265(.a(new_n114), .b(new_n116), .c(new_n115), .out0(new_n361));
  oaib12aa1n02x5               g266(.a(new_n360), .b(new_n359), .c(new_n361), .out0(\s[6] ));
  oai012aa1n02x5               g267(.a(new_n114), .b(new_n116), .c(new_n115), .o1(new_n363));
  nanp02aa1n02x5               g268(.a(new_n151), .b(new_n118), .o1(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n113), .b(new_n364), .c(new_n363), .out0(\s[7] ));
  aob012aa1n02x5               g270(.a(new_n113), .b(new_n364), .c(new_n363), .out0(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n110), .b(new_n366), .c(new_n124), .out0(\s[8] ));
  aoi113aa1n02x5               g272(.a(new_n125), .b(new_n129), .c(new_n121), .d(new_n122), .e(new_n123), .o1(new_n368));
  aoi022aa1n02x5               g273(.a(new_n127), .b(new_n129), .c(new_n154), .d(new_n368), .o1(\s[9] ));
endmodule


