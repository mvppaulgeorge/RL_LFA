// Benchmark "adder" written by ABC on Wed Jul 17 14:01:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n310,
    new_n313, new_n314, new_n316, new_n317, new_n318, new_n320;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor042aa1n06x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand22aa1n09x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  and002aa1n12x5               g005(.a(\b[3] ), .b(\a[4] ), .o(new_n101));
  inv040aa1d32x5               g006(.a(\a[3] ), .o1(new_n102));
  inv040aa1d28x5               g007(.a(\b[2] ), .o1(new_n103));
  nand02aa1n08x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nand02aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1d04x5               g010(.a(new_n104), .b(new_n105), .o1(new_n106));
  nand42aa1d28x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nor042aa1d18x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nand02aa1d28x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  oai012aa1d24x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\a[4] ), .o1(new_n111));
  aboi22aa1d24x5               g016(.a(\b[3] ), .b(new_n111), .c(new_n102), .d(new_n103), .out0(new_n112));
  oaoi13aa1n12x5               g017(.a(new_n101), .b(new_n112), .c(new_n110), .d(new_n106), .o1(new_n113));
  nor042aa1n06x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand02aa1d24x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  norb02aa1n06x5               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  nor002aa1d32x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nand02aa1d28x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nanb02aa1d36x5               g023(.a(new_n117), .b(new_n118), .out0(new_n119));
  nor042aa1n04x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nand02aa1d20x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  norb02aa1n06x4               g026(.a(new_n121), .b(new_n120), .out0(new_n122));
  xnrc02aa1n12x5               g027(.a(\b[4] ), .b(\a[5] ), .out0(new_n123));
  nano23aa1n09x5               g028(.a(new_n123), .b(new_n119), .c(new_n116), .d(new_n122), .out0(new_n124));
  nanp02aa1n02x5               g029(.a(new_n113), .b(new_n124), .o1(new_n125));
  nano23aa1n03x7               g030(.a(new_n114), .b(new_n117), .c(new_n118), .d(new_n115), .out0(new_n126));
  orn002aa1n03x5               g031(.a(\a[5] ), .b(\b[4] ), .o(new_n127));
  oaoi03aa1n06x5               g032(.a(\a[6] ), .b(\b[5] ), .c(new_n127), .o1(new_n128));
  oaih12aa1n02x5               g033(.a(new_n115), .b(new_n117), .c(new_n114), .o1(new_n129));
  aobi12aa1n06x5               g034(.a(new_n129), .b(new_n126), .c(new_n128), .out0(new_n130));
  oai112aa1n06x5               g035(.a(new_n125), .b(new_n130), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  xobna2aa1n03x5               g036(.a(new_n99), .b(new_n131), .c(new_n100), .out0(\s[10] ));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nand42aa1d28x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv000aa1n09x5               g040(.a(new_n98), .o1(new_n136));
  aoai13aa1n06x5               g041(.a(new_n136), .b(new_n97), .c(new_n131), .d(new_n100), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n134), .c(new_n135), .out0(\s[11] ));
  nanb02aa1n02x5               g043(.a(new_n133), .b(new_n135), .out0(new_n139));
  nor002aa1d24x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(new_n142));
  oai112aa1n03x5               g047(.a(new_n134), .b(new_n142), .c(new_n137), .d(new_n139), .o1(new_n143));
  oaoi13aa1n06x5               g048(.a(new_n142), .b(new_n134), .c(new_n137), .d(new_n139), .o1(new_n144));
  norb02aa1n03x4               g049(.a(new_n143), .b(new_n144), .out0(\s[12] ));
  xnrc02aa1n12x5               g050(.a(\b[12] ), .b(\a[13] ), .out0(new_n146));
  nona23aa1d18x5               g051(.a(new_n141), .b(new_n135), .c(new_n133), .d(new_n140), .out0(new_n147));
  nor022aa1n16x5               g052(.a(\b[8] ), .b(\a[9] ), .o1(new_n148));
  oai012aa1n12x5               g053(.a(new_n136), .b(new_n148), .c(new_n97), .o1(new_n149));
  oai012aa1d24x5               g054(.a(new_n141), .b(new_n140), .c(new_n133), .o1(new_n150));
  oai012aa1n18x5               g055(.a(new_n150), .b(new_n147), .c(new_n149), .o1(new_n151));
  inv040aa1n03x5               g056(.a(new_n151), .o1(new_n152));
  aob012aa1n06x5               g057(.a(new_n129), .b(new_n126), .c(new_n128), .out0(new_n153));
  nano23aa1d15x5               g058(.a(new_n133), .b(new_n140), .c(new_n141), .d(new_n135), .out0(new_n154));
  norb02aa1n12x5               g059(.a(new_n100), .b(new_n148), .out0(new_n155));
  nand23aa1d12x5               g060(.a(new_n154), .b(new_n99), .c(new_n155), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n153), .c(new_n113), .d(new_n124), .o1(new_n158));
  xobna2aa1n03x5               g063(.a(new_n146), .b(new_n158), .c(new_n152), .out0(\s[13] ));
  orn002aa1n02x7               g064(.a(\a[13] ), .b(\b[12] ), .o(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n146), .c(new_n158), .d(new_n152), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xnrc02aa1n12x5               g067(.a(\b[13] ), .b(\a[14] ), .out0(new_n163));
  nor042aa1n04x5               g068(.a(new_n163), .b(new_n146), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  oao003aa1n03x5               g070(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .carry(new_n166));
  aoai13aa1n04x5               g071(.a(new_n166), .b(new_n165), .c(new_n158), .d(new_n152), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n09x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand02aa1d28x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nor042aa1n06x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nand02aa1d20x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoi112aa1n03x5               g078(.a(new_n173), .b(new_n169), .c(new_n167), .d(new_n170), .o1(new_n174));
  aoai13aa1n03x5               g079(.a(new_n173), .b(new_n169), .c(new_n167), .d(new_n170), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[16] ));
  nano23aa1d15x5               g081(.a(new_n169), .b(new_n171), .c(new_n172), .d(new_n170), .out0(new_n177));
  nona22aa1n12x5               g082(.a(new_n177), .b(new_n163), .c(new_n146), .out0(new_n178));
  nor042aa1n09x5               g083(.a(new_n178), .b(new_n156), .o1(new_n179));
  aoai13aa1n12x5               g084(.a(new_n179), .b(new_n153), .c(new_n113), .d(new_n124), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n172), .b(new_n171), .c(new_n169), .o1(new_n181));
  oaib12aa1n09x5               g086(.a(new_n181), .b(new_n166), .c(new_n177), .out0(new_n182));
  aoi013aa1n09x5               g087(.a(new_n182), .b(new_n151), .c(new_n164), .d(new_n177), .o1(new_n183));
  nanp02aa1n09x5               g088(.a(new_n180), .b(new_n183), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g090(.a(\a[18] ), .o1(new_n186));
  inv040aa1d32x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  oaoi03aa1n03x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n186), .out0(\s[18] ));
  xroi22aa1d06x4               g095(.a(new_n187), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(new_n188), .b(new_n187), .o1(new_n192));
  oaoi03aa1n09x5               g097(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n193));
  nor002aa1d32x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand02aa1d06x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n193), .c(new_n184), .d(new_n191), .o1(new_n197));
  aoi112aa1n02x5               g102(.a(new_n196), .b(new_n193), .c(new_n184), .d(new_n191), .o1(new_n198));
  norb02aa1n02x7               g103(.a(new_n197), .b(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n12x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand02aa1n06x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  nona22aa1n02x5               g108(.a(new_n197), .b(new_n203), .c(new_n194), .out0(new_n204));
  inv040aa1n08x5               g109(.a(new_n194), .o1(new_n205));
  aobi12aa1n06x5               g110(.a(new_n203), .b(new_n197), .c(new_n205), .out0(new_n206));
  norb02aa1n03x4               g111(.a(new_n204), .b(new_n206), .out0(\s[20] ));
  nano23aa1n03x7               g112(.a(new_n194), .b(new_n201), .c(new_n202), .d(new_n195), .out0(new_n208));
  nanp02aa1n02x5               g113(.a(new_n191), .b(new_n208), .o1(new_n209));
  oaih22aa1n06x5               g114(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n210));
  oaib12aa1n18x5               g115(.a(new_n210), .b(new_n186), .c(\b[17] ), .out0(new_n211));
  nona23aa1n12x5               g116(.a(new_n202), .b(new_n195), .c(new_n194), .d(new_n201), .out0(new_n212));
  oaoi03aa1n06x5               g117(.a(\a[20] ), .b(\b[19] ), .c(new_n205), .o1(new_n213));
  inv040aa1n03x5               g118(.a(new_n213), .o1(new_n214));
  oai012aa1d24x5               g119(.a(new_n214), .b(new_n212), .c(new_n211), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n04x5               g121(.a(new_n216), .b(new_n209), .c(new_n180), .d(new_n183), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[21] ), .b(\b[20] ), .out0(new_n220));
  xorc02aa1n02x5               g125(.a(\a[22] ), .b(\b[21] ), .out0(new_n221));
  aoi112aa1n02x5               g126(.a(new_n219), .b(new_n221), .c(new_n217), .d(new_n220), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n221), .b(new_n219), .c(new_n217), .d(new_n220), .o1(new_n223));
  norb02aa1n03x4               g128(.a(new_n223), .b(new_n222), .out0(\s[22] ));
  inv000aa1d42x5               g129(.a(\a[21] ), .o1(new_n225));
  inv040aa1d32x5               g130(.a(\a[22] ), .o1(new_n226));
  xroi22aa1d06x4               g131(.a(new_n225), .b(\b[20] ), .c(new_n226), .d(\b[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(\b[21] ), .o1(new_n228));
  oao003aa1n02x5               g133(.a(new_n226), .b(new_n228), .c(new_n219), .carry(new_n229));
  aoi012aa1n02x5               g134(.a(new_n229), .b(new_n215), .c(new_n227), .o1(new_n230));
  nanp03aa1n02x5               g135(.a(new_n227), .b(new_n191), .c(new_n208), .o1(new_n231));
  aoai13aa1n06x5               g136(.a(new_n230), .b(new_n231), .c(new_n180), .d(new_n183), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  xorc02aa1n02x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  xorc02aa1n02x5               g140(.a(\a[24] ), .b(\b[23] ), .out0(new_n236));
  aoi112aa1n02x5               g141(.a(new_n234), .b(new_n236), .c(new_n232), .d(new_n235), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n234), .c(new_n232), .d(new_n235), .o1(new_n238));
  norb02aa1n03x4               g143(.a(new_n238), .b(new_n237), .out0(\s[24] ));
  inv000aa1d42x5               g144(.a(\a[23] ), .o1(new_n240));
  inv040aa1d32x5               g145(.a(\a[24] ), .o1(new_n241));
  xroi22aa1d06x4               g146(.a(new_n240), .b(\b[22] ), .c(new_n241), .d(\b[23] ), .out0(new_n242));
  nano22aa1n02x4               g147(.a(new_n209), .b(new_n227), .c(new_n242), .out0(new_n243));
  aoai13aa1n03x5               g148(.a(new_n227), .b(new_n213), .c(new_n208), .d(new_n193), .o1(new_n244));
  inv000aa1n02x5               g149(.a(new_n229), .o1(new_n245));
  inv000aa1n02x5               g150(.a(new_n242), .o1(new_n246));
  oai022aa1n02x5               g151(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n247));
  oaib12aa1n02x5               g152(.a(new_n247), .b(new_n241), .c(\b[23] ), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n246), .c(new_n244), .d(new_n245), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[25] ), .b(\b[24] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(new_n184), .d(new_n243), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(new_n250), .b(new_n249), .c(new_n184), .d(new_n243), .o1(new_n252));
  norb02aa1n02x7               g157(.a(new_n251), .b(new_n252), .out0(\s[25] ));
  nor042aa1n03x5               g158(.a(\b[24] ), .b(\a[25] ), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[26] ), .b(\b[25] ), .out0(new_n255));
  nona22aa1n02x5               g160(.a(new_n251), .b(new_n255), .c(new_n254), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n254), .o1(new_n257));
  aobi12aa1n06x5               g162(.a(new_n255), .b(new_n251), .c(new_n257), .out0(new_n258));
  norb02aa1n03x4               g163(.a(new_n256), .b(new_n258), .out0(\s[26] ));
  nanp02aa1n02x5               g164(.a(new_n125), .b(new_n130), .o1(new_n260));
  oabi12aa1n02x5               g165(.a(new_n182), .b(new_n152), .c(new_n178), .out0(new_n261));
  inv020aa1d32x5               g166(.a(\a[25] ), .o1(new_n262));
  inv020aa1n04x5               g167(.a(\a[26] ), .o1(new_n263));
  xroi22aa1d06x4               g168(.a(new_n262), .b(\b[24] ), .c(new_n263), .d(\b[25] ), .out0(new_n264));
  nano32aa1n03x7               g169(.a(new_n209), .b(new_n264), .c(new_n227), .d(new_n242), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n261), .c(new_n260), .d(new_n179), .o1(new_n266));
  oao003aa1n02x5               g171(.a(\a[26] ), .b(\b[25] ), .c(new_n257), .carry(new_n267));
  aobi12aa1n06x5               g172(.a(new_n267), .b(new_n249), .c(new_n264), .out0(new_n268));
  nor042aa1n04x5               g173(.a(\b[26] ), .b(\a[27] ), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n270), .b(new_n269), .out0(new_n271));
  xnbna2aa1n03x5               g176(.a(new_n271), .b(new_n268), .c(new_n266), .out0(\s[27] ));
  xorc02aa1n02x5               g177(.a(\a[28] ), .b(\b[27] ), .out0(new_n273));
  aobi12aa1n06x5               g178(.a(new_n265), .b(new_n180), .c(new_n183), .out0(new_n274));
  aoai13aa1n02x5               g179(.a(new_n242), .b(new_n229), .c(new_n215), .d(new_n227), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n264), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n267), .b(new_n276), .c(new_n275), .d(new_n248), .o1(new_n277));
  norp03aa1n03x5               g182(.a(new_n277), .b(new_n274), .c(new_n269), .o1(new_n278));
  nano22aa1n03x7               g183(.a(new_n278), .b(new_n270), .c(new_n273), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n269), .o1(new_n280));
  nanp03aa1n03x5               g185(.a(new_n268), .b(new_n266), .c(new_n280), .o1(new_n281));
  aoi012aa1n03x5               g186(.a(new_n273), .b(new_n281), .c(new_n270), .o1(new_n282));
  nor042aa1n03x5               g187(.a(new_n282), .b(new_n279), .o1(\s[28] ));
  and002aa1n02x5               g188(.a(new_n273), .b(new_n271), .o(new_n284));
  oaih12aa1n02x5               g189(.a(new_n284), .b(new_n277), .c(new_n274), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[28] ), .b(\a[29] ), .out0(new_n287));
  tech160nm_fiaoi012aa1n02p5x5 g192(.a(new_n287), .b(new_n285), .c(new_n286), .o1(new_n288));
  aobi12aa1n02x7               g193(.a(new_n284), .b(new_n268), .c(new_n266), .out0(new_n289));
  nano22aa1n02x4               g194(.a(new_n289), .b(new_n286), .c(new_n287), .out0(new_n290));
  norp02aa1n03x5               g195(.a(new_n288), .b(new_n290), .o1(\s[29] ));
  xorb03aa1n02x5               g196(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g197(.a(new_n287), .b(new_n273), .c(new_n271), .out0(new_n293));
  oaih12aa1n02x5               g198(.a(new_n293), .b(new_n277), .c(new_n274), .o1(new_n294));
  oao003aa1n02x5               g199(.a(\a[29] ), .b(\b[28] ), .c(new_n286), .carry(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[29] ), .b(\a[30] ), .out0(new_n296));
  tech160nm_fiaoi012aa1n02p5x5 g201(.a(new_n296), .b(new_n294), .c(new_n295), .o1(new_n297));
  aobi12aa1n02x7               g202(.a(new_n293), .b(new_n268), .c(new_n266), .out0(new_n298));
  nano22aa1n03x5               g203(.a(new_n298), .b(new_n295), .c(new_n296), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[30] ));
  nano23aa1n02x4               g205(.a(new_n296), .b(new_n287), .c(new_n273), .d(new_n271), .out0(new_n301));
  aobi12aa1n02x7               g206(.a(new_n301), .b(new_n268), .c(new_n266), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n295), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  nano22aa1n02x4               g209(.a(new_n302), .b(new_n303), .c(new_n304), .out0(new_n305));
  oaih12aa1n02x5               g210(.a(new_n301), .b(new_n277), .c(new_n274), .o1(new_n306));
  tech160nm_fiaoi012aa1n02p5x5 g211(.a(new_n304), .b(new_n306), .c(new_n303), .o1(new_n307));
  norp02aa1n03x5               g212(.a(new_n307), .b(new_n305), .o1(\s[31] ));
  xnbna2aa1n03x5               g213(.a(new_n110), .b(new_n104), .c(new_n105), .out0(\s[3] ));
  oaoi03aa1n02x5               g214(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g216(.a(new_n113), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1n03x5               g217(.a(new_n113), .o1(new_n313));
  oaoi03aa1n02x5               g218(.a(\a[5] ), .b(\b[4] ), .c(new_n313), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g220(.a(new_n119), .o1(new_n316));
  oai112aa1n03x5               g221(.a(new_n316), .b(new_n121), .c(new_n314), .d(new_n120), .o1(new_n317));
  oaoi13aa1n02x5               g222(.a(new_n316), .b(new_n121), .c(new_n314), .d(new_n120), .o1(new_n318));
  norb02aa1n02x5               g223(.a(new_n317), .b(new_n318), .out0(\s[7] ));
  inv000aa1d42x5               g224(.a(new_n117), .o1(new_n320));
  xnbna2aa1n03x5               g225(.a(new_n116), .b(new_n317), .c(new_n320), .out0(\s[8] ));
  xnbna2aa1n03x5               g226(.a(new_n155), .b(new_n125), .c(new_n130), .out0(\s[9] ));
endmodule


