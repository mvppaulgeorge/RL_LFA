// Benchmark "adder" written by ABC on Thu Jul 18 07:19:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n316, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n337,
    new_n338, new_n339, new_n340, new_n342, new_n344, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n352, new_n353, new_n355, new_n356,
    new_n358, new_n359, new_n360;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n16x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand23aa1n06x5               g005(.a(new_n100), .b(\a[1] ), .c(\b[0] ), .o1(new_n101));
  aoi022aa1d24x5               g006(.a(\b[2] ), .b(\a[3] ), .c(\a[2] ), .d(\b[1] ), .o1(new_n102));
  nor002aa1n20x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1d28x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb03aa1d15x5               g010(.a(new_n105), .b(new_n103), .c(new_n104), .out0(new_n106));
  oai112aa1n06x5               g011(.a(new_n106), .b(new_n102), .c(new_n101), .d(new_n99), .o1(new_n107));
  tech160nm_fioai012aa1n03p5x5 g012(.a(new_n105), .b(new_n104), .c(new_n103), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1d28x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor042aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand42aa1n10x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nano23aa1n03x5               g017(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n113));
  nor002aa1n03x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  tech160nm_finand02aa1n05x5   g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nor042aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand42aa1n08x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nano23aa1n02x5               g022(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n118));
  nand02aa1n02x5               g023(.a(new_n118), .b(new_n113), .o1(new_n119));
  aoi112aa1n09x5               g024(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n120));
  oai022aa1d18x5               g025(.a(\a[6] ), .b(\b[5] ), .c(\b[6] ), .d(\a[7] ), .o1(new_n121));
  aoi022aa1n06x5               g026(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n122));
  oaoi13aa1n09x5               g027(.a(new_n114), .b(new_n122), .c(new_n120), .d(new_n121), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n123), .b(new_n119), .c(new_n107), .d(new_n108), .o1(new_n124));
  nand42aa1n08x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n03x5               g030(.a(new_n125), .b(new_n97), .out0(new_n126));
  nanp02aa1n02x5               g031(.a(new_n124), .b(new_n126), .o1(new_n127));
  nor002aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1n06x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n03x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  aoai13aa1n06x5               g036(.a(new_n130), .b(new_n97), .c(new_n124), .d(new_n125), .o1(new_n132));
  oai012aa1n02x5               g037(.a(new_n129), .b(new_n128), .c(new_n97), .o1(new_n133));
  nor042aa1n09x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n12x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n132), .c(new_n133), .out0(\s[11] ));
  nand22aa1n03x5               g042(.a(new_n132), .b(new_n133), .o1(new_n138));
  nor002aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n134), .c(new_n138), .d(new_n136), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(new_n138), .b(new_n136), .o1(new_n143));
  nona22aa1n02x4               g048(.a(new_n143), .b(new_n141), .c(new_n134), .out0(new_n144));
  nanp02aa1n02x5               g049(.a(new_n144), .b(new_n142), .o1(\s[12] ));
  nano32aa1n02x4               g050(.a(new_n141), .b(new_n136), .c(new_n130), .d(new_n126), .out0(new_n146));
  nand22aa1n03x5               g051(.a(new_n124), .b(new_n146), .o1(new_n147));
  tech160nm_fioaoi03aa1n03p5x5 g052(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n148));
  nano23aa1n06x5               g053(.a(new_n134), .b(new_n139), .c(new_n140), .d(new_n135), .out0(new_n149));
  oai012aa1n03x5               g054(.a(new_n140), .b(new_n139), .c(new_n134), .o1(new_n150));
  aobi12aa1n06x5               g055(.a(new_n150), .b(new_n149), .c(new_n148), .out0(new_n151));
  nanp02aa1n03x5               g056(.a(new_n147), .b(new_n151), .o1(new_n152));
  nor002aa1n10x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand02aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  nanp02aa1n02x5               g060(.a(new_n149), .b(new_n148), .o1(new_n156));
  nano22aa1n02x4               g061(.a(new_n155), .b(new_n156), .c(new_n150), .out0(new_n157));
  aoi022aa1n02x5               g062(.a(new_n152), .b(new_n155), .c(new_n147), .d(new_n157), .o1(\s[13] ));
  tech160nm_fiaoi012aa1n05x5   g063(.a(new_n153), .b(new_n152), .c(new_n154), .o1(new_n159));
  xnrb03aa1n03x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nanp02aa1n02x5               g065(.a(new_n156), .b(new_n150), .o1(new_n161));
  nor002aa1n04x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nanp02aa1n04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nano23aa1n09x5               g068(.a(new_n153), .b(new_n162), .c(new_n163), .d(new_n154), .out0(new_n164));
  aoai13aa1n03x5               g069(.a(new_n164), .b(new_n161), .c(new_n124), .d(new_n146), .o1(new_n165));
  oai012aa1n04x7               g070(.a(new_n163), .b(new_n162), .c(new_n153), .o1(new_n166));
  nor042aa1n06x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n04x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n165), .c(new_n166), .out0(\s[15] ));
  nanp02aa1n03x5               g075(.a(new_n165), .b(new_n166), .o1(new_n171));
  nor042aa1n06x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  aoai13aa1n03x5               g079(.a(new_n174), .b(new_n167), .c(new_n171), .d(new_n169), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n171), .b(new_n169), .o1(new_n176));
  nona22aa1n02x4               g081(.a(new_n176), .b(new_n174), .c(new_n167), .out0(new_n177));
  nanp02aa1n02x5               g082(.a(new_n177), .b(new_n175), .o1(\s[16] ));
  nano23aa1n09x5               g083(.a(new_n167), .b(new_n172), .c(new_n173), .d(new_n168), .out0(new_n179));
  nand02aa1d04x5               g084(.a(new_n179), .b(new_n164), .o1(new_n180));
  nano32aa1n06x5               g085(.a(new_n180), .b(new_n149), .c(new_n130), .d(new_n126), .out0(new_n181));
  nanp02aa1n09x5               g086(.a(new_n124), .b(new_n181), .o1(new_n182));
  inv000aa1n02x5               g087(.a(new_n180), .o1(new_n183));
  nona23aa1n03x5               g088(.a(new_n173), .b(new_n168), .c(new_n167), .d(new_n172), .out0(new_n184));
  tech160nm_fioai012aa1n03p5x5 g089(.a(new_n173), .b(new_n172), .c(new_n167), .o1(new_n185));
  tech160nm_fioai012aa1n04x5   g090(.a(new_n185), .b(new_n184), .c(new_n166), .o1(new_n186));
  aoi012aa1n06x5               g091(.a(new_n186), .b(new_n161), .c(new_n183), .o1(new_n187));
  nand02aa1d10x5               g092(.a(new_n182), .b(new_n187), .o1(new_n188));
  nor042aa1n12x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  nand42aa1d28x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n190), .b(new_n189), .out0(new_n191));
  oaib12aa1n02x5               g096(.a(new_n185), .b(new_n189), .c(new_n190), .out0(new_n192));
  oabi12aa1n02x5               g097(.a(new_n192), .b(new_n166), .c(new_n184), .out0(new_n193));
  aoi012aa1n02x5               g098(.a(new_n193), .b(new_n161), .c(new_n183), .o1(new_n194));
  aoi022aa1n02x5               g099(.a(new_n188), .b(new_n191), .c(new_n182), .d(new_n194), .o1(\s[17] ));
  tech160nm_fiaoi012aa1n05x5   g100(.a(new_n189), .b(new_n188), .c(new_n191), .o1(new_n196));
  xnrb03aa1n03x5               g101(.a(new_n196), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  oabi12aa1n09x5               g102(.a(new_n186), .b(new_n151), .c(new_n180), .out0(new_n198));
  nor042aa1n09x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nand42aa1n20x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nano23aa1d15x5               g105(.a(new_n189), .b(new_n199), .c(new_n200), .d(new_n190), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n198), .c(new_n124), .d(new_n181), .o1(new_n202));
  nor042aa1n03x5               g107(.a(new_n199), .b(new_n189), .o1(new_n203));
  norb02aa1n06x4               g108(.a(new_n200), .b(new_n203), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  nor002aa1n06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand42aa1n06x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  norb02aa1n09x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n202), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g115(.a(new_n202), .b(new_n205), .o1(new_n211));
  nor042aa1n09x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nanp02aa1n24x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanb02aa1n12x5               g118(.a(new_n212), .b(new_n213), .out0(new_n214));
  aoai13aa1n02x7               g119(.a(new_n214), .b(new_n206), .c(new_n211), .d(new_n207), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n208), .b(new_n204), .c(new_n188), .d(new_n201), .o1(new_n216));
  nona22aa1n03x5               g121(.a(new_n216), .b(new_n214), .c(new_n206), .out0(new_n217));
  nanp02aa1n03x5               g122(.a(new_n215), .b(new_n217), .o1(\s[20] ));
  nanb03aa1d24x5               g123(.a(new_n214), .b(new_n201), .c(new_n208), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n198), .c(new_n124), .d(new_n181), .o1(new_n221));
  oai012aa1n09x5               g126(.a(new_n213), .b(new_n212), .c(new_n206), .o1(new_n222));
  nanb03aa1n02x5               g127(.a(new_n212), .b(new_n213), .c(new_n207), .out0(new_n223));
  oai022aa1n02x5               g128(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n224));
  oai112aa1n02x5               g129(.a(new_n224), .b(new_n200), .c(\b[18] ), .d(\a[19] ), .o1(new_n225));
  tech160nm_fioai012aa1n03p5x5 g130(.a(new_n222), .b(new_n225), .c(new_n223), .o1(new_n226));
  nanb02aa1n02x5               g131(.a(new_n226), .b(new_n221), .out0(new_n227));
  xorc02aa1n12x5               g132(.a(\a[21] ), .b(\b[20] ), .out0(new_n228));
  inv040aa1n03x5               g133(.a(new_n222), .o1(new_n229));
  nano22aa1n12x5               g134(.a(new_n212), .b(new_n207), .c(new_n213), .out0(new_n230));
  oai012aa1n06x5               g135(.a(new_n200), .b(\b[18] ), .c(\a[19] ), .o1(new_n231));
  oab012aa1n02x4               g136(.a(new_n231), .b(new_n189), .c(new_n199), .out0(new_n232));
  aoi112aa1n02x5               g137(.a(new_n228), .b(new_n229), .c(new_n232), .d(new_n230), .o1(new_n233));
  aoi022aa1n02x5               g138(.a(new_n227), .b(new_n228), .c(new_n221), .d(new_n233), .o1(\s[21] ));
  nor042aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  tech160nm_fixnrc02aa1n05x5   g140(.a(\b[21] ), .b(\a[22] ), .out0(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n235), .c(new_n227), .d(new_n228), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n228), .b(new_n226), .c(new_n188), .d(new_n220), .o1(new_n238));
  nona22aa1n02x4               g143(.a(new_n238), .b(new_n236), .c(new_n235), .out0(new_n239));
  nanp02aa1n02x5               g144(.a(new_n237), .b(new_n239), .o1(\s[22] ));
  nanb02aa1n12x5               g145(.a(new_n236), .b(new_n228), .out0(new_n241));
  nor042aa1n02x5               g146(.a(new_n219), .b(new_n241), .o1(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n198), .c(new_n124), .d(new_n181), .o1(new_n243));
  nona22aa1n09x5               g148(.a(new_n230), .b(new_n203), .c(new_n231), .out0(new_n244));
  inv000aa1d42x5               g149(.a(\a[22] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\b[21] ), .o1(new_n246));
  oao003aa1n09x5               g151(.a(new_n245), .b(new_n246), .c(new_n235), .carry(new_n247));
  inv040aa1n06x5               g152(.a(new_n247), .o1(new_n248));
  aoai13aa1n12x5               g153(.a(new_n248), .b(new_n241), .c(new_n244), .d(new_n222), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  nanp02aa1n02x5               g155(.a(new_n243), .b(new_n250), .o1(new_n251));
  xorc02aa1n12x5               g156(.a(\a[23] ), .b(\b[22] ), .out0(new_n252));
  xnrc02aa1n02x5               g157(.a(\b[20] ), .b(\a[21] ), .out0(new_n253));
  nor042aa1n03x5               g158(.a(new_n236), .b(new_n253), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n252), .b(new_n247), .c(new_n226), .d(new_n254), .o1(new_n255));
  aoi022aa1n02x5               g160(.a(new_n251), .b(new_n252), .c(new_n243), .d(new_n255), .o1(\s[23] ));
  nor002aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  xnrc02aa1n02x5               g162(.a(\b[23] ), .b(\a[24] ), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n257), .c(new_n251), .d(new_n252), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n252), .b(new_n249), .c(new_n188), .d(new_n242), .o1(new_n260));
  nona22aa1n03x5               g165(.a(new_n260), .b(new_n258), .c(new_n257), .out0(new_n261));
  nanp02aa1n02x5               g166(.a(new_n259), .b(new_n261), .o1(\s[24] ));
  norb02aa1n03x5               g167(.a(new_n252), .b(new_n258), .out0(new_n263));
  nano22aa1n03x7               g168(.a(new_n219), .b(new_n263), .c(new_n254), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n198), .c(new_n124), .d(new_n181), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n254), .b(new_n229), .c(new_n232), .d(new_n230), .o1(new_n266));
  inv000aa1n02x5               g171(.a(new_n263), .o1(new_n267));
  inv000aa1d42x5               g172(.a(\a[24] ), .o1(new_n268));
  inv000aa1d42x5               g173(.a(\b[23] ), .o1(new_n269));
  oao003aa1n02x5               g174(.a(new_n268), .b(new_n269), .c(new_n257), .carry(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n267), .c(new_n266), .d(new_n248), .o1(new_n272));
  nanb02aa1n02x5               g177(.a(new_n272), .b(new_n265), .out0(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoi112aa1n02x5               g179(.a(new_n274), .b(new_n270), .c(new_n249), .d(new_n263), .o1(new_n275));
  aoi022aa1n02x5               g180(.a(new_n273), .b(new_n274), .c(new_n265), .d(new_n275), .o1(\s[25] ));
  norp02aa1n02x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  nor002aa1n02x5               g182(.a(\b[25] ), .b(\a[26] ), .o1(new_n278));
  nand42aa1n02x5               g183(.a(\b[25] ), .b(\a[26] ), .o1(new_n279));
  nanb02aa1n06x5               g184(.a(new_n278), .b(new_n279), .out0(new_n280));
  aoai13aa1n02x7               g185(.a(new_n280), .b(new_n277), .c(new_n273), .d(new_n274), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n274), .b(new_n272), .c(new_n188), .d(new_n264), .o1(new_n282));
  nona22aa1n02x4               g187(.a(new_n282), .b(new_n280), .c(new_n277), .out0(new_n283));
  nanp02aa1n02x5               g188(.a(new_n281), .b(new_n283), .o1(\s[26] ));
  norb02aa1n06x4               g189(.a(new_n274), .b(new_n280), .out0(new_n285));
  inv000aa1n02x5               g190(.a(new_n285), .o1(new_n286));
  nano23aa1d15x5               g191(.a(new_n286), .b(new_n219), .c(new_n263), .d(new_n254), .out0(new_n287));
  aoai13aa1n09x5               g192(.a(new_n287), .b(new_n198), .c(new_n124), .d(new_n181), .o1(new_n288));
  oai012aa1n02x5               g193(.a(new_n279), .b(new_n278), .c(new_n277), .o1(new_n289));
  aobi12aa1n06x5               g194(.a(new_n289), .b(new_n272), .c(new_n285), .out0(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnbna2aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n288), .out0(\s[27] ));
  aoai13aa1n04x5               g197(.a(new_n285), .b(new_n270), .c(new_n249), .d(new_n263), .o1(new_n293));
  nand23aa1n04x5               g198(.a(new_n288), .b(new_n293), .c(new_n289), .o1(new_n294));
  nor002aa1d32x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  nor042aa1n06x5               g200(.a(\b[27] ), .b(\a[28] ), .o1(new_n296));
  nand42aa1n08x5               g201(.a(\b[27] ), .b(\a[28] ), .o1(new_n297));
  nanb02aa1n02x5               g202(.a(new_n296), .b(new_n297), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n295), .c(new_n294), .d(new_n291), .o1(new_n299));
  aoai13aa1n02x5               g204(.a(new_n263), .b(new_n247), .c(new_n226), .d(new_n254), .o1(new_n300));
  aoai13aa1n02x7               g205(.a(new_n289), .b(new_n286), .c(new_n300), .d(new_n271), .o1(new_n301));
  aoai13aa1n02x5               g206(.a(new_n291), .b(new_n301), .c(new_n188), .d(new_n287), .o1(new_n302));
  nona22aa1n02x4               g207(.a(new_n302), .b(new_n298), .c(new_n295), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n299), .b(new_n303), .o1(\s[28] ));
  norb02aa1n02x7               g209(.a(new_n291), .b(new_n298), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n301), .c(new_n188), .d(new_n287), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n305), .o1(new_n307));
  oai012aa1n06x5               g212(.a(new_n297), .b(new_n296), .c(new_n295), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n307), .c(new_n290), .d(new_n288), .o1(new_n309));
  norp02aa1n02x5               g214(.a(\b[28] ), .b(\a[29] ), .o1(new_n310));
  nand42aa1n03x5               g215(.a(\b[28] ), .b(\a[29] ), .o1(new_n311));
  norb02aa1n03x5               g216(.a(new_n311), .b(new_n310), .out0(new_n312));
  oai022aa1n02x5               g217(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n313));
  aboi22aa1n03x5               g218(.a(new_n310), .b(new_n311), .c(new_n313), .d(new_n297), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n309), .b(new_n312), .c(new_n306), .d(new_n314), .o1(\s[29] ));
  nanp02aa1n02x5               g220(.a(\b[0] ), .b(\a[1] ), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g222(.a(new_n298), .b(new_n291), .c(new_n312), .out0(new_n318));
  nanb02aa1n03x5               g223(.a(new_n318), .b(new_n294), .out0(new_n319));
  tech160nm_fioaoi03aa1n02p5x5 g224(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n318), .c(new_n290), .d(new_n288), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  aoi113aa1n02x5               g228(.a(new_n323), .b(new_n310), .c(new_n313), .d(new_n311), .e(new_n297), .o1(new_n324));
  aoi022aa1n03x5               g229(.a(new_n322), .b(new_n323), .c(new_n319), .d(new_n324), .o1(\s[30] ));
  inv000aa1d42x5               g230(.a(new_n312), .o1(new_n326));
  nona23aa1n02x4               g231(.a(new_n291), .b(new_n323), .c(new_n326), .d(new_n298), .out0(new_n327));
  nanb02aa1n03x5               g232(.a(new_n327), .b(new_n294), .out0(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  inv000aa1d42x5               g234(.a(\a[30] ), .o1(new_n330));
  inv000aa1d42x5               g235(.a(\b[29] ), .o1(new_n331));
  oabi12aa1n02x5               g236(.a(new_n329), .b(\a[30] ), .c(\b[29] ), .out0(new_n332));
  oaoi13aa1n02x5               g237(.a(new_n332), .b(new_n320), .c(new_n330), .d(new_n331), .o1(new_n333));
  oaoi03aa1n02x5               g238(.a(new_n330), .b(new_n331), .c(new_n320), .o1(new_n334));
  aoai13aa1n02x7               g239(.a(new_n334), .b(new_n327), .c(new_n290), .d(new_n288), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n335), .b(new_n329), .c(new_n328), .d(new_n333), .o1(\s[31] ));
  norb03aa1n03x5               g241(.a(new_n100), .b(new_n99), .c(new_n316), .out0(new_n337));
  xorc02aa1n02x5               g242(.a(\a[3] ), .b(\b[2] ), .out0(new_n338));
  aoai13aa1n02x5               g243(.a(new_n338), .b(new_n337), .c(\a[2] ), .d(\b[1] ), .o1(new_n339));
  nona22aa1n02x4               g244(.a(new_n100), .b(new_n338), .c(new_n337), .out0(new_n340));
  nanp02aa1n02x5               g245(.a(new_n340), .b(new_n339), .o1(\s[3] ));
  aboi22aa1n03x5               g246(.a(new_n103), .b(new_n105), .c(\a[3] ), .d(\b[2] ), .out0(new_n342));
  ao0022aa1n03x5               g247(.a(new_n339), .b(new_n342), .c(new_n107), .d(new_n106), .o(\s[4] ));
  norb02aa1n02x5               g248(.a(new_n112), .b(new_n111), .out0(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n344), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  nona23aa1n02x4               g250(.a(new_n102), .b(new_n105), .c(new_n104), .d(new_n103), .out0(new_n346));
  oaih12aa1n02x5               g251(.a(new_n108), .b(new_n346), .c(new_n337), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n117), .b(new_n116), .out0(new_n348));
  aoai13aa1n03x5               g253(.a(new_n348), .b(new_n111), .c(new_n347), .d(new_n112), .o1(new_n349));
  aoi112aa1n02x5               g254(.a(new_n111), .b(new_n348), .c(new_n347), .d(new_n344), .o1(new_n350));
  norb02aa1n02x5               g255(.a(new_n349), .b(new_n350), .out0(\s[6] ));
  norb02aa1n02x5               g256(.a(new_n110), .b(new_n109), .out0(new_n352));
  aoi012aa1n02x5               g257(.a(new_n116), .b(new_n111), .c(new_n117), .o1(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n352), .b(new_n349), .c(new_n353), .out0(\s[7] ));
  nanp02aa1n03x5               g259(.a(new_n349), .b(new_n353), .o1(new_n355));
  aoi012aa1n03x5               g260(.a(new_n109), .b(new_n355), .c(new_n110), .o1(new_n356));
  xnrb03aa1n03x5               g261(.a(new_n356), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  nanb02aa1n02x5               g262(.a(new_n119), .b(new_n347), .out0(new_n358));
  obai22aa1n02x7               g263(.a(new_n125), .b(new_n97), .c(\a[8] ), .d(\b[7] ), .out0(new_n359));
  oaoi13aa1n02x5               g264(.a(new_n359), .b(new_n122), .c(new_n120), .d(new_n121), .o1(new_n360));
  aoi022aa1n02x5               g265(.a(new_n124), .b(new_n126), .c(new_n358), .d(new_n360), .o1(\s[9] ));
endmodule


