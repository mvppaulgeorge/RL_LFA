// Benchmark "adder" written by ABC on Thu Jul 18 11:23:50 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n306, new_n309, new_n310, new_n312, new_n314;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n03p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n09x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n03x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  oai012aa1n02x7               g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oai012aa1n04x7               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nor042aa1n09x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n06x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nor042aa1n03x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand02aa1n03x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nano23aa1n03x7               g018(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n114));
  nand02aa1n10x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor022aa1n08x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  orn002aa1n02x5               g021(.a(\a[8] ), .b(\b[7] ), .o(new_n117));
  and002aa1n12x5               g022(.a(\b[7] ), .b(\a[8] ), .o(new_n118));
  nona23aa1n03x5               g023(.a(new_n117), .b(new_n115), .c(new_n118), .d(new_n116), .out0(new_n119));
  norb02aa1n03x5               g024(.a(new_n114), .b(new_n119), .out0(new_n120));
  inv000aa1d42x5               g025(.a(new_n110), .o1(new_n121));
  aoai13aa1n04x5               g026(.a(new_n111), .b(new_n116), .c(new_n112), .d(new_n115), .o1(new_n122));
  aoai13aa1n06x5               g027(.a(new_n117), .b(new_n118), .c(new_n122), .d(new_n121), .o1(new_n123));
  tech160nm_fixorc02aa1n02p5x5 g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(new_n120), .d(new_n109), .o1(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n97), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  nand02aa1n03x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n10x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  nor042aa1n03x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nanb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  oai022aa1d18x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n131), .b(new_n125), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n130), .b(new_n132), .c(new_n127), .out0(\s[11] ));
  inv000aa1d42x5               g038(.a(\a[12] ), .o1(new_n134));
  aoi013aa1n02x4               g039(.a(new_n129), .b(new_n132), .c(new_n127), .d(new_n128), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[11] ), .c(new_n134), .out0(\s[12] ));
  oao003aa1n02x5               g041(.a(new_n99), .b(new_n100), .c(new_n101), .carry(new_n137));
  nano23aa1n02x4               g042(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n138));
  aobi12aa1n02x5               g043(.a(new_n108), .b(new_n138), .c(new_n137), .out0(new_n139));
  nanb02aa1d24x5               g044(.a(new_n116), .b(new_n115), .out0(new_n140));
  nona23aa1n03x5               g045(.a(new_n114), .b(new_n117), .c(new_n118), .d(new_n140), .out0(new_n141));
  oabi12aa1n06x5               g046(.a(new_n123), .b(new_n139), .c(new_n141), .out0(new_n142));
  norp02aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n03x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nano23aa1n03x7               g049(.a(new_n143), .b(new_n129), .c(new_n144), .d(new_n128), .out0(new_n145));
  and003aa1n02x5               g050(.a(new_n145), .b(new_n124), .c(new_n97), .o(new_n146));
  aoi022aa1n09x5               g051(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n147));
  aoai13aa1n03x5               g052(.a(new_n147), .b(new_n129), .c(new_n131), .d(new_n127), .o1(new_n148));
  oaib12aa1n09x5               g053(.a(new_n148), .b(\b[11] ), .c(new_n134), .out0(new_n149));
  aoi012aa1n03x5               g054(.a(new_n149), .b(new_n142), .c(new_n146), .o1(new_n150));
  xnrb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n03x5               g056(.a(\a[13] ), .b(\b[12] ), .c(new_n150), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand42aa1n03x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nor022aa1n08x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nand42aa1n08x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nano23aa1n06x5               g062(.a(new_n154), .b(new_n156), .c(new_n157), .d(new_n155), .out0(new_n158));
  aoai13aa1n03x5               g063(.a(new_n158), .b(new_n149), .c(new_n142), .d(new_n146), .o1(new_n159));
  oai012aa1n02x5               g064(.a(new_n157), .b(new_n156), .c(new_n154), .o1(new_n160));
  nor002aa1n04x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n159), .c(new_n160), .out0(\s[15] ));
  nanp02aa1n03x5               g069(.a(new_n159), .b(new_n160), .o1(new_n165));
  nor042aa1n02x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand42aa1n06x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n161), .c(new_n165), .d(new_n162), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(new_n165), .b(new_n163), .o1(new_n170));
  nona22aa1n02x4               g075(.a(new_n170), .b(new_n168), .c(new_n161), .out0(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n169), .o1(\s[16] ));
  nano23aa1n06x5               g077(.a(new_n161), .b(new_n166), .c(new_n167), .d(new_n162), .out0(new_n173));
  nand42aa1n04x5               g078(.a(new_n173), .b(new_n158), .o1(new_n174));
  nano32aa1n03x7               g079(.a(new_n174), .b(new_n145), .c(new_n124), .d(new_n97), .out0(new_n175));
  aoai13aa1n12x5               g080(.a(new_n175), .b(new_n123), .c(new_n120), .d(new_n109), .o1(new_n176));
  and002aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o(new_n177));
  oaoi13aa1n06x5               g082(.a(new_n161), .b(new_n157), .c(new_n154), .d(new_n156), .o1(new_n178));
  oai022aa1n03x5               g083(.a(new_n178), .b(new_n177), .c(\b[15] ), .d(\a[16] ), .o1(new_n179));
  aboi22aa1n12x5               g084(.a(new_n174), .b(new_n149), .c(new_n179), .d(new_n167), .out0(new_n180));
  nand02aa1d10x5               g085(.a(new_n176), .b(new_n180), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g087(.a(\a[18] ), .o1(new_n183));
  inv040aa1d32x5               g088(.a(\a[17] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\b[16] ), .o1(new_n185));
  oaoi03aa1n02x5               g090(.a(new_n184), .b(new_n185), .c(new_n181), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[17] ), .c(new_n183), .out0(\s[18] ));
  xroi22aa1d06x4               g092(.a(new_n184), .b(\b[16] ), .c(new_n183), .d(\b[17] ), .out0(new_n188));
  nand42aa1n02x5               g093(.a(new_n185), .b(new_n184), .o1(new_n189));
  oaoi03aa1n12x5               g094(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n190));
  nor042aa1n12x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nand22aa1n09x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n190), .c(new_n181), .d(new_n188), .o1(new_n195));
  aoi112aa1n02x5               g100(.a(new_n194), .b(new_n190), .c(new_n181), .d(new_n188), .o1(new_n196));
  norb02aa1n02x5               g101(.a(new_n195), .b(new_n196), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand22aa1n12x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  tech160nm_fioai012aa1n03p5x5 g106(.a(new_n195), .b(\b[18] ), .c(\a[19] ), .o1(new_n202));
  nanp02aa1n03x5               g107(.a(new_n202), .b(new_n201), .o1(new_n203));
  nona22aa1n02x4               g108(.a(new_n195), .b(new_n201), .c(new_n191), .out0(new_n204));
  nanp02aa1n03x5               g109(.a(new_n203), .b(new_n204), .o1(\s[20] ));
  nano23aa1n06x5               g110(.a(new_n191), .b(new_n199), .c(new_n200), .d(new_n192), .out0(new_n206));
  nanp02aa1n02x5               g111(.a(new_n188), .b(new_n206), .o1(new_n207));
  oai022aa1n04x5               g112(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n208));
  oaib12aa1n06x5               g113(.a(new_n208), .b(new_n183), .c(\b[17] ), .out0(new_n209));
  nona23aa1n09x5               g114(.a(new_n200), .b(new_n192), .c(new_n191), .d(new_n199), .out0(new_n210));
  aoi012aa1n06x5               g115(.a(new_n199), .b(new_n191), .c(new_n200), .o1(new_n211));
  oai012aa1n18x5               g116(.a(new_n211), .b(new_n210), .c(new_n209), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  aoai13aa1n04x5               g118(.a(new_n213), .b(new_n207), .c(new_n176), .d(new_n180), .o1(new_n214));
  xorb03aa1n02x5               g119(.a(new_n214), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  xorc02aa1n02x5               g121(.a(\a[21] ), .b(\b[20] ), .out0(new_n217));
  xorc02aa1n02x5               g122(.a(\a[22] ), .b(\b[21] ), .out0(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n216), .c(new_n214), .d(new_n217), .o1(new_n220));
  aoi112aa1n03x5               g125(.a(new_n216), .b(new_n219), .c(new_n214), .d(new_n217), .o1(new_n221));
  nanb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(\s[22] ));
  inv000aa1d42x5               g127(.a(\a[21] ), .o1(new_n223));
  inv040aa1d32x5               g128(.a(\a[22] ), .o1(new_n224));
  xroi22aa1d06x4               g129(.a(new_n223), .b(\b[20] ), .c(new_n224), .d(\b[21] ), .out0(new_n225));
  nanp03aa1n02x5               g130(.a(new_n225), .b(new_n188), .c(new_n206), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[21] ), .o1(new_n227));
  oao003aa1n02x5               g132(.a(new_n224), .b(new_n227), .c(new_n216), .carry(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n212), .c(new_n225), .o1(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n226), .c(new_n176), .d(new_n180), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .o1(new_n232));
  xorc02aa1n12x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[23] ), .b(\a[24] ), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n235));
  aoi112aa1n03x5               g140(.a(new_n232), .b(new_n234), .c(new_n230), .d(new_n233), .o1(new_n236));
  nanb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(\s[24] ));
  norb02aa1n06x4               g142(.a(new_n233), .b(new_n234), .out0(new_n238));
  nano22aa1n02x4               g143(.a(new_n207), .b(new_n238), .c(new_n225), .out0(new_n239));
  inv020aa1n03x5               g144(.a(new_n211), .o1(new_n240));
  aoai13aa1n06x5               g145(.a(new_n225), .b(new_n240), .c(new_n206), .d(new_n190), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n228), .o1(new_n242));
  inv000aa1n02x5               g147(.a(new_n238), .o1(new_n243));
  oai022aa1n02x5               g148(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n244));
  aob012aa1n02x5               g149(.a(new_n244), .b(\b[23] ), .c(\a[24] ), .out0(new_n245));
  aoai13aa1n12x5               g150(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n242), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aob012aa1n03x5               g152(.a(new_n247), .b(new_n181), .c(new_n239), .out0(new_n248));
  xorb03aa1n02x5               g153(.a(new_n248), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g154(.a(\b[24] ), .b(\a[25] ), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[25] ), .b(\b[24] ), .out0(new_n251));
  nor002aa1n03x5               g156(.a(\b[25] ), .b(\a[26] ), .o1(new_n252));
  nand02aa1d06x5               g157(.a(\b[25] ), .b(\a[26] ), .o1(new_n253));
  norb02aa1n09x5               g158(.a(new_n253), .b(new_n252), .out0(new_n254));
  inv040aa1n03x5               g159(.a(new_n254), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n250), .c(new_n248), .d(new_n251), .o1(new_n256));
  aoai13aa1n02x5               g161(.a(new_n251), .b(new_n246), .c(new_n181), .d(new_n239), .o1(new_n257));
  nona22aa1n02x4               g162(.a(new_n257), .b(new_n255), .c(new_n250), .out0(new_n258));
  nanp02aa1n03x5               g163(.a(new_n256), .b(new_n258), .o1(\s[26] ));
  norb02aa1n15x5               g164(.a(new_n251), .b(new_n255), .out0(new_n260));
  nano22aa1n06x5               g165(.a(new_n226), .b(new_n238), .c(new_n260), .out0(new_n261));
  nand02aa1d04x5               g166(.a(new_n181), .b(new_n261), .o1(new_n262));
  oai012aa1n02x5               g167(.a(new_n253), .b(new_n252), .c(new_n250), .o1(new_n263));
  aobi12aa1n12x5               g168(.a(new_n263), .b(new_n246), .c(new_n260), .out0(new_n264));
  xorc02aa1n02x5               g169(.a(\a[27] ), .b(\b[26] ), .out0(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n264), .c(new_n262), .out0(\s[27] ));
  nanp02aa1n06x5               g171(.a(new_n264), .b(new_n262), .o1(new_n267));
  norp02aa1n02x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  norp02aa1n02x5               g173(.a(\b[27] ), .b(\a[28] ), .o1(new_n269));
  nand42aa1n03x5               g174(.a(\b[27] ), .b(\a[28] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n270), .b(new_n269), .out0(new_n271));
  inv040aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n268), .c(new_n267), .d(new_n265), .o1(new_n273));
  aobi12aa1n09x5               g178(.a(new_n261), .b(new_n176), .c(new_n180), .out0(new_n274));
  aoai13aa1n02x7               g179(.a(new_n238), .b(new_n228), .c(new_n212), .d(new_n225), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n260), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n263), .b(new_n276), .c(new_n275), .d(new_n245), .o1(new_n277));
  oai012aa1n02x5               g182(.a(new_n265), .b(new_n277), .c(new_n274), .o1(new_n278));
  nona22aa1n02x5               g183(.a(new_n278), .b(new_n272), .c(new_n268), .out0(new_n279));
  nanp02aa1n03x5               g184(.a(new_n273), .b(new_n279), .o1(\s[28] ));
  norb02aa1n02x5               g185(.a(new_n265), .b(new_n272), .out0(new_n281));
  tech160nm_fioai012aa1n04x5   g186(.a(new_n281), .b(new_n277), .c(new_n274), .o1(new_n282));
  xorc02aa1n02x5               g187(.a(\a[29] ), .b(\b[28] ), .out0(new_n283));
  aoi012aa1n02x5               g188(.a(new_n269), .b(new_n268), .c(new_n270), .o1(new_n284));
  norb02aa1n02x5               g189(.a(new_n284), .b(new_n283), .out0(new_n285));
  nanp02aa1n03x5               g190(.a(new_n282), .b(new_n284), .o1(new_n286));
  aoi022aa1n02x7               g191(.a(new_n286), .b(new_n283), .c(new_n282), .d(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g193(.a(new_n265), .b(new_n283), .c(new_n271), .o(new_n289));
  tech160nm_fioai012aa1n05x5   g194(.a(new_n289), .b(new_n277), .c(new_n274), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[30] ), .b(\b[29] ), .out0(new_n291));
  oao003aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .carry(new_n292));
  norb02aa1n02x5               g197(.a(new_n292), .b(new_n291), .out0(new_n293));
  nanp02aa1n03x5               g198(.a(new_n290), .b(new_n292), .o1(new_n294));
  aoi022aa1n02x7               g199(.a(new_n294), .b(new_n291), .c(new_n290), .d(new_n293), .o1(\s[30] ));
  nanb02aa1n02x5               g200(.a(\b[30] ), .b(\a[31] ), .out0(new_n296));
  nanb02aa1n02x5               g201(.a(\a[31] ), .b(\b[30] ), .out0(new_n297));
  and003aa1n02x5               g202(.a(new_n281), .b(new_n291), .c(new_n283), .o(new_n298));
  oaih12aa1n02x5               g203(.a(new_n298), .b(new_n277), .c(new_n274), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[30] ), .b(\b[29] ), .c(new_n292), .carry(new_n300));
  aoi022aa1n02x7               g205(.a(new_n299), .b(new_n300), .c(new_n297), .d(new_n296), .o1(new_n301));
  aobi12aa1n06x5               g206(.a(new_n298), .b(new_n264), .c(new_n262), .out0(new_n302));
  nano32aa1n03x7               g207(.a(new_n302), .b(new_n300), .c(new_n296), .d(new_n297), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[31] ));
  xnrb03aa1n02x5               g209(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g210(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n306));
  xorb03aa1n02x5               g211(.a(new_n306), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g212(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g213(.a(new_n140), .o1(new_n309));
  aoi012aa1n03x5               g214(.a(new_n112), .b(new_n109), .c(new_n113), .o1(new_n310));
  xnrc02aa1n02x5               g215(.a(new_n310), .b(new_n309), .out0(\s[6] ));
  aob012aa1n03x5               g216(.a(new_n115), .b(new_n310), .c(new_n309), .out0(new_n312));
  xnbna2aa1n03x5               g217(.a(new_n312), .b(new_n121), .c(new_n111), .out0(\s[7] ));
  oaoi03aa1n03x5               g218(.a(\a[7] ), .b(\b[6] ), .c(new_n312), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g220(.a(new_n142), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


