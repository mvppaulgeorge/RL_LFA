// Benchmark "adder" written by ABC on Thu Jul 18 13:04:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n317, new_n319, new_n320,
    new_n321, new_n323, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1n02x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nor022aa1n16x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  norp02aa1n06x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  oai012aa1n02x7               g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n12x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nor022aa1n03x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  tech160nm_fioai012aa1n05x5   g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  nand42aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n99), .b(new_n107), .c(new_n101), .d(new_n100), .out0(new_n108));
  oaih12aa1n06x5               g013(.a(new_n102), .b(new_n108), .c(new_n106), .o1(new_n109));
  nor022aa1n12x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nand22aa1n06x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor022aa1n16x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  xnrc02aa1n12x5               g019(.a(\b[7] ), .b(\a[8] ), .out0(new_n115));
  xnrc02aa1n12x5               g020(.a(\b[6] ), .b(\a[7] ), .out0(new_n116));
  nor043aa1n03x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  norp02aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  tech160nm_fioai012aa1n03p5x5 g024(.a(new_n118), .b(new_n115), .c(new_n119), .o1(new_n120));
  tech160nm_fiaoi012aa1n05x5   g025(.a(new_n110), .b(new_n112), .c(new_n111), .o1(new_n121));
  oai013aa1n09x5               g026(.a(new_n120), .b(new_n121), .c(new_n115), .d(new_n116), .o1(new_n122));
  tech160nm_fixorc02aa1n05x5   g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  aoai13aa1n02x5               g028(.a(new_n123), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n124));
  nor042aa1n04x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nand42aa1n08x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  norb02aa1n15x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n127), .b(new_n124), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g033(.a(new_n127), .o1(new_n129));
  aoi012aa1n06x5               g034(.a(new_n125), .b(new_n97), .c(new_n126), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n129), .c(new_n124), .d(new_n98), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n06x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1n08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nano22aa1n02x4               g039(.a(new_n133), .b(new_n131), .c(new_n134), .out0(new_n135));
  nor042aa1n04x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand42aa1n08x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aoi012aa1n02x5               g043(.a(new_n133), .b(new_n131), .c(new_n134), .o1(new_n139));
  nona22aa1n02x4               g044(.a(new_n137), .b(new_n136), .c(new_n133), .out0(new_n140));
  oai022aa1n02x5               g045(.a(new_n135), .b(new_n140), .c(new_n139), .d(new_n138), .o1(\s[12] ));
  aoi012aa1n12x5               g046(.a(new_n122), .b(new_n109), .c(new_n117), .o1(new_n142));
  nano23aa1n06x5               g047(.a(new_n133), .b(new_n136), .c(new_n137), .d(new_n134), .out0(new_n143));
  nand23aa1n04x5               g048(.a(new_n143), .b(new_n123), .c(new_n127), .o1(new_n144));
  nona23aa1n02x4               g049(.a(new_n137), .b(new_n134), .c(new_n133), .d(new_n136), .out0(new_n145));
  oa0012aa1n03x5               g050(.a(new_n137), .b(new_n136), .c(new_n133), .o(new_n146));
  inv040aa1n03x5               g051(.a(new_n146), .o1(new_n147));
  oai012aa1n02x5               g052(.a(new_n147), .b(new_n145), .c(new_n130), .o1(new_n148));
  oabi12aa1n02x5               g053(.a(new_n148), .b(new_n142), .c(new_n144), .out0(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n04x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  tech160nm_finand02aa1n03p5x5 g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  aoi012aa1n03x5               g057(.a(new_n151), .b(new_n149), .c(new_n152), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  tech160nm_finand02aa1n03p5x5 g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nor042aa1n02x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nano23aa1n09x5               g061(.a(new_n151), .b(new_n156), .c(new_n155), .d(new_n152), .out0(new_n157));
  oai022aa1n02x5               g062(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n158));
  aoi022aa1n02x5               g063(.a(new_n148), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n159));
  nona22aa1n09x5               g064(.a(new_n157), .b(new_n142), .c(new_n144), .out0(new_n160));
  nor002aa1n16x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nand42aa1d28x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(new_n161), .b(new_n162), .out0(new_n163));
  xobna2aa1n03x5               g068(.a(new_n163), .b(new_n160), .c(new_n159), .out0(\s[15] ));
  inv000aa1d42x5               g069(.a(new_n161), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n163), .c(new_n160), .d(new_n159), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor002aa1n04x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  nand42aa1n16x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nano23aa1d15x5               g074(.a(new_n161), .b(new_n168), .c(new_n169), .d(new_n162), .out0(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  nano22aa1d15x5               g076(.a(new_n144), .b(new_n157), .c(new_n170), .out0(new_n172));
  aoai13aa1n12x5               g077(.a(new_n172), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n173));
  oai012aa1n02x7               g078(.a(new_n169), .b(new_n168), .c(new_n161), .o1(new_n174));
  oai112aa1n06x5               g079(.a(new_n173), .b(new_n174), .c(new_n159), .d(new_n171), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g081(.a(\a[18] ), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n173), .o1(new_n178));
  inv040aa1n02x5               g083(.a(new_n130), .o1(new_n179));
  aoai13aa1n04x5               g084(.a(new_n157), .b(new_n146), .c(new_n143), .d(new_n179), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n155), .b(new_n156), .c(new_n151), .o1(new_n181));
  aoai13aa1n12x5               g086(.a(new_n174), .b(new_n171), .c(new_n180), .d(new_n181), .o1(new_n182));
  norp02aa1n02x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  xorc02aa1n02x5               g088(.a(\a[17] ), .b(\b[16] ), .out0(new_n184));
  oaoi13aa1n02x5               g089(.a(new_n183), .b(new_n184), .c(new_n178), .d(new_n182), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n177), .out0(\s[18] ));
  inv000aa1d42x5               g091(.a(new_n182), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\a[17] ), .o1(new_n188));
  xroi22aa1d06x4               g093(.a(new_n188), .b(\b[16] ), .c(new_n177), .d(\b[17] ), .out0(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[17] ), .o1(new_n191));
  oai022aa1d24x5               g096(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n192));
  oaib12aa1n09x5               g097(.a(new_n192), .b(new_n191), .c(\a[18] ), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n190), .c(new_n187), .d(new_n173), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n12x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanp02aa1n04x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nor002aa1n06x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1n06x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  aoai13aa1n02x5               g106(.a(new_n201), .b(new_n197), .c(new_n194), .d(new_n198), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n142), .o1(new_n203));
  aoai13aa1n02x5               g108(.a(new_n189), .b(new_n182), .c(new_n203), .d(new_n172), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n197), .b(new_n198), .out0(new_n205));
  norb03aa1n02x5               g110(.a(new_n200), .b(new_n197), .c(new_n199), .out0(new_n206));
  aoai13aa1n02x5               g111(.a(new_n206), .b(new_n205), .c(new_n204), .d(new_n193), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n202), .b(new_n207), .o1(\s[20] ));
  nano23aa1n09x5               g113(.a(new_n197), .b(new_n199), .c(new_n200), .d(new_n198), .out0(new_n209));
  nand22aa1n12x5               g114(.a(new_n189), .b(new_n209), .o1(new_n210));
  nona23aa1n09x5               g115(.a(new_n200), .b(new_n198), .c(new_n197), .d(new_n199), .out0(new_n211));
  oai012aa1n12x5               g116(.a(new_n200), .b(new_n199), .c(new_n197), .o1(new_n212));
  oai012aa1d24x5               g117(.a(new_n212), .b(new_n211), .c(new_n193), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  aoai13aa1n04x5               g119(.a(new_n214), .b(new_n210), .c(new_n187), .d(new_n173), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xorc02aa1n12x5               g123(.a(\a[22] ), .b(\b[21] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n02x5               g125(.a(new_n220), .b(new_n217), .c(new_n215), .d(new_n218), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n210), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n218), .b(new_n213), .c(new_n175), .d(new_n222), .o1(new_n223));
  nona22aa1n03x5               g128(.a(new_n223), .b(new_n220), .c(new_n217), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n221), .b(new_n224), .o1(\s[22] ));
  nano32aa1n03x7               g130(.a(new_n190), .b(new_n219), .c(new_n209), .d(new_n218), .out0(new_n226));
  inv000aa1n02x5               g131(.a(new_n226), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv040aa1d32x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(\b[21] ), .o1(new_n231));
  oao003aa1n02x5               g136(.a(new_n229), .b(new_n231), .c(new_n217), .carry(new_n232));
  aoi012aa1d18x5               g137(.a(new_n232), .b(new_n213), .c(new_n230), .o1(new_n233));
  aoai13aa1n04x5               g138(.a(new_n233), .b(new_n227), .c(new_n187), .d(new_n173), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  xorc02aa1n06x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  xnrc02aa1n02x5               g142(.a(\b[23] ), .b(\a[24] ), .out0(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n236), .c(new_n234), .d(new_n237), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n233), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n237), .b(new_n240), .c(new_n175), .d(new_n226), .o1(new_n241));
  nona22aa1n03x5               g146(.a(new_n241), .b(new_n238), .c(new_n236), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n239), .b(new_n242), .o1(\s[24] ));
  norb02aa1n03x5               g148(.a(new_n237), .b(new_n238), .out0(new_n244));
  nano22aa1n03x7               g149(.a(new_n210), .b(new_n244), .c(new_n230), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n182), .c(new_n203), .d(new_n172), .o1(new_n246));
  inv030aa1n02x5               g151(.a(new_n193), .o1(new_n247));
  inv000aa1n02x5               g152(.a(new_n212), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n230), .b(new_n248), .c(new_n209), .d(new_n247), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n232), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n244), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\a[24] ), .o1(new_n252));
  inv000aa1d42x5               g157(.a(\b[23] ), .o1(new_n253));
  oao003aa1n02x5               g158(.a(new_n252), .b(new_n253), .c(new_n236), .carry(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  aoai13aa1n12x5               g160(.a(new_n255), .b(new_n251), .c(new_n249), .d(new_n250), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  tech160nm_fixorc02aa1n05x5   g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  xnbna2aa1n03x5               g163(.a(new_n258), .b(new_n246), .c(new_n257), .out0(\s[25] ));
  nand02aa1n03x5               g164(.a(new_n246), .b(new_n257), .o1(new_n260));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  norp02aa1n02x5               g166(.a(\b[25] ), .b(\a[26] ), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(\b[25] ), .b(\a[26] ), .o1(new_n263));
  norb02aa1n02x5               g168(.a(new_n263), .b(new_n262), .out0(new_n264));
  inv040aa1n03x5               g169(.a(new_n264), .o1(new_n265));
  aoai13aa1n02x5               g170(.a(new_n265), .b(new_n261), .c(new_n260), .d(new_n258), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n258), .b(new_n256), .c(new_n175), .d(new_n245), .o1(new_n267));
  nona22aa1n03x5               g172(.a(new_n267), .b(new_n265), .c(new_n261), .out0(new_n268));
  nanp02aa1n03x5               g173(.a(new_n266), .b(new_n268), .o1(\s[26] ));
  norb02aa1n03x5               g174(.a(new_n258), .b(new_n265), .out0(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  nano23aa1d15x5               g176(.a(new_n210), .b(new_n271), .c(new_n244), .d(new_n230), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n182), .c(new_n203), .d(new_n172), .o1(new_n273));
  oai012aa1n02x5               g178(.a(new_n263), .b(new_n262), .c(new_n261), .o1(new_n274));
  aobi12aa1n12x5               g179(.a(new_n274), .b(new_n256), .c(new_n270), .out0(new_n275));
  xorc02aa1n02x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n273), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  inv040aa1n03x5               g183(.a(new_n278), .o1(new_n279));
  aoai13aa1n02x5               g184(.a(new_n244), .b(new_n232), .c(new_n213), .d(new_n230), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n274), .b(new_n271), .c(new_n280), .d(new_n255), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n276), .b(new_n281), .c(new_n175), .d(new_n272), .o1(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n283), .b(new_n282), .c(new_n279), .o1(new_n284));
  aobi12aa1n02x7               g189(.a(new_n276), .b(new_n275), .c(new_n273), .out0(new_n285));
  nano22aa1n02x4               g190(.a(new_n285), .b(new_n279), .c(new_n283), .out0(new_n286));
  norp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[28] ));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  norb02aa1n02x5               g193(.a(new_n276), .b(new_n283), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n281), .c(new_n175), .d(new_n272), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n279), .carry(new_n291));
  aoi012aa1n02x7               g196(.a(new_n288), .b(new_n290), .c(new_n291), .o1(new_n292));
  aobi12aa1n02x7               g197(.a(new_n289), .b(new_n275), .c(new_n273), .out0(new_n293));
  nano22aa1n02x4               g198(.a(new_n293), .b(new_n288), .c(new_n291), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g201(.a(\b[29] ), .b(\a[30] ), .out0(new_n297));
  norb03aa1n02x5               g202(.a(new_n276), .b(new_n288), .c(new_n283), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n281), .c(new_n175), .d(new_n272), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n297), .b(new_n299), .c(new_n300), .o1(new_n301));
  aobi12aa1n02x7               g206(.a(new_n298), .b(new_n275), .c(new_n273), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n297), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[30] ));
  norb02aa1n02x5               g209(.a(new_n298), .b(new_n297), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n281), .c(new_n175), .d(new_n272), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  aobi12aa1n02x7               g214(.a(new_n305), .b(new_n275), .c(new_n273), .out0(new_n310));
  nano22aa1n02x4               g215(.a(new_n310), .b(new_n307), .c(new_n308), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[31] ));
  xnrb03aa1n02x5               g217(.a(new_n106), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g218(.a(\a[3] ), .b(\b[2] ), .c(new_n106), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g220(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g221(.a(new_n112), .b(new_n109), .c(new_n113), .o1(new_n317));
  xnrb03aa1n02x5               g222(.a(new_n317), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g223(.a(new_n110), .b(new_n111), .out0(new_n319));
  oaoi13aa1n02x5               g224(.a(new_n116), .b(new_n121), .c(new_n317), .d(new_n319), .o1(new_n320));
  oai112aa1n02x5               g225(.a(new_n121), .b(new_n116), .c(new_n317), .d(new_n319), .o1(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(\s[7] ));
  oabi12aa1n02x5               g227(.a(new_n115), .b(\a[7] ), .c(\b[6] ), .out0(new_n323));
  oai012aa1n02x5               g228(.a(new_n115), .b(new_n320), .c(new_n119), .o1(new_n324));
  oai012aa1n02x5               g229(.a(new_n324), .b(new_n320), .c(new_n323), .o1(\s[8] ));
  xnrc02aa1n02x5               g230(.a(new_n142), .b(new_n123), .out0(\s[9] ));
endmodule


