// Benchmark "adder" written by ABC on Thu Jul 18 10:16:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n316, new_n317, new_n318, new_n320,
    new_n322;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor042aa1n04x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  norp02aa1n04x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n101), .b(new_n104), .c(new_n103), .d(new_n102), .out0(new_n105));
  nor002aa1n03x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nand42aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  aoi012aa1n02x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  oai012aa1n02x5               g014(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n110));
  tech160nm_fioai012aa1n04x5   g015(.a(new_n110), .b(new_n105), .c(new_n109), .o1(new_n111));
  inv000aa1n02x5               g016(.a(new_n111), .o1(new_n112));
  norp02aa1n02x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand02aa1n02x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  tech160nm_fiaoi012aa1n05x5   g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nor022aa1n04x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  nand42aa1n02x5               g022(.a(\b[3] ), .b(\a[4] ), .o1(new_n118));
  nor022aa1n16x5               g023(.a(\b[2] ), .b(\a[3] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  nona23aa1n03x5               g025(.a(new_n120), .b(new_n118), .c(new_n117), .d(new_n119), .out0(new_n121));
  oai012aa1n02x5               g026(.a(new_n118), .b(new_n119), .c(new_n117), .o1(new_n122));
  tech160nm_fioai012aa1n05x5   g027(.a(new_n122), .b(new_n121), .c(new_n116), .o1(new_n123));
  nanb02aa1n02x5               g028(.a(new_n106), .b(new_n108), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .out0(new_n125));
  nor003aa1n03x5               g030(.a(new_n105), .b(new_n124), .c(new_n125), .o1(new_n126));
  nanp02aa1n03x5               g031(.a(new_n123), .b(new_n126), .o1(new_n127));
  nanp02aa1n06x5               g032(.a(new_n127), .b(new_n112), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  tech160nm_fiaoi012aa1n05x5   g034(.a(new_n100), .b(new_n128), .c(new_n129), .o1(new_n130));
  xnrc02aa1n02x5               g035(.a(new_n130), .b(new_n99), .out0(\s[10] ));
  nanp02aa1n03x5               g036(.a(new_n130), .b(new_n99), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb02aa1n12x5               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n132), .c(new_n98), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n98), .o1(new_n137));
  nona22aa1n02x4               g042(.a(new_n132), .b(new_n135), .c(new_n137), .out0(new_n138));
  nor002aa1n20x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand22aa1n02x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n06x4               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  nona22aa1n02x4               g046(.a(new_n138), .b(new_n141), .c(new_n133), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n133), .o1(new_n143));
  nanb02aa1n06x5               g048(.a(new_n139), .b(new_n140), .out0(new_n144));
  tech160nm_fiaoi012aa1n02p5x5 g049(.a(new_n144), .b(new_n138), .c(new_n143), .o1(new_n145));
  norb02aa1n02x7               g050(.a(new_n142), .b(new_n145), .out0(\s[12] ));
  nano23aa1n02x5               g051(.a(new_n97), .b(new_n100), .c(new_n129), .d(new_n98), .out0(new_n147));
  nona22aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n135), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n139), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n133), .b(new_n140), .o1(new_n150));
  oai022aa1n02x5               g055(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n151));
  nano23aa1n02x4               g056(.a(new_n144), .b(new_n135), .c(new_n151), .d(new_n98), .out0(new_n152));
  nano22aa1n03x7               g057(.a(new_n152), .b(new_n149), .c(new_n150), .out0(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n148), .c(new_n127), .d(new_n112), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1n06x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n156), .b(new_n154), .c(new_n157), .o1(new_n158));
  nor042aa1n04x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nand02aa1d10x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  xnrc02aa1n02x5               g066(.a(new_n158), .b(new_n161), .out0(\s[14] ));
  nor002aa1n03x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nand42aa1n06x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  nano23aa1n09x5               g070(.a(new_n156), .b(new_n159), .c(new_n160), .d(new_n157), .out0(new_n166));
  aoi012aa1d18x5               g071(.a(new_n159), .b(new_n156), .c(new_n160), .o1(new_n167));
  inv000aa1n02x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n06x5               g073(.a(new_n165), .b(new_n168), .c(new_n154), .d(new_n166), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n165), .b(new_n168), .c(new_n154), .d(new_n166), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[15] ));
  nor022aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  nona22aa1n03x5               g079(.a(new_n169), .b(new_n174), .c(new_n163), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n174), .o1(new_n176));
  oaoi13aa1n04x5               g081(.a(new_n176), .b(new_n169), .c(\a[15] ), .d(\b[14] ), .o1(new_n177));
  norb02aa1n03x4               g082(.a(new_n175), .b(new_n177), .out0(\s[16] ));
  norb02aa1n02x5               g083(.a(new_n134), .b(new_n133), .out0(new_n179));
  nor002aa1n02x5               g084(.a(new_n100), .b(new_n97), .o1(new_n180));
  nona23aa1n03x5               g085(.a(new_n141), .b(new_n179), .c(new_n180), .d(new_n137), .out0(new_n181));
  nand23aa1n03x5               g086(.a(new_n181), .b(new_n149), .c(new_n150), .o1(new_n182));
  nano23aa1n09x5               g087(.a(new_n163), .b(new_n172), .c(new_n173), .d(new_n164), .out0(new_n183));
  nand02aa1d04x5               g088(.a(new_n183), .b(new_n166), .o1(new_n184));
  inv020aa1n02x5               g089(.a(new_n184), .o1(new_n185));
  oai012aa1n02x5               g090(.a(new_n173), .b(new_n172), .c(new_n163), .o1(new_n186));
  aob012aa1n06x5               g091(.a(new_n186), .b(new_n183), .c(new_n168), .out0(new_n187));
  aoi012aa1d18x5               g092(.a(new_n187), .b(new_n182), .c(new_n185), .o1(new_n188));
  nor042aa1n06x5               g093(.a(new_n148), .b(new_n184), .o1(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n111), .c(new_n123), .d(new_n126), .o1(new_n190));
  nanp02aa1n09x5               g095(.a(new_n188), .b(new_n190), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g097(.a(\a[18] ), .o1(new_n193));
  inv040aa1d28x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  oaoi03aa1n03x5               g100(.a(new_n194), .b(new_n195), .c(new_n191), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  xroi22aa1d06x4               g102(.a(new_n194), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  norp02aa1n02x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nand22aa1n06x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  aoi013aa1n06x4               g106(.a(new_n200), .b(new_n201), .c(new_n194), .d(new_n195), .o1(new_n202));
  aoai13aa1n04x5               g107(.a(new_n202), .b(new_n199), .c(new_n188), .d(new_n190), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand02aa1d28x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nor002aa1d32x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand42aa1n20x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi112aa1n02x5               g115(.a(new_n206), .b(new_n210), .c(new_n203), .d(new_n207), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n210), .b(new_n206), .c(new_n203), .d(new_n207), .o1(new_n212));
  norb02aa1n02x7               g117(.a(new_n212), .b(new_n211), .out0(\s[20] ));
  nano23aa1n09x5               g118(.a(new_n206), .b(new_n208), .c(new_n209), .d(new_n207), .out0(new_n214));
  nand02aa1d04x5               g119(.a(new_n198), .b(new_n214), .o1(new_n215));
  nona23aa1n09x5               g120(.a(new_n209), .b(new_n207), .c(new_n206), .d(new_n208), .out0(new_n216));
  oai012aa1n04x7               g121(.a(new_n209), .b(new_n208), .c(new_n206), .o1(new_n217));
  oai012aa1n12x5               g122(.a(new_n217), .b(new_n216), .c(new_n202), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n04x5               g124(.a(new_n219), .b(new_n215), .c(new_n188), .d(new_n190), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n04x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[21] ), .b(\b[20] ), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[22] ), .b(\b[21] ), .out0(new_n224));
  aoi112aa1n03x5               g129(.a(new_n222), .b(new_n224), .c(new_n220), .d(new_n223), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n224), .b(new_n222), .c(new_n220), .d(new_n223), .o1(new_n226));
  norb02aa1n02x7               g131(.a(new_n226), .b(new_n225), .out0(\s[22] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv040aa1d32x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  nand23aa1n06x5               g135(.a(new_n230), .b(new_n198), .c(new_n214), .o1(new_n231));
  nona22aa1n02x4               g136(.a(new_n201), .b(\b[16] ), .c(\a[17] ), .out0(new_n232));
  oaib12aa1n06x5               g137(.a(new_n232), .b(\b[17] ), .c(new_n193), .out0(new_n233));
  inv000aa1n02x5               g138(.a(new_n217), .o1(new_n234));
  aoai13aa1n06x5               g139(.a(new_n230), .b(new_n234), .c(new_n214), .d(new_n233), .o1(new_n235));
  inv000aa1d42x5               g140(.a(\b[21] ), .o1(new_n236));
  oao003aa1n02x5               g141(.a(new_n229), .b(new_n236), .c(new_n222), .carry(new_n237));
  inv030aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  nanp02aa1n02x5               g143(.a(new_n235), .b(new_n238), .o1(new_n239));
  inv000aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  aoai13aa1n04x5               g145(.a(new_n240), .b(new_n231), .c(new_n188), .d(new_n190), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  tech160nm_fixorc02aa1n05x5   g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  xorc02aa1n03x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoi112aa1n02x5               g150(.a(new_n243), .b(new_n245), .c(new_n241), .d(new_n244), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n247));
  norb02aa1n02x7               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  and002aa1n02x5               g153(.a(new_n245), .b(new_n244), .o(new_n249));
  nanb03aa1n03x5               g154(.a(new_n215), .b(new_n249), .c(new_n230), .out0(new_n250));
  inv000aa1n02x5               g155(.a(new_n249), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  oai022aa1n02x5               g157(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n253), .b(new_n252), .o1(new_n254));
  aoai13aa1n12x5               g159(.a(new_n254), .b(new_n251), .c(new_n235), .d(new_n238), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n04x5               g161(.a(new_n256), .b(new_n250), .c(new_n188), .d(new_n190), .o1(new_n257));
  xorb03aa1n02x5               g162(.a(new_n257), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  xorc02aa1n02x5               g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  xorc02aa1n02x5               g165(.a(\a[26] ), .b(\b[25] ), .out0(new_n261));
  aoi112aa1n02x5               g166(.a(new_n259), .b(new_n261), .c(new_n257), .d(new_n260), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n261), .b(new_n259), .c(new_n257), .d(new_n260), .o1(new_n263));
  norb02aa1n02x7               g168(.a(new_n263), .b(new_n262), .out0(\s[26] ));
  oabi12aa1n03x5               g169(.a(new_n187), .b(new_n153), .c(new_n184), .out0(new_n265));
  and002aa1n12x5               g170(.a(new_n261), .b(new_n260), .o(new_n266));
  nano22aa1n03x7               g171(.a(new_n231), .b(new_n249), .c(new_n266), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n265), .c(new_n128), .d(new_n189), .o1(new_n268));
  oai022aa1n02x5               g173(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n269));
  aob012aa1n02x5               g174(.a(new_n269), .b(\b[25] ), .c(\a[26] ), .out0(new_n270));
  aobi12aa1n12x5               g175(.a(new_n270), .b(new_n255), .c(new_n266), .out0(new_n271));
  xorc02aa1n02x5               g176(.a(\a[27] ), .b(\b[26] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n268), .out0(\s[27] ));
  nor042aa1n03x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n274), .o1(new_n275));
  aobi12aa1n02x7               g180(.a(new_n272), .b(new_n271), .c(new_n268), .out0(new_n276));
  xnrc02aa1n02x5               g181(.a(\b[27] ), .b(\a[28] ), .out0(new_n277));
  nano22aa1n03x5               g182(.a(new_n276), .b(new_n275), .c(new_n277), .out0(new_n278));
  inv020aa1n02x5               g183(.a(new_n267), .o1(new_n279));
  aoi012aa1n06x5               g184(.a(new_n279), .b(new_n188), .c(new_n190), .o1(new_n280));
  aoai13aa1n02x7               g185(.a(new_n249), .b(new_n237), .c(new_n218), .d(new_n230), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n266), .o1(new_n282));
  aoai13aa1n04x5               g187(.a(new_n270), .b(new_n282), .c(new_n281), .d(new_n254), .o1(new_n283));
  oaih12aa1n02x5               g188(.a(new_n272), .b(new_n283), .c(new_n280), .o1(new_n284));
  tech160nm_fiaoi012aa1n03p5x5 g189(.a(new_n277), .b(new_n284), .c(new_n275), .o1(new_n285));
  norp02aa1n03x5               g190(.a(new_n285), .b(new_n278), .o1(\s[28] ));
  norb02aa1n02x5               g191(.a(new_n272), .b(new_n277), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n283), .c(new_n280), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n275), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[28] ), .b(\a[29] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  aobi12aa1n02x7               g196(.a(new_n287), .b(new_n271), .c(new_n268), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g200(.a(new_n272), .b(new_n290), .c(new_n277), .out0(new_n296));
  oaih12aa1n02x5               g201(.a(new_n296), .b(new_n283), .c(new_n280), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[29] ), .b(\a[30] ), .out0(new_n299));
  tech160nm_fiaoi012aa1n03p5x5 g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n296), .b(new_n271), .c(new_n268), .out0(new_n301));
  nano22aa1n02x4               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[30] ));
  norb02aa1n02x5               g208(.a(new_n296), .b(new_n299), .out0(new_n304));
  aobi12aa1n02x7               g209(.a(new_n304), .b(new_n271), .c(new_n268), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  nano22aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n307), .out0(new_n308));
  oaih12aa1n02x5               g213(.a(new_n304), .b(new_n283), .c(new_n280), .o1(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n307), .b(new_n309), .c(new_n306), .o1(new_n310));
  norp02aa1n03x5               g215(.a(new_n310), .b(new_n308), .o1(\s[31] ));
  xnrb03aa1n02x5               g216(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g217(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g219(.a(new_n123), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi13aa1n02x5               g220(.a(new_n125), .b(new_n122), .c(new_n121), .d(new_n116), .o1(new_n316));
  oai012aa1n02x5               g221(.a(new_n124), .b(new_n316), .c(new_n107), .o1(new_n317));
  orn003aa1n02x5               g222(.a(new_n316), .b(new_n107), .c(new_n124), .o(new_n318));
  nanp02aa1n02x5               g223(.a(new_n318), .b(new_n317), .o1(\s[6] ));
  oai013aa1n02x4               g224(.a(new_n108), .b(new_n316), .c(new_n106), .d(new_n107), .o1(new_n320));
  xnrb03aa1n02x5               g225(.a(new_n320), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g226(.a(\a[7] ), .b(\b[6] ), .c(new_n320), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g228(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


