// Benchmark "adder" written by ABC on Wed Jul 17 21:50:14 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n324,
    new_n327, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1n06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor042aa1n06x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor042aa1n04x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nand42aa1n20x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano23aa1n02x4               g009(.a(new_n101), .b(new_n103), .c(new_n104), .d(new_n102), .out0(new_n105));
  inv000aa1d42x5               g010(.a(\a[2] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[1] ), .o1(new_n107));
  nand22aa1n03x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  oao003aa1n02x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .carry(new_n109));
  aoi012aa1n02x5               g014(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n110));
  aobi12aa1n06x5               g015(.a(new_n110), .b(new_n105), .c(new_n109), .out0(new_n111));
  nor002aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1d28x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n08x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand02aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  nona22aa1n03x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\a[5] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[4] ), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  tech160nm_fiao0012aa1n02p5x5 g028(.a(new_n112), .b(new_n114), .c(new_n113), .o(new_n124));
  aoi012aa1n06x5               g029(.a(new_n124), .b(new_n116), .c(new_n123), .o1(new_n125));
  oai012aa1n03x5               g030(.a(new_n125), .b(new_n111), .c(new_n119), .o1(new_n126));
  tech160nm_finand02aa1n03p5x5 g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  tech160nm_fiaoi012aa1n05x5   g032(.a(new_n100), .b(new_n126), .c(new_n127), .o1(new_n128));
  xnrc02aa1n02x5               g033(.a(new_n128), .b(new_n99), .out0(\s[10] ));
  nanp02aa1n06x5               g034(.a(new_n128), .b(new_n99), .o1(new_n130));
  nor002aa1d32x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanp02aa1n06x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  xobna2aa1n03x5               g038(.a(new_n133), .b(new_n130), .c(new_n98), .out0(\s[11] ));
  nor002aa1d32x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nand42aa1n04x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  aoi113aa1n02x5               g042(.a(new_n137), .b(new_n131), .c(new_n130), .d(new_n133), .e(new_n98), .o1(new_n138));
  inv040aa1n03x5               g043(.a(new_n131), .o1(new_n139));
  nanp03aa1n02x5               g044(.a(new_n130), .b(new_n98), .c(new_n133), .o1(new_n140));
  aobi12aa1n02x7               g045(.a(new_n137), .b(new_n140), .c(new_n139), .out0(new_n141));
  nor002aa1n02x5               g046(.a(new_n141), .b(new_n138), .o1(\s[12] ));
  nona23aa1n02x4               g047(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n143));
  oaoi03aa1n02x5               g048(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n144));
  oaih12aa1n02x5               g049(.a(new_n110), .b(new_n143), .c(new_n144), .o1(new_n145));
  nona23aa1n03x5               g050(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n146));
  nor003aa1n02x5               g051(.a(new_n146), .b(new_n117), .c(new_n118), .o1(new_n147));
  nanp02aa1n03x5               g052(.a(new_n145), .b(new_n147), .o1(new_n148));
  nona23aa1d18x5               g053(.a(new_n136), .b(new_n132), .c(new_n131), .d(new_n135), .out0(new_n149));
  tech160nm_fioai012aa1n05x5   g054(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n150));
  oaoi03aa1n09x5               g055(.a(\a[12] ), .b(\b[11] ), .c(new_n139), .o1(new_n151));
  oabi12aa1n12x5               g056(.a(new_n151), .b(new_n149), .c(new_n150), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  nano23aa1n09x5               g058(.a(new_n131), .b(new_n135), .c(new_n136), .d(new_n132), .out0(new_n154));
  nano23aa1n02x5               g059(.a(new_n97), .b(new_n100), .c(new_n127), .d(new_n98), .out0(new_n155));
  nand02aa1n02x5               g060(.a(new_n155), .b(new_n154), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n153), .b(new_n156), .c(new_n148), .d(new_n125), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g063(.a(\a[14] ), .o1(new_n159));
  nor042aa1n03x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  xnrc02aa1n12x5               g065(.a(\b[12] ), .b(\a[13] ), .out0(new_n161));
  aoib12aa1n02x5               g066(.a(new_n160), .b(new_n157), .c(new_n161), .out0(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[13] ), .c(new_n159), .out0(\s[14] ));
  nor042aa1d18x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand42aa1d28x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  tech160nm_fixnrc02aa1n02p5x5 g072(.a(\b[13] ), .b(\a[14] ), .out0(new_n168));
  nor042aa1n04x5               g073(.a(new_n168), .b(new_n161), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\b[13] ), .o1(new_n170));
  tech160nm_fioaoi03aa1n03p5x5 g075(.a(new_n159), .b(new_n170), .c(new_n160), .o1(new_n171));
  inv000aa1n02x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n167), .b(new_n172), .c(new_n157), .d(new_n169), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n167), .b(new_n172), .c(new_n157), .d(new_n169), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(\s[15] ));
  inv000aa1d42x5               g080(.a(new_n164), .o1(new_n176));
  nor042aa1n09x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand42aa1d28x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n173), .c(new_n176), .out0(\s[16] ));
  inv000aa1n02x5               g086(.a(new_n125), .o1(new_n182));
  nano23aa1d15x5               g087(.a(new_n164), .b(new_n177), .c(new_n178), .d(new_n165), .out0(new_n183));
  nano22aa1n03x5               g088(.a(new_n156), .b(new_n169), .c(new_n183), .out0(new_n184));
  aoai13aa1n04x5               g089(.a(new_n184), .b(new_n182), .c(new_n145), .d(new_n147), .o1(new_n185));
  aoai13aa1n09x5               g090(.a(new_n183), .b(new_n172), .c(new_n152), .d(new_n169), .o1(new_n186));
  aoi012aa1d24x5               g091(.a(new_n177), .b(new_n164), .c(new_n178), .o1(new_n187));
  nand23aa1n06x5               g092(.a(new_n185), .b(new_n186), .c(new_n187), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g094(.a(\a[18] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\a[17] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[16] ), .o1(new_n192));
  oaoi03aa1n03x5               g097(.a(new_n191), .b(new_n192), .c(new_n188), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[17] ), .c(new_n190), .out0(\s[18] ));
  nona23aa1n03x5               g099(.a(new_n127), .b(new_n98), .c(new_n97), .d(new_n100), .out0(new_n195));
  nona23aa1d18x5               g100(.a(new_n169), .b(new_n183), .c(new_n195), .d(new_n149), .out0(new_n196));
  oaoi13aa1n12x5               g101(.a(new_n196), .b(new_n125), .c(new_n111), .d(new_n119), .o1(new_n197));
  inv000aa1d42x5               g102(.a(new_n183), .o1(new_n198));
  inv030aa1n04x5               g103(.a(new_n150), .o1(new_n199));
  aoai13aa1n04x5               g104(.a(new_n169), .b(new_n151), .c(new_n154), .d(new_n199), .o1(new_n200));
  aoai13aa1n09x5               g105(.a(new_n187), .b(new_n198), .c(new_n200), .d(new_n171), .o1(new_n201));
  xroi22aa1d06x4               g106(.a(new_n191), .b(\b[16] ), .c(new_n190), .d(\b[17] ), .out0(new_n202));
  tech160nm_fioai012aa1n03p5x5 g107(.a(new_n202), .b(new_n201), .c(new_n197), .o1(new_n203));
  oai022aa1n04x5               g108(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n204));
  oaib12aa1n09x5               g109(.a(new_n204), .b(new_n190), .c(\b[17] ), .out0(new_n205));
  nor042aa1d18x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand02aa1n06x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nanb02aa1n02x5               g112(.a(new_n206), .b(new_n207), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n203), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g116(.a(new_n206), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n208), .b(new_n203), .c(new_n205), .o1(new_n213));
  nor042aa1n06x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand02aa1d08x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nanb02aa1n02x5               g120(.a(new_n214), .b(new_n215), .out0(new_n216));
  nano22aa1n03x5               g121(.a(new_n213), .b(new_n212), .c(new_n216), .out0(new_n217));
  nanp02aa1n02x5               g122(.a(new_n192), .b(new_n191), .o1(new_n218));
  oaoi03aa1n02x5               g123(.a(\a[18] ), .b(\b[17] ), .c(new_n218), .o1(new_n219));
  oaoi13aa1n03x5               g124(.a(new_n219), .b(new_n202), .c(new_n201), .d(new_n197), .o1(new_n220));
  oaoi13aa1n02x7               g125(.a(new_n216), .b(new_n212), .c(new_n220), .d(new_n208), .o1(new_n221));
  norp02aa1n03x5               g126(.a(new_n221), .b(new_n217), .o1(\s[20] ));
  nano23aa1n09x5               g127(.a(new_n206), .b(new_n214), .c(new_n215), .d(new_n207), .out0(new_n223));
  nand02aa1n03x5               g128(.a(new_n202), .b(new_n223), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  tech160nm_fioai012aa1n03p5x5 g130(.a(new_n225), .b(new_n201), .c(new_n197), .o1(new_n226));
  nona23aa1n09x5               g131(.a(new_n215), .b(new_n207), .c(new_n206), .d(new_n214), .out0(new_n227));
  aoi012aa1d18x5               g132(.a(new_n214), .b(new_n206), .c(new_n215), .o1(new_n228));
  oai012aa1n18x5               g133(.a(new_n228), .b(new_n227), .c(new_n205), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  nor042aa1n06x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  nanp02aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n226), .c(new_n230), .out0(\s[21] ));
  inv000aa1d42x5               g139(.a(new_n231), .o1(new_n235));
  aobi12aa1n06x5               g140(.a(new_n233), .b(new_n226), .c(new_n230), .out0(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[21] ), .b(\a[22] ), .out0(new_n237));
  nano22aa1n02x4               g142(.a(new_n236), .b(new_n235), .c(new_n237), .out0(new_n238));
  aoai13aa1n03x5               g143(.a(new_n233), .b(new_n229), .c(new_n188), .d(new_n225), .o1(new_n239));
  tech160nm_fiaoi012aa1n02p5x5 g144(.a(new_n237), .b(new_n239), .c(new_n235), .o1(new_n240));
  norp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[22] ));
  nano22aa1n03x7               g146(.a(new_n237), .b(new_n235), .c(new_n232), .out0(new_n242));
  and003aa1n02x5               g147(.a(new_n202), .b(new_n242), .c(new_n223), .o(new_n243));
  tech160nm_fioai012aa1n03p5x5 g148(.a(new_n243), .b(new_n201), .c(new_n197), .o1(new_n244));
  oao003aa1n12x5               g149(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .carry(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  tech160nm_fiaoi012aa1n02p5x5 g151(.a(new_n246), .b(new_n229), .c(new_n242), .o1(new_n247));
  xnrc02aa1n12x5               g152(.a(\b[22] ), .b(\a[23] ), .out0(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  xnbna2aa1n03x5               g154(.a(new_n249), .b(new_n244), .c(new_n247), .out0(\s[23] ));
  nor042aa1n03x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  tech160nm_fiaoi012aa1n02p5x5 g157(.a(new_n248), .b(new_n244), .c(new_n247), .o1(new_n253));
  xnrc02aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n253), .b(new_n252), .c(new_n254), .out0(new_n255));
  inv030aa1n02x5               g160(.a(new_n247), .o1(new_n256));
  oaoi13aa1n03x5               g161(.a(new_n256), .b(new_n243), .c(new_n201), .d(new_n197), .o1(new_n257));
  oaoi13aa1n02x7               g162(.a(new_n254), .b(new_n252), .c(new_n257), .d(new_n248), .o1(new_n258));
  norp02aa1n03x5               g163(.a(new_n258), .b(new_n255), .o1(\s[24] ));
  nor042aa1n02x5               g164(.a(new_n254), .b(new_n248), .o1(new_n260));
  nano22aa1n03x5               g165(.a(new_n224), .b(new_n242), .c(new_n260), .out0(new_n261));
  oaih12aa1n02x5               g166(.a(new_n261), .b(new_n201), .c(new_n197), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n228), .o1(new_n263));
  aoai13aa1n03x5               g168(.a(new_n242), .b(new_n263), .c(new_n223), .d(new_n219), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n260), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n252), .carry(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n265), .c(new_n264), .d(new_n245), .o1(new_n267));
  xnrc02aa1n12x5               g172(.a(\b[24] ), .b(\a[25] ), .out0(new_n268));
  aoib12aa1n06x5               g173(.a(new_n268), .b(new_n262), .c(new_n267), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n268), .o1(new_n270));
  aoi112aa1n02x5               g175(.a(new_n270), .b(new_n267), .c(new_n188), .d(new_n261), .o1(new_n271));
  norp02aa1n02x5               g176(.a(new_n269), .b(new_n271), .o1(\s[25] ));
  nor042aa1n03x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  nano22aa1n03x5               g180(.a(new_n269), .b(new_n274), .c(new_n275), .out0(new_n276));
  oaoi13aa1n03x5               g181(.a(new_n267), .b(new_n261), .c(new_n201), .d(new_n197), .o1(new_n277));
  oaoi13aa1n02x7               g182(.a(new_n275), .b(new_n274), .c(new_n277), .d(new_n268), .o1(new_n278));
  norp02aa1n03x5               g183(.a(new_n278), .b(new_n276), .o1(\s[26] ));
  nor042aa1n04x5               g184(.a(new_n275), .b(new_n268), .o1(new_n280));
  nano32aa1n03x7               g185(.a(new_n224), .b(new_n280), .c(new_n242), .d(new_n260), .out0(new_n281));
  oai012aa1n06x5               g186(.a(new_n281), .b(new_n201), .c(new_n197), .o1(new_n282));
  oao003aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .c(new_n274), .carry(new_n283));
  aobi12aa1n06x5               g188(.a(new_n283), .b(new_n267), .c(new_n280), .out0(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n282), .c(new_n284), .out0(\s[27] ));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  inv040aa1n03x5               g192(.a(new_n287), .o1(new_n288));
  aobi12aa1n02x7               g193(.a(new_n285), .b(new_n282), .c(new_n284), .out0(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[27] ), .b(\a[28] ), .out0(new_n290));
  nano22aa1n03x5               g195(.a(new_n289), .b(new_n288), .c(new_n290), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n260), .b(new_n246), .c(new_n229), .d(new_n242), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n280), .o1(new_n293));
  aoai13aa1n04x5               g198(.a(new_n283), .b(new_n293), .c(new_n292), .d(new_n266), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n285), .b(new_n294), .c(new_n188), .d(new_n281), .o1(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n290), .b(new_n295), .c(new_n288), .o1(new_n296));
  norp02aa1n03x5               g201(.a(new_n296), .b(new_n291), .o1(\s[28] ));
  norb02aa1n02x5               g202(.a(new_n285), .b(new_n290), .out0(new_n298));
  aobi12aa1n02x7               g203(.a(new_n298), .b(new_n282), .c(new_n284), .out0(new_n299));
  oao003aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .c(new_n288), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[28] ), .b(\a[29] ), .out0(new_n301));
  nano22aa1n03x5               g206(.a(new_n299), .b(new_n300), .c(new_n301), .out0(new_n302));
  aoai13aa1n02x5               g207(.a(new_n298), .b(new_n294), .c(new_n188), .d(new_n281), .o1(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n301), .b(new_n303), .c(new_n300), .o1(new_n304));
  norp02aa1n03x5               g209(.a(new_n304), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g211(.a(new_n285), .b(new_n301), .c(new_n290), .out0(new_n307));
  aobi12aa1n02x7               g212(.a(new_n307), .b(new_n282), .c(new_n284), .out0(new_n308));
  oao003aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[29] ), .b(\a[30] ), .out0(new_n310));
  nano22aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n310), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n307), .b(new_n294), .c(new_n188), .d(new_n281), .o1(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n310), .b(new_n312), .c(new_n309), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n313), .b(new_n311), .o1(\s[30] ));
  norb02aa1n02x5               g219(.a(new_n307), .b(new_n310), .out0(new_n315));
  aobi12aa1n02x7               g220(.a(new_n315), .b(new_n282), .c(new_n284), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  nano22aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n318), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n315), .b(new_n294), .c(new_n188), .d(new_n281), .o1(new_n320));
  tech160nm_fiaoi012aa1n02p5x5 g225(.a(new_n318), .b(new_n320), .c(new_n317), .o1(new_n321));
  norp02aa1n03x5               g226(.a(new_n321), .b(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g227(.a(new_n144), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g228(.a(\a[3] ), .b(\b[2] ), .c(new_n144), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n145), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g231(.a(new_n120), .b(new_n121), .c(new_n145), .o1(new_n327));
  xnrb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g233(.a(\a[6] ), .b(\b[5] ), .c(new_n327), .o1(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g235(.a(new_n114), .b(new_n329), .c(new_n115), .o1(new_n331));
  xnrb03aa1n02x5               g236(.a(new_n331), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g237(.a(new_n126), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


