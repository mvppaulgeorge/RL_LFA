// Benchmark "adder" written by ABC on Wed Jul 17 23:02:58 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n322, new_n324,
    new_n327, new_n328, new_n329, new_n331, new_n333;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n24x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor002aa1n03x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[8] ), .o1(new_n101));
  xnrc02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .out0(new_n102));
  nanp02aa1n02x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  norb03aa1n03x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n106));
  nor002aa1n20x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nanb03aa1n06x5               g013(.a(new_n107), .b(new_n108), .c(new_n104), .out0(new_n109));
  inv000aa1d42x5               g014(.a(new_n107), .o1(new_n110));
  oao003aa1n02x5               g015(.a(\a[4] ), .b(\b[3] ), .c(new_n110), .carry(new_n111));
  oai013aa1n03x5               g016(.a(new_n111), .b(new_n106), .c(new_n109), .d(new_n102), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  inv000aa1d42x5               g022(.a(\b[5] ), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(\a[6] ), .b(new_n118), .out0(new_n119));
  nand42aa1n03x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  oai112aa1n02x5               g025(.a(new_n119), .b(new_n120), .c(\b[4] ), .d(\a[5] ), .o1(new_n121));
  aoi112aa1n03x5               g026(.a(new_n117), .b(new_n121), .c(\a[5] ), .d(\b[4] ), .o1(new_n122));
  nand02aa1n04x5               g027(.a(new_n112), .b(new_n122), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n113), .o1(new_n124));
  aoi112aa1n06x5               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  nano22aa1n02x4               g031(.a(new_n117), .b(new_n121), .c(new_n120), .out0(new_n127));
  nano22aa1n03x7               g032(.a(new_n127), .b(new_n124), .c(new_n126), .out0(new_n128));
  nanp02aa1n06x5               g033(.a(new_n123), .b(new_n128), .o1(new_n129));
  tech160nm_fioaoi03aa1n03p5x5 g034(.a(new_n100), .b(new_n101), .c(new_n129), .o1(new_n130));
  xnrc02aa1n02x5               g035(.a(new_n130), .b(new_n99), .out0(\s[10] ));
  inv040aa1n02x5               g036(.a(new_n98), .o1(new_n132));
  nanp02aa1n03x5               g037(.a(new_n130), .b(new_n99), .o1(new_n133));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanp02aa1n03x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n133), .c(new_n132), .out0(\s[11] ));
  nona22aa1n03x5               g042(.a(new_n133), .b(new_n136), .c(new_n98), .out0(new_n138));
  nor042aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  nona22aa1n02x5               g047(.a(new_n138), .b(new_n142), .c(new_n134), .out0(new_n143));
  inv000aa1d42x5               g048(.a(new_n134), .o1(new_n144));
  tech160nm_fiaoi012aa1n03p5x5 g049(.a(new_n141), .b(new_n138), .c(new_n144), .o1(new_n145));
  norb02aa1n03x4               g050(.a(new_n143), .b(new_n145), .out0(\s[12] ));
  xorc02aa1n02x5               g051(.a(\a[9] ), .b(\b[8] ), .out0(new_n147));
  nona23aa1n09x5               g052(.a(new_n140), .b(new_n135), .c(new_n134), .d(new_n139), .out0(new_n148));
  norb02aa1n02x5               g053(.a(new_n99), .b(new_n148), .out0(new_n149));
  nand23aa1n03x5               g054(.a(new_n129), .b(new_n147), .c(new_n149), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n132), .b(new_n97), .c(new_n100), .d(new_n101), .o1(new_n151));
  oaoi03aa1n02x5               g056(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n152));
  oabi12aa1n09x5               g057(.a(new_n152), .b(new_n151), .c(new_n148), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  xnrc02aa1n12x5               g059(.a(\b[12] ), .b(\a[13] ), .out0(new_n155));
  xobna2aa1n03x5               g060(.a(new_n155), .b(new_n150), .c(new_n154), .out0(\s[13] ));
  tech160nm_fiao0012aa1n02p5x5 g061(.a(new_n155), .b(new_n150), .c(new_n154), .o(new_n157));
  inv000aa1d42x5               g062(.a(\a[14] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(\b[13] ), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(new_n159), .b(new_n158), .o1(new_n160));
  nor002aa1n02x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  oaoi03aa1n12x5               g066(.a(new_n158), .b(new_n159), .c(new_n161), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nano22aa1d15x5               g068(.a(new_n155), .b(new_n160), .c(new_n163), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n162), .b(new_n165), .c(new_n150), .d(new_n154), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n161), .b(new_n160), .c(new_n163), .o1(new_n167));
  aoi022aa1n02x5               g072(.a(new_n157), .b(new_n167), .c(new_n166), .d(new_n160), .o1(\s[14] ));
  xorb03aa1n02x5               g073(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  xnrc02aa1n12x5               g074(.a(\b[14] ), .b(\a[15] ), .out0(new_n170));
  nanb02aa1n02x5               g075(.a(new_n170), .b(new_n166), .out0(new_n171));
  inv000aa1d42x5               g076(.a(\a[16] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(\b[15] ), .o1(new_n173));
  nand42aa1n03x5               g078(.a(new_n173), .b(new_n172), .o1(new_n174));
  norp02aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n175), .b(new_n174), .c(new_n176), .o1(new_n177));
  nano23aa1n02x4               g082(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n178));
  nanp03aa1n02x5               g083(.a(new_n178), .b(new_n120), .c(new_n121), .o1(new_n179));
  nona22aa1n02x4               g084(.a(new_n179), .b(new_n125), .c(new_n113), .out0(new_n180));
  nano22aa1n09x5               g085(.a(new_n170), .b(new_n174), .c(new_n176), .out0(new_n181));
  nano23aa1n06x5               g086(.a(new_n134), .b(new_n139), .c(new_n140), .d(new_n135), .out0(new_n182));
  nand23aa1n03x5               g087(.a(new_n182), .b(new_n99), .c(new_n147), .o1(new_n183));
  nano22aa1n03x7               g088(.a(new_n183), .b(new_n164), .c(new_n181), .out0(new_n184));
  aoai13aa1n03x5               g089(.a(new_n184), .b(new_n180), .c(new_n112), .d(new_n122), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n162), .o1(new_n186));
  aoai13aa1n04x5               g091(.a(new_n181), .b(new_n186), .c(new_n153), .d(new_n164), .o1(new_n187));
  oaoi03aa1n02x5               g092(.a(new_n172), .b(new_n173), .c(new_n175), .o1(new_n188));
  nand03aa1n04x5               g093(.a(new_n185), .b(new_n187), .c(new_n188), .o1(new_n189));
  aoi022aa1n02x5               g094(.a(new_n171), .b(new_n177), .c(new_n174), .d(new_n189), .o1(\s[16] ));
  inv040aa1d30x5               g095(.a(\a[17] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n181), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(new_n101), .b(new_n100), .o1(new_n193));
  oaoi03aa1n02x5               g098(.a(\a[10] ), .b(\b[9] ), .c(new_n193), .o1(new_n194));
  aoai13aa1n09x5               g099(.a(new_n164), .b(new_n152), .c(new_n182), .d(new_n194), .o1(new_n195));
  aoai13aa1n12x5               g100(.a(new_n188), .b(new_n192), .c(new_n195), .d(new_n162), .o1(new_n196));
  tech160nm_fiaoi012aa1n05x5   g101(.a(new_n196), .b(new_n129), .c(new_n184), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[16] ), .c(new_n191), .out0(\s[17] ));
  nor002aa1n16x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nanb03aa1n02x5               g104(.a(new_n183), .b(new_n164), .c(new_n181), .out0(new_n200));
  aoi012aa1n06x5               g105(.a(new_n200), .b(new_n123), .c(new_n128), .o1(new_n201));
  inv040aa1d32x5               g106(.a(\a[18] ), .o1(new_n202));
  xroi22aa1d06x4               g107(.a(new_n191), .b(\b[16] ), .c(new_n202), .d(\b[17] ), .out0(new_n203));
  inv000aa1d42x5               g108(.a(\b[16] ), .o1(new_n204));
  nand42aa1n08x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  aoai13aa1n12x5               g110(.a(new_n205), .b(new_n199), .c(new_n191), .d(new_n204), .o1(new_n206));
  inv020aa1n02x5               g111(.a(new_n206), .o1(new_n207));
  oaoi13aa1n06x5               g112(.a(new_n207), .b(new_n203), .c(new_n201), .d(new_n196), .o1(new_n208));
  xorc02aa1n02x5               g113(.a(\a[17] ), .b(\b[16] ), .out0(new_n209));
  obai22aa1n02x7               g114(.a(new_n205), .b(new_n199), .c(\a[17] ), .d(\b[16] ), .out0(new_n210));
  oaoi13aa1n02x5               g115(.a(new_n210), .b(new_n209), .c(new_n201), .d(new_n196), .o1(new_n211));
  oab012aa1n02x4               g116(.a(new_n211), .b(new_n208), .c(new_n199), .out0(\s[18] ));
  nor002aa1d24x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nand42aa1n04x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n208), .b(new_n215), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g122(.a(new_n203), .o1(new_n218));
  nanb02aa1n06x5               g123(.a(new_n213), .b(new_n215), .out0(new_n219));
  oaoi13aa1n02x5               g124(.a(new_n219), .b(new_n206), .c(new_n197), .d(new_n218), .o1(new_n220));
  nor042aa1n04x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1d08x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanb02aa1n12x5               g127(.a(new_n221), .b(new_n222), .out0(new_n223));
  nano22aa1n02x4               g128(.a(new_n220), .b(new_n214), .c(new_n223), .out0(new_n224));
  oaoi13aa1n03x5               g129(.a(new_n223), .b(new_n214), .c(new_n208), .d(new_n219), .o1(new_n225));
  norp02aa1n02x5               g130(.a(new_n225), .b(new_n224), .o1(\s[20] ));
  nano23aa1d15x5               g131(.a(new_n213), .b(new_n221), .c(new_n222), .d(new_n215), .out0(new_n227));
  nand22aa1n12x5               g132(.a(new_n203), .b(new_n227), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoi012aa1d18x5               g134(.a(new_n221), .b(new_n213), .c(new_n222), .o1(new_n230));
  oai013aa1d12x5               g135(.a(new_n230), .b(new_n206), .c(new_n219), .d(new_n223), .o1(new_n231));
  oaoi13aa1n06x5               g136(.a(new_n231), .b(new_n229), .c(new_n201), .d(new_n196), .o1(new_n232));
  xnrb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  inv040aa1n03x5               g139(.a(new_n234), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n231), .o1(new_n236));
  xnrc02aa1n02x5               g141(.a(\b[20] ), .b(\a[21] ), .out0(new_n237));
  oaoi13aa1n02x7               g142(.a(new_n237), .b(new_n236), .c(new_n197), .d(new_n228), .o1(new_n238));
  tech160nm_fixnrc02aa1n02p5x5 g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  nano22aa1n03x7               g144(.a(new_n238), .b(new_n235), .c(new_n239), .out0(new_n240));
  oaoi13aa1n02x5               g145(.a(new_n239), .b(new_n235), .c(new_n232), .d(new_n237), .o1(new_n241));
  norp02aa1n02x5               g146(.a(new_n241), .b(new_n240), .o1(\s[22] ));
  nor002aa1n04x5               g147(.a(new_n239), .b(new_n237), .o1(new_n243));
  nano22aa1n02x4               g148(.a(new_n218), .b(new_n243), .c(new_n227), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n196), .c(new_n129), .d(new_n184), .o1(new_n245));
  oao003aa1n12x5               g150(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .carry(new_n246));
  inv040aa1d30x5               g151(.a(new_n246), .o1(new_n247));
  aoi012aa1n02x5               g152(.a(new_n247), .b(new_n231), .c(new_n243), .o1(new_n248));
  xnrc02aa1n12x5               g153(.a(\b[22] ), .b(\a[23] ), .out0(new_n249));
  xobna2aa1n03x5               g154(.a(new_n249), .b(new_n245), .c(new_n248), .out0(\s[23] ));
  nor042aa1n03x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  tech160nm_fiaoi012aa1n02p5x5 g157(.a(new_n249), .b(new_n245), .c(new_n248), .o1(new_n253));
  xnrc02aa1n06x5               g158(.a(\b[23] ), .b(\a[24] ), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n253), .b(new_n252), .c(new_n254), .out0(new_n255));
  inv000aa1n03x5               g160(.a(new_n248), .o1(new_n256));
  oaoi13aa1n02x5               g161(.a(new_n256), .b(new_n244), .c(new_n201), .d(new_n196), .o1(new_n257));
  oaoi13aa1n02x5               g162(.a(new_n254), .b(new_n252), .c(new_n257), .d(new_n249), .o1(new_n258));
  norp02aa1n02x5               g163(.a(new_n258), .b(new_n255), .o1(\s[24] ));
  nor002aa1n02x5               g164(.a(new_n254), .b(new_n249), .o1(new_n260));
  nano22aa1n03x7               g165(.a(new_n228), .b(new_n243), .c(new_n260), .out0(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n196), .c(new_n129), .d(new_n184), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n230), .o1(new_n263));
  aoai13aa1n06x5               g168(.a(new_n243), .b(new_n263), .c(new_n227), .d(new_n207), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n260), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n252), .carry(new_n266));
  aoai13aa1n12x5               g171(.a(new_n266), .b(new_n265), .c(new_n264), .d(new_n246), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  tech160nm_fixnrc02aa1n05x5   g173(.a(\b[24] ), .b(\a[25] ), .out0(new_n269));
  xobna2aa1n03x5               g174(.a(new_n269), .b(new_n262), .c(new_n268), .out0(\s[25] ));
  nor042aa1n03x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  tech160nm_fiaoi012aa1n05x5   g177(.a(new_n269), .b(new_n262), .c(new_n268), .o1(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[25] ), .b(\a[26] ), .out0(new_n274));
  nano22aa1n03x7               g179(.a(new_n273), .b(new_n272), .c(new_n274), .out0(new_n275));
  oaoi13aa1n02x5               g180(.a(new_n267), .b(new_n261), .c(new_n201), .d(new_n196), .o1(new_n276));
  oaoi13aa1n02x5               g181(.a(new_n274), .b(new_n272), .c(new_n276), .d(new_n269), .o1(new_n277));
  norp02aa1n02x5               g182(.a(new_n277), .b(new_n275), .o1(\s[26] ));
  nor042aa1n03x5               g183(.a(new_n274), .b(new_n269), .o1(new_n279));
  nano32aa1d12x5               g184(.a(new_n228), .b(new_n279), .c(new_n243), .d(new_n260), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n196), .c(new_n129), .d(new_n184), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[26] ), .b(\b[25] ), .c(new_n272), .carry(new_n282));
  aobi12aa1n12x5               g187(.a(new_n282), .b(new_n267), .c(new_n279), .out0(new_n283));
  xorc02aa1n02x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  xnbna2aa1n03x5               g189(.a(new_n284), .b(new_n281), .c(new_n283), .out0(\s[27] ));
  norp02aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  inv040aa1n03x5               g191(.a(new_n286), .o1(new_n287));
  aobi12aa1n02x7               g192(.a(new_n284), .b(new_n281), .c(new_n283), .out0(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[27] ), .b(\a[28] ), .out0(new_n289));
  nano22aa1n03x5               g194(.a(new_n288), .b(new_n287), .c(new_n289), .out0(new_n290));
  aoai13aa1n03x5               g195(.a(new_n260), .b(new_n247), .c(new_n231), .d(new_n243), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n279), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n282), .b(new_n292), .c(new_n291), .d(new_n266), .o1(new_n293));
  aoai13aa1n02x5               g198(.a(new_n284), .b(new_n293), .c(new_n189), .d(new_n280), .o1(new_n294));
  tech160nm_fiaoi012aa1n02p5x5 g199(.a(new_n289), .b(new_n294), .c(new_n287), .o1(new_n295));
  norp02aa1n03x5               g200(.a(new_n295), .b(new_n290), .o1(\s[28] ));
  xnrc02aa1n02x5               g201(.a(\b[28] ), .b(\a[29] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n284), .b(new_n289), .out0(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n293), .c(new_n189), .d(new_n280), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n297), .b(new_n299), .c(new_n300), .o1(new_n301));
  aobi12aa1n03x5               g206(.a(new_n298), .b(new_n281), .c(new_n283), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n297), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g210(.a(new_n284), .b(new_n297), .c(new_n289), .out0(new_n306));
  aoai13aa1n02x5               g211(.a(new_n306), .b(new_n293), .c(new_n189), .d(new_n280), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[29] ), .b(\a[30] ), .out0(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  aobi12aa1n02x7               g215(.a(new_n306), .b(new_n281), .c(new_n283), .out0(new_n311));
  nano22aa1n03x5               g216(.a(new_n311), .b(new_n308), .c(new_n309), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n310), .b(new_n312), .o1(\s[30] ));
  xnrc02aa1n02x5               g218(.a(\b[30] ), .b(\a[31] ), .out0(new_n314));
  norb02aa1n02x5               g219(.a(new_n306), .b(new_n309), .out0(new_n315));
  aobi12aa1n06x5               g220(.a(new_n315), .b(new_n281), .c(new_n283), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n317));
  nano22aa1n03x5               g222(.a(new_n316), .b(new_n314), .c(new_n317), .out0(new_n318));
  aoai13aa1n02x5               g223(.a(new_n315), .b(new_n293), .c(new_n189), .d(new_n280), .o1(new_n319));
  aoi012aa1n03x5               g224(.a(new_n314), .b(new_n319), .c(new_n317), .o1(new_n320));
  norp02aa1n02x5               g225(.a(new_n320), .b(new_n318), .o1(\s[31] ));
  aboi22aa1n03x5               g226(.a(new_n106), .b(new_n104), .c(new_n108), .d(new_n110), .out0(new_n322));
  oab012aa1n02x4               g227(.a(new_n322), .b(new_n106), .c(new_n109), .out0(\s[3] ));
  oai012aa1n02x5               g228(.a(new_n110), .b(new_n106), .c(new_n109), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g231(.a(\a[5] ), .o1(new_n327));
  inv000aa1d42x5               g232(.a(\b[4] ), .o1(new_n328));
  oaoi03aa1n02x5               g233(.a(new_n327), .b(new_n328), .c(new_n112), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n329), .b(new_n119), .c(new_n120), .out0(\s[6] ));
  oaoi03aa1n02x5               g235(.a(\a[6] ), .b(\b[5] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g237(.a(new_n115), .b(new_n331), .c(new_n116), .o1(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n124), .c(new_n114), .out0(\s[8] ));
  xnbna2aa1n03x5               g239(.a(new_n147), .b(new_n123), .c(new_n128), .out0(\s[9] ));
endmodule


