// Benchmark "adder" written by ABC on Thu Jul 11 12:55:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n307, new_n309, new_n311, new_n313,
    new_n315;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nanp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  and002aa1n02x5               g003(.a(\b[3] ), .b(\a[4] ), .o(new_n99));
  160nm_ficinv00aa1n08x5       g004(.clk(\a[3] ), .clkout(new_n100));
  160nm_ficinv00aa1n08x5       g005(.clk(\b[2] ), .clkout(new_n101));
  nanp02aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(new_n102), .b(new_n103), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  norp02aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  oai012aa1n02x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .o1(new_n108));
  oa0022aa1n02x5               g013(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n109));
  oai012aa1n02x5               g014(.a(new_n109), .b(new_n108), .c(new_n104), .o1(new_n110));
  norp02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  norp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n02x4               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  norp02aa1n02x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  nona23aa1n02x4               g023(.a(new_n110), .b(new_n118), .c(new_n115), .d(new_n99), .out0(new_n119));
  nano23aa1n02x4               g024(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n120));
  orn002aa1n02x5               g025(.a(\a[5] ), .b(\b[4] ), .o(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  oai012aa1n02x5               g027(.a(new_n112), .b(new_n113), .c(new_n111), .o1(new_n123));
  aobi12aa1n02x5               g028(.a(new_n123), .b(new_n120), .c(new_n122), .out0(new_n124));
  oai112aa1n02x5               g029(.a(new_n119), .b(new_n124), .c(\b[8] ), .d(\a[9] ), .o1(new_n125));
  xobna2aa1n03x5               g030(.a(new_n97), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  orn002aa1n02x5               g031(.a(\a[10] ), .b(\b[9] ), .o(new_n127));
  and002aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  nanp02aa1n02x5               g033(.a(new_n125), .b(new_n98), .o1(new_n129));
  norp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  160nm_ficinv00aa1n08x5       g037(.clk(new_n132), .clkout(new_n133));
  aoi112aa1n02x5               g038(.a(new_n133), .b(new_n128), .c(new_n129), .d(new_n127), .o1(new_n134));
  aoai13aa1n02x5               g039(.a(new_n133), .b(new_n128), .c(new_n129), .d(new_n127), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(\s[11] ));
  norp02aa1n02x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanp02aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(new_n139));
  oai012aa1n02x5               g044(.a(new_n139), .b(new_n134), .c(new_n130), .o1(new_n140));
  norp03aa1n02x5               g045(.a(new_n134), .b(new_n139), .c(new_n130), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(\s[12] ));
  nano23aa1n02x4               g047(.a(new_n130), .b(new_n137), .c(new_n138), .d(new_n131), .out0(new_n143));
  oaoi13aa1n02x5               g048(.a(new_n128), .b(new_n127), .c(\a[9] ), .d(\b[8] ), .o1(new_n144));
  oa0012aa1n02x5               g049(.a(new_n138), .b(new_n137), .c(new_n130), .o(new_n145));
  aoi012aa1n02x5               g050(.a(new_n145), .b(new_n143), .c(new_n144), .o1(new_n146));
  xorc02aa1n02x5               g051(.a(\a[9] ), .b(\b[8] ), .out0(new_n147));
  nanp03aa1n02x5               g052(.a(new_n143), .b(new_n97), .c(new_n147), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n146), .b(new_n148), .c(new_n119), .d(new_n124), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  160nm_ficinv00aa1n08x5       g055(.clk(\a[14] ), .clkout(new_n151));
  norp02aa1n02x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  xnrc02aa1n02x5               g057(.a(\b[12] ), .b(\a[13] ), .out0(new_n153));
  aoib12aa1n02x5               g058(.a(new_n152), .b(new_n149), .c(new_n153), .out0(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(new_n151), .out0(\s[14] ));
  xnrc02aa1n02x5               g060(.a(\b[13] ), .b(\a[14] ), .out0(new_n156));
  norp02aa1n02x5               g061(.a(new_n156), .b(new_n153), .o1(new_n157));
  160nm_ficinv00aa1n08x5       g062(.clk(\b[13] ), .clkout(new_n158));
  oao003aa1n02x5               g063(.a(new_n151), .b(new_n158), .c(new_n152), .carry(new_n159));
  160nm_fiao0012aa1n02p5x5     g064(.a(new_n159), .b(new_n149), .c(new_n157), .o(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  xnrc02aa1n02x5               g067(.a(\b[14] ), .b(\a[15] ), .out0(new_n163));
  160nm_ficinv00aa1n08x5       g068(.clk(new_n163), .clkout(new_n164));
  norp02aa1n02x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n162), .c(new_n160), .d(new_n164), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n164), .b(new_n159), .c(new_n149), .d(new_n157), .o1(new_n169));
  nona22aa1n02x4               g074(.a(new_n169), .b(new_n167), .c(new_n162), .out0(new_n170));
  nanp02aa1n02x5               g075(.a(new_n168), .b(new_n170), .o1(\s[16] ));
  nanp02aa1n02x5               g076(.a(new_n119), .b(new_n124), .o1(new_n172));
  norp02aa1n02x5               g077(.a(new_n163), .b(new_n167), .o1(new_n173));
  nano22aa1n02x4               g078(.a(new_n148), .b(new_n157), .c(new_n173), .out0(new_n174));
  nanp02aa1n02x5               g079(.a(new_n172), .b(new_n174), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n157), .b(new_n173), .o1(new_n176));
  oai022aa1n02x5               g081(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n177));
  aoi022aa1n02x5               g082(.a(new_n173), .b(new_n159), .c(new_n166), .d(new_n177), .o1(new_n178));
  oai012aa1n02x5               g083(.a(new_n178), .b(new_n146), .c(new_n176), .o1(new_n179));
  160nm_ficinv00aa1n08x5       g084(.clk(new_n179), .clkout(new_n180));
  xorc02aa1n02x5               g085(.a(\a[17] ), .b(\b[16] ), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n175), .c(new_n180), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g087(.clk(\a[17] ), .clkout(new_n183));
  nanb02aa1n02x5               g088(.a(\b[16] ), .b(new_n183), .out0(new_n184));
  aoai13aa1n02x5               g089(.a(new_n181), .b(new_n179), .c(new_n172), .d(new_n174), .o1(new_n185));
  xnrc02aa1n02x5               g090(.a(\b[17] ), .b(\a[18] ), .out0(new_n186));
  xobna2aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n184), .out0(\s[18] ));
  160nm_ficinv00aa1n08x5       g092(.clk(\a[18] ), .clkout(new_n188));
  xroi22aa1d04x5               g093(.a(new_n183), .b(\b[16] ), .c(new_n188), .d(\b[17] ), .out0(new_n189));
  aoai13aa1n02x5               g094(.a(new_n189), .b(new_n179), .c(new_n172), .d(new_n174), .o1(new_n190));
  oai022aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n191));
  oaib12aa1n02x5               g096(.a(new_n191), .b(new_n188), .c(\b[17] ), .out0(new_n192));
  norp02aa1n02x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  160nm_ficinv00aa1n08x5       g100(.clk(new_n195), .clkout(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n190), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g103(.a(new_n190), .b(new_n192), .o1(new_n199));
  norp02aa1n02x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(new_n200), .b(new_n201), .out0(new_n202));
  aoai13aa1n02x5               g107(.a(new_n202), .b(new_n193), .c(new_n199), .d(new_n196), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n199), .b(new_n196), .o1(new_n204));
  nona22aa1n02x4               g109(.a(new_n204), .b(new_n202), .c(new_n193), .out0(new_n205));
  nanp02aa1n02x5               g110(.a(new_n205), .b(new_n203), .o1(\s[20] ));
  nona23aa1n02x4               g111(.a(new_n201), .b(new_n194), .c(new_n193), .d(new_n200), .out0(new_n207));
  oai012aa1n02x5               g112(.a(new_n201), .b(new_n200), .c(new_n193), .o1(new_n208));
  oai012aa1n02x5               g113(.a(new_n208), .b(new_n207), .c(new_n192), .o1(new_n209));
  160nm_ficinv00aa1n08x5       g114(.clk(new_n209), .clkout(new_n210));
  nano23aa1n02x4               g115(.a(new_n193), .b(new_n200), .c(new_n201), .d(new_n194), .out0(new_n211));
  nanb03aa1n02x5               g116(.a(new_n186), .b(new_n211), .c(new_n181), .out0(new_n212));
  aoai13aa1n02x5               g117(.a(new_n210), .b(new_n212), .c(new_n175), .d(new_n180), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  xorc02aa1n02x5               g121(.a(\a[22] ), .b(\b[21] ), .out0(new_n217));
  160nm_ficinv00aa1n08x5       g122(.clk(new_n217), .clkout(new_n218));
  aoai13aa1n02x5               g123(.a(new_n218), .b(new_n215), .c(new_n213), .d(new_n216), .o1(new_n219));
  nanp02aa1n02x5               g124(.a(new_n213), .b(new_n216), .o1(new_n220));
  nona22aa1n02x4               g125(.a(new_n220), .b(new_n218), .c(new_n215), .out0(new_n221));
  nanp02aa1n02x5               g126(.a(new_n221), .b(new_n219), .o1(\s[22] ));
  160nm_ficinv00aa1n08x5       g127(.clk(\a[21] ), .clkout(new_n223));
  160nm_ficinv00aa1n08x5       g128(.clk(\a[22] ), .clkout(new_n224));
  xroi22aa1d04x5               g129(.a(new_n223), .b(\b[20] ), .c(new_n224), .d(\b[21] ), .out0(new_n225));
  160nm_ficinv00aa1n08x5       g130(.clk(\b[21] ), .clkout(new_n226));
  oao003aa1n02x5               g131(.a(new_n224), .b(new_n226), .c(new_n215), .carry(new_n227));
  aoi012aa1n02x5               g132(.a(new_n227), .b(new_n209), .c(new_n225), .o1(new_n228));
  nanp03aa1n02x5               g133(.a(new_n225), .b(new_n189), .c(new_n211), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n228), .b(new_n229), .c(new_n175), .d(new_n180), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  xnrc02aa1n02x5               g138(.a(\b[23] ), .b(\a[24] ), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n235));
  nanp02aa1n02x5               g140(.a(new_n230), .b(new_n233), .o1(new_n236));
  nona22aa1n02x4               g141(.a(new_n236), .b(new_n234), .c(new_n232), .out0(new_n237));
  nanp02aa1n02x5               g142(.a(new_n237), .b(new_n235), .o1(\s[24] ));
  norb02aa1n02x5               g143(.a(new_n233), .b(new_n234), .out0(new_n239));
  nano22aa1n02x4               g144(.a(new_n212), .b(new_n239), .c(new_n225), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n179), .c(new_n172), .d(new_n174), .o1(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[18] ), .b(\b[17] ), .c(new_n184), .o1(new_n242));
  160nm_ficinv00aa1n08x5       g147(.clk(new_n208), .clkout(new_n243));
  aoai13aa1n02x5               g148(.a(new_n225), .b(new_n243), .c(new_n211), .d(new_n242), .o1(new_n244));
  160nm_ficinv00aa1n08x5       g149(.clk(new_n227), .clkout(new_n245));
  160nm_ficinv00aa1n08x5       g150(.clk(new_n239), .clkout(new_n246));
  oai022aa1n02x5               g151(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n247));
  aob012aa1n02x5               g152(.a(new_n247), .b(\b[23] ), .c(\a[24] ), .out0(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n246), .c(new_n244), .d(new_n245), .o1(new_n249));
  nanb02aa1n02x5               g154(.a(new_n249), .b(new_n241), .out0(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[25] ), .b(\b[24] ), .out0(new_n253));
  norp02aa1n02x5               g158(.a(\b[25] ), .b(\a[26] ), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(\b[25] ), .b(\a[26] ), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n255), .b(new_n254), .out0(new_n256));
  160nm_ficinv00aa1n08x5       g161(.clk(new_n256), .clkout(new_n257));
  aoai13aa1n02x5               g162(.a(new_n257), .b(new_n252), .c(new_n250), .d(new_n253), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(new_n175), .b(new_n180), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n253), .b(new_n249), .c(new_n259), .d(new_n240), .o1(new_n260));
  nona22aa1n02x4               g165(.a(new_n260), .b(new_n257), .c(new_n252), .out0(new_n261));
  nanp02aa1n02x5               g166(.a(new_n258), .b(new_n261), .o1(\s[26] ));
  norb02aa1n02x5               g167(.a(new_n253), .b(new_n257), .out0(new_n263));
  nano22aa1n02x4               g168(.a(new_n229), .b(new_n239), .c(new_n263), .out0(new_n264));
  aoai13aa1n02x5               g169(.a(new_n264), .b(new_n179), .c(new_n172), .d(new_n174), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(new_n249), .b(new_n263), .o1(new_n266));
  oai012aa1n02x5               g171(.a(new_n255), .b(new_n254), .c(new_n252), .o1(new_n267));
  nanp03aa1n02x5               g172(.a(new_n265), .b(new_n266), .c(new_n267), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[27] ), .b(\b[26] ), .out0(new_n271));
  xnrc02aa1n02x5               g176(.a(\b[27] ), .b(\a[28] ), .out0(new_n272));
  aoai13aa1n02x5               g177(.a(new_n272), .b(new_n270), .c(new_n268), .d(new_n271), .o1(new_n273));
  aoai13aa1n02x5               g178(.a(new_n239), .b(new_n227), .c(new_n209), .d(new_n225), .o1(new_n274));
  160nm_ficinv00aa1n08x5       g179(.clk(new_n263), .clkout(new_n275));
  aoai13aa1n02x5               g180(.a(new_n267), .b(new_n275), .c(new_n274), .d(new_n248), .o1(new_n276));
  aoai13aa1n02x5               g181(.a(new_n271), .b(new_n276), .c(new_n259), .d(new_n264), .o1(new_n277));
  nona22aa1n02x4               g182(.a(new_n277), .b(new_n272), .c(new_n270), .out0(new_n278));
  nanp02aa1n02x5               g183(.a(new_n273), .b(new_n278), .o1(\s[28] ));
  norb02aa1n02x5               g184(.a(new_n271), .b(new_n272), .out0(new_n280));
  aoai13aa1n02x5               g185(.a(new_n280), .b(new_n276), .c(new_n259), .d(new_n264), .o1(new_n281));
  160nm_ficinv00aa1n08x5       g186(.clk(new_n270), .clkout(new_n282));
  oaoi03aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .o1(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[28] ), .b(\a[29] ), .out0(new_n284));
  nona22aa1n02x4               g189(.a(new_n281), .b(new_n283), .c(new_n284), .out0(new_n285));
  aoai13aa1n02x5               g190(.a(new_n284), .b(new_n283), .c(new_n268), .d(new_n280), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(new_n286), .b(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g193(.a(new_n271), .b(new_n284), .c(new_n272), .out0(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .carry(new_n290));
  oaoi03aa1n02x5               g195(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[30] ), .b(\b[29] ), .out0(new_n292));
  160nm_ficinv00aa1n08x5       g197(.clk(new_n292), .clkout(new_n293));
  aoai13aa1n02x5               g198(.a(new_n293), .b(new_n291), .c(new_n268), .d(new_n289), .o1(new_n294));
  aoai13aa1n02x5               g199(.a(new_n289), .b(new_n276), .c(new_n259), .d(new_n264), .o1(new_n295));
  nona22aa1n02x4               g200(.a(new_n295), .b(new_n291), .c(new_n293), .out0(new_n296));
  nanp02aa1n02x5               g201(.a(new_n294), .b(new_n296), .o1(\s[30] ));
  nano23aa1n02x4               g202(.a(new_n284), .b(new_n272), .c(new_n292), .d(new_n271), .out0(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n276), .c(new_n259), .d(new_n264), .o1(new_n299));
  nanp02aa1n02x5               g204(.a(new_n291), .b(new_n292), .o1(new_n300));
  oai012aa1n02x5               g205(.a(new_n300), .b(\b[29] ), .c(\a[30] ), .o1(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[30] ), .b(\a[31] ), .out0(new_n302));
  nona22aa1n02x4               g207(.a(new_n299), .b(new_n301), .c(new_n302), .out0(new_n303));
  aoai13aa1n02x5               g208(.a(new_n302), .b(new_n301), .c(new_n268), .d(new_n298), .o1(new_n304));
  nanp02aa1n02x5               g209(.a(new_n304), .b(new_n303), .o1(\s[31] ));
  xnbna2aa1n03x5               g210(.a(new_n108), .b(new_n102), .c(new_n103), .out0(\s[3] ));
  oaoi03aa1n02x5               g211(.a(\a[3] ), .b(\b[2] ), .c(new_n108), .o1(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  oaoi13aa1n02x5               g213(.a(new_n99), .b(new_n109), .c(new_n108), .d(new_n104), .o1(new_n309));
  xorb03aa1n02x5               g214(.a(new_n309), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nona22aa1n02x4               g215(.a(new_n110), .b(new_n117), .c(new_n99), .out0(new_n311));
  xobna2aa1n03x5               g216(.a(new_n116), .b(new_n311), .c(new_n121), .out0(\s[6] ));
  aoi012aa1n02x5               g217(.a(new_n122), .b(new_n309), .c(new_n118), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g219(.a(\a[7] ), .b(\b[6] ), .c(new_n313), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g221(.a(new_n147), .b(new_n119), .c(new_n124), .out0(\s[9] ));
endmodule


