// Benchmark "adder" written by ABC on Wed Jul 17 12:27:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n319,
    new_n320, new_n322, new_n323, new_n324, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  and002aa1n24x5               g001(.a(\b[8] ), .b(\a[9] ), .o(new_n97));
  inv040aa1d32x5               g002(.a(\a[9] ), .o1(new_n98));
  inv040aa1d28x5               g003(.a(\b[8] ), .o1(new_n99));
  nand02aa1n03x5               g004(.a(new_n99), .b(new_n98), .o1(new_n100));
  inv000aa1n03x5               g005(.a(new_n100), .o1(new_n101));
  and002aa1n12x5               g006(.a(\b[1] ), .b(\a[2] ), .o(new_n102));
  nand02aa1d16x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor002aa1n10x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oab012aa1d18x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .out0(new_n105));
  xorc02aa1n12x5               g010(.a(\a[4] ), .b(\b[3] ), .out0(new_n106));
  nor042aa1d18x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nanp03aa1d12x5               g014(.a(new_n105), .b(new_n106), .c(new_n109), .o1(new_n110));
  inv030aa1n02x5               g015(.a(new_n107), .o1(new_n111));
  oao003aa1n06x5               g016(.a(\a[4] ), .b(\b[3] ), .c(new_n111), .carry(new_n112));
  nor042aa1n03x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1d28x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor042aa1d18x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1d28x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n09x5               g021(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n117));
  tech160nm_fixorc02aa1n04x5   g022(.a(\a[6] ), .b(\b[5] ), .out0(new_n118));
  xorc02aa1n12x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nand23aa1n03x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  inv040aa1d28x5               g025(.a(\a[6] ), .o1(new_n121));
  inv040aa1d32x5               g026(.a(\b[5] ), .o1(new_n122));
  nor022aa1n16x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  oao003aa1n03x5               g028(.a(new_n121), .b(new_n122), .c(new_n123), .carry(new_n124));
  inv000aa1n02x5               g029(.a(new_n115), .o1(new_n125));
  oaoi03aa1n03x5               g030(.a(\a[8] ), .b(\b[7] ), .c(new_n125), .o1(new_n126));
  aoi012aa1n06x5               g031(.a(new_n126), .b(new_n117), .c(new_n124), .o1(new_n127));
  aoai13aa1n12x5               g032(.a(new_n127), .b(new_n120), .c(new_n110), .d(new_n112), .o1(new_n128));
  oab012aa1n02x4               g033(.a(new_n97), .b(new_n128), .c(new_n101), .out0(new_n129));
  xorb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1n08x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nor042aa1n06x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  norb02aa1n15x5               g037(.a(new_n131), .b(new_n132), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n97), .o1(new_n135));
  oaoi13aa1n03x5               g040(.a(new_n134), .b(new_n135), .c(new_n128), .d(new_n101), .o1(new_n136));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand42aa1d28x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  nano22aa1n03x5               g044(.a(new_n136), .b(new_n131), .c(new_n139), .out0(new_n140));
  oaoi13aa1n02x5               g045(.a(new_n139), .b(new_n131), .c(new_n129), .d(new_n134), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n141), .b(new_n140), .o1(\s[11] ));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n16x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  oai012aa1n02x5               g050(.a(new_n145), .b(new_n140), .c(new_n137), .o1(new_n146));
  orn003aa1n03x5               g051(.a(new_n140), .b(new_n137), .c(new_n145), .o(new_n147));
  nanp02aa1n03x5               g052(.a(new_n147), .b(new_n146), .o1(\s[12] ));
  nona23aa1n03x5               g053(.a(new_n144), .b(new_n138), .c(new_n137), .d(new_n143), .out0(new_n149));
  aoai13aa1n03x5               g054(.a(new_n131), .b(new_n132), .c(new_n98), .d(new_n99), .o1(new_n150));
  oa0012aa1n03x5               g055(.a(new_n144), .b(new_n143), .c(new_n137), .o(new_n151));
  oabi12aa1n06x5               g056(.a(new_n151), .b(new_n149), .c(new_n150), .out0(new_n152));
  nano23aa1d15x5               g057(.a(new_n137), .b(new_n143), .c(new_n144), .d(new_n138), .out0(new_n153));
  nona23aa1d16x5               g058(.a(new_n153), .b(new_n133), .c(new_n97), .d(new_n101), .out0(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  xnrc02aa1n12x5               g060(.a(\b[12] ), .b(\a[13] ), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n152), .c(new_n128), .d(new_n155), .o1(new_n158));
  aoi112aa1n02x5               g063(.a(new_n152), .b(new_n157), .c(new_n128), .d(new_n155), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(\s[13] ));
  nor042aa1n03x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  inv000aa1n03x5               g066(.a(new_n161), .o1(new_n162));
  tech160nm_fixnrc02aa1n04x5   g067(.a(\b[13] ), .b(\a[14] ), .out0(new_n163));
  xobna2aa1n03x5               g068(.a(new_n163), .b(new_n158), .c(new_n162), .out0(\s[14] ));
  nor042aa1n09x5               g069(.a(new_n163), .b(new_n156), .o1(new_n165));
  tech160nm_fioaoi03aa1n02p5x5 g070(.a(\a[14] ), .b(\b[13] ), .c(new_n162), .o1(new_n166));
  tech160nm_fiaoi012aa1n04x5   g071(.a(new_n166), .b(new_n152), .c(new_n165), .o1(new_n167));
  nona32aa1n09x5               g072(.a(new_n128), .b(new_n163), .c(new_n156), .d(new_n154), .out0(new_n168));
  xnrc02aa1n12x5               g073(.a(\b[14] ), .b(\a[15] ), .out0(new_n169));
  xobna2aa1n03x5               g074(.a(new_n169), .b(new_n168), .c(new_n167), .out0(\s[15] ));
  nor002aa1n03x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  ao0012aa1n03x5               g076(.a(new_n169), .b(new_n168), .c(new_n167), .o(new_n172));
  xnrc02aa1n12x5               g077(.a(\b[15] ), .b(\a[16] ), .out0(new_n173));
  oaib12aa1n03x5               g078(.a(new_n173), .b(new_n171), .c(new_n172), .out0(new_n174));
  nona22aa1n02x4               g079(.a(new_n172), .b(new_n173), .c(new_n171), .out0(new_n175));
  nanp02aa1n03x5               g080(.a(new_n174), .b(new_n175), .o1(\s[16] ));
  inv040aa1d32x5               g081(.a(\a[17] ), .o1(new_n177));
  nor042aa1n04x5               g082(.a(new_n173), .b(new_n169), .o1(new_n178));
  nano22aa1d15x5               g083(.a(new_n154), .b(new_n165), .c(new_n178), .out0(new_n179));
  inv000aa1d42x5               g084(.a(\a[16] ), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\b[15] ), .o1(new_n181));
  oao003aa1n12x5               g086(.a(new_n180), .b(new_n181), .c(new_n171), .carry(new_n182));
  oaoi03aa1n02x5               g087(.a(\a[10] ), .b(\b[9] ), .c(new_n100), .o1(new_n183));
  aoai13aa1n03x5               g088(.a(new_n165), .b(new_n151), .c(new_n153), .d(new_n183), .o1(new_n184));
  inv000aa1n02x5               g089(.a(new_n166), .o1(new_n185));
  inv000aa1n02x5               g090(.a(new_n178), .o1(new_n186));
  aoi012aa1n06x5               g091(.a(new_n186), .b(new_n184), .c(new_n185), .o1(new_n187));
  aoi112aa1n09x5               g092(.a(new_n187), .b(new_n182), .c(new_n128), .d(new_n179), .o1(new_n188));
  xorb03aa1n03x5               g093(.a(new_n188), .b(\b[16] ), .c(new_n177), .out0(\s[17] ));
  oaoi03aa1n03x5               g094(.a(\a[17] ), .b(\b[16] ), .c(new_n188), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g096(.a(\a[18] ), .o1(new_n192));
  xroi22aa1d06x4               g097(.a(new_n177), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n193));
  inv000aa1n02x5               g098(.a(new_n193), .o1(new_n194));
  oai022aa1n04x7               g099(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n195));
  oaib12aa1n09x5               g100(.a(new_n195), .b(new_n192), .c(\b[17] ), .out0(new_n196));
  tech160nm_fioai012aa1n05x5   g101(.a(new_n196), .b(new_n188), .c(new_n194), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g103(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand02aa1d16x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(new_n200), .b(new_n201), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  norp02aa1n24x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand22aa1n12x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  aoai13aa1n02x7               g111(.a(new_n206), .b(new_n200), .c(new_n197), .d(new_n203), .o1(new_n207));
  tech160nm_finand02aa1n05x5   g112(.a(new_n128), .b(new_n179), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n182), .o1(new_n209));
  oai112aa1n06x5               g114(.a(new_n208), .b(new_n209), .c(new_n167), .d(new_n186), .o1(new_n210));
  nanb02aa1n02x5               g115(.a(\b[16] ), .b(new_n177), .out0(new_n211));
  oaoi03aa1n12x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n211), .o1(new_n212));
  aoai13aa1n02x7               g117(.a(new_n203), .b(new_n212), .c(new_n210), .d(new_n193), .o1(new_n213));
  nona22aa1n03x5               g118(.a(new_n213), .b(new_n206), .c(new_n200), .out0(new_n214));
  nanp02aa1n03x5               g119(.a(new_n207), .b(new_n214), .o1(\s[20] ));
  nona23aa1n09x5               g120(.a(new_n205), .b(new_n201), .c(new_n200), .d(new_n204), .out0(new_n216));
  oa0012aa1n03x5               g121(.a(new_n205), .b(new_n204), .c(new_n200), .o(new_n217));
  inv040aa1n03x5               g122(.a(new_n217), .o1(new_n218));
  oai012aa1n18x5               g123(.a(new_n218), .b(new_n216), .c(new_n196), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  nano23aa1n06x5               g125(.a(new_n200), .b(new_n204), .c(new_n205), .d(new_n201), .out0(new_n221));
  nand02aa1d06x5               g126(.a(new_n193), .b(new_n221), .o1(new_n222));
  tech160nm_fioai012aa1n05x5   g127(.a(new_n220), .b(new_n188), .c(new_n222), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  aoai13aa1n02x7               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n222), .o1(new_n230));
  aoai13aa1n02x7               g135(.a(new_n227), .b(new_n219), .c(new_n210), .d(new_n230), .o1(new_n231));
  nona22aa1n03x5               g136(.a(new_n231), .b(new_n228), .c(new_n225), .out0(new_n232));
  nanp02aa1n03x5               g137(.a(new_n229), .b(new_n232), .o1(\s[22] ));
  nor042aa1n06x5               g138(.a(new_n228), .b(new_n226), .o1(new_n234));
  inv000aa1n09x5               g139(.a(\a[22] ), .o1(new_n235));
  inv040aa1d32x5               g140(.a(\b[21] ), .o1(new_n236));
  oao003aa1n06x5               g141(.a(new_n235), .b(new_n236), .c(new_n225), .carry(new_n237));
  aoi012aa1d18x5               g142(.a(new_n237), .b(new_n219), .c(new_n234), .o1(new_n238));
  nano22aa1n06x5               g143(.a(new_n194), .b(new_n234), .c(new_n221), .out0(new_n239));
  inv000aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  tech160nm_fioai012aa1n05x5   g145(.a(new_n238), .b(new_n188), .c(new_n240), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  tech160nm_fixnrc02aa1n05x5   g149(.a(\b[23] ), .b(\a[24] ), .out0(new_n245));
  aoai13aa1n02x7               g150(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n238), .o1(new_n247));
  aoai13aa1n02x7               g152(.a(new_n244), .b(new_n247), .c(new_n210), .d(new_n239), .o1(new_n248));
  nona22aa1n03x5               g153(.a(new_n248), .b(new_n245), .c(new_n243), .out0(new_n249));
  nanp02aa1n03x5               g154(.a(new_n246), .b(new_n249), .o1(\s[24] ));
  norb02aa1n02x7               g155(.a(new_n244), .b(new_n245), .out0(new_n251));
  inv030aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  nano32aa1n03x7               g157(.a(new_n252), .b(new_n193), .c(new_n234), .d(new_n221), .out0(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n234), .b(new_n217), .c(new_n221), .d(new_n212), .o1(new_n255));
  inv030aa1n02x5               g160(.a(new_n237), .o1(new_n256));
  oai022aa1n02x5               g161(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n257));
  aob012aa1n02x5               g162(.a(new_n257), .b(\b[23] ), .c(\a[24] ), .out0(new_n258));
  aoai13aa1n02x7               g163(.a(new_n258), .b(new_n252), .c(new_n255), .d(new_n256), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  tech160nm_fioai012aa1n05x5   g165(.a(new_n260), .b(new_n188), .c(new_n254), .o1(new_n261));
  xorb03aa1n02x5               g166(.a(new_n261), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  xorc02aa1n03x5               g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  xnrc02aa1n12x5               g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  aoai13aa1n02x7               g170(.a(new_n265), .b(new_n263), .c(new_n261), .d(new_n264), .o1(new_n266));
  aoai13aa1n02x7               g171(.a(new_n264), .b(new_n259), .c(new_n210), .d(new_n253), .o1(new_n267));
  nona22aa1n03x5               g172(.a(new_n267), .b(new_n265), .c(new_n263), .out0(new_n268));
  nanp02aa1n03x5               g173(.a(new_n266), .b(new_n268), .o1(\s[26] ));
  norb02aa1n09x5               g174(.a(new_n264), .b(new_n265), .out0(new_n270));
  nano23aa1n06x5               g175(.a(new_n222), .b(new_n252), .c(new_n270), .d(new_n234), .out0(new_n271));
  inv000aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .o1(new_n273));
  oai022aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n274));
  aoi022aa1n02x7               g179(.a(new_n259), .b(new_n270), .c(new_n273), .d(new_n274), .o1(new_n275));
  tech160nm_fioai012aa1n05x5   g180(.a(new_n275), .b(new_n188), .c(new_n272), .o1(new_n276));
  xorb03aa1n03x5               g181(.a(new_n276), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[27] ), .b(\a[28] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n278), .c(new_n276), .d(new_n279), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n251), .b(new_n237), .c(new_n219), .d(new_n234), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n270), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n274), .b(new_n273), .o1(new_n284));
  aoai13aa1n04x5               g189(.a(new_n284), .b(new_n283), .c(new_n282), .d(new_n258), .o1(new_n285));
  aoai13aa1n02x7               g190(.a(new_n279), .b(new_n285), .c(new_n210), .d(new_n271), .o1(new_n286));
  nona22aa1n02x4               g191(.a(new_n286), .b(new_n280), .c(new_n278), .out0(new_n287));
  nanp02aa1n03x5               g192(.a(new_n281), .b(new_n287), .o1(\s[28] ));
  norb02aa1n02x5               g193(.a(new_n279), .b(new_n280), .out0(new_n289));
  aoai13aa1n02x7               g194(.a(new_n289), .b(new_n285), .c(new_n210), .d(new_n271), .o1(new_n290));
  inv000aa1n03x5               g195(.a(new_n278), .o1(new_n291));
  oaoi03aa1n02x5               g196(.a(\a[28] ), .b(\b[27] ), .c(new_n291), .o1(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  nona22aa1n02x4               g198(.a(new_n290), .b(new_n292), .c(new_n293), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n293), .b(new_n292), .c(new_n276), .d(new_n289), .o1(new_n295));
  nanp02aa1n03x5               g200(.a(new_n295), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g202(.a(new_n279), .b(new_n293), .c(new_n280), .out0(new_n298));
  oao003aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .c(new_n291), .carry(new_n299));
  oaoi03aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n299), .o1(new_n300));
  tech160nm_fixorc02aa1n03p5x5 g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n300), .c(new_n276), .d(new_n298), .o1(new_n303));
  aoai13aa1n02x7               g208(.a(new_n298), .b(new_n285), .c(new_n210), .d(new_n271), .o1(new_n304));
  nona22aa1n02x4               g209(.a(new_n304), .b(new_n300), .c(new_n302), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n303), .b(new_n305), .o1(\s[30] ));
  nano23aa1n02x4               g211(.a(new_n293), .b(new_n280), .c(new_n301), .d(new_n279), .out0(new_n307));
  aoai13aa1n02x7               g212(.a(new_n307), .b(new_n285), .c(new_n210), .d(new_n271), .o1(new_n308));
  nanp02aa1n02x5               g213(.a(new_n300), .b(new_n301), .o1(new_n309));
  oai012aa1n02x5               g214(.a(new_n309), .b(\b[29] ), .c(\a[30] ), .o1(new_n310));
  xnrc02aa1n02x5               g215(.a(\b[30] ), .b(\a[31] ), .out0(new_n311));
  nona22aa1n02x4               g216(.a(new_n308), .b(new_n310), .c(new_n311), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n311), .b(new_n310), .c(new_n276), .d(new_n307), .o1(new_n313));
  nanp02aa1n03x5               g218(.a(new_n313), .b(new_n312), .o1(\s[31] ));
  xobna2aa1n03x5               g219(.a(new_n105), .b(new_n108), .c(new_n111), .out0(\s[3] ));
  oai012aa1n02x5               g220(.a(new_n108), .b(new_n105), .c(new_n107), .o1(new_n316));
  xnrb03aa1n02x5               g221(.a(new_n316), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnbna2aa1n03x5               g222(.a(new_n119), .b(new_n110), .c(new_n112), .out0(\s[5] ));
  nanp02aa1n02x5               g223(.a(new_n110), .b(new_n112), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n123), .b(new_n319), .c(new_n119), .o1(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[5] ), .c(new_n121), .out0(\s[6] ));
  norb02aa1n02x5               g226(.a(new_n116), .b(new_n115), .out0(new_n322));
  nanp02aa1n02x5               g227(.a(new_n320), .b(new_n118), .o1(new_n323));
  oai112aa1n02x5               g228(.a(new_n323), .b(new_n322), .c(new_n122), .d(new_n121), .o1(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n322), .b(new_n323), .c(new_n121), .d(new_n122), .o1(new_n325));
  norb02aa1n02x5               g230(.a(new_n324), .b(new_n325), .out0(\s[7] ));
  norb02aa1n02x5               g231(.a(new_n114), .b(new_n113), .out0(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n327), .b(new_n324), .c(new_n125), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


