// Benchmark "adder" written by ABC on Thu Jul 18 10:49:18 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n329, new_n331, new_n332, new_n333, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oao003aa1n02x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n101));
  norp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano23aa1n02x4               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  oa0012aa1n02x5               g011(.a(new_n103), .b(new_n104), .c(new_n102), .o(new_n107));
  nand02aa1d04x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor042aa1n03x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand02aa1n03x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb03aa1d18x5               g015(.a(new_n109), .b(new_n110), .c(new_n108), .out0(new_n111));
  xnrc02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .out0(new_n112));
  inv000aa1d42x5               g017(.a(\a[5] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[4] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(new_n114), .b(new_n113), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  oai112aa1n02x5               g021(.a(new_n115), .b(new_n116), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  nor043aa1n03x5               g022(.a(new_n117), .b(new_n111), .c(new_n112), .o1(new_n118));
  aoai13aa1n02x5               g023(.a(new_n118), .b(new_n107), .c(new_n101), .d(new_n106), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n111), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\a[6] ), .o1(new_n121));
  aboi22aa1n06x5               g026(.a(\b[5] ), .b(new_n121), .c(new_n113), .d(new_n114), .out0(new_n122));
  norp02aa1n02x5               g027(.a(new_n112), .b(new_n122), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\a[8] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[7] ), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(new_n124), .b(new_n125), .c(new_n109), .o1(new_n126));
  aobi12aa1n02x5               g031(.a(new_n126), .b(new_n123), .c(new_n120), .out0(new_n127));
  nanp02aa1n06x5               g032(.a(new_n119), .b(new_n127), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  aoi012aa1n02x5               g034(.a(new_n97), .b(new_n128), .c(new_n129), .o1(new_n130));
  xnrb03aa1n02x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand22aa1n03x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  norp02aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  nano23aa1n03x7               g038(.a(new_n97), .b(new_n133), .c(new_n132), .d(new_n129), .out0(new_n134));
  oai022aa1n02x5               g039(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n135));
  ao0022aa1n03x5               g040(.a(new_n128), .b(new_n134), .c(new_n135), .d(new_n132), .o(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  aoi022aa1n02x5               g042(.a(new_n128), .b(new_n134), .c(new_n132), .d(new_n135), .o1(new_n138));
  oaoi03aa1n02x5               g043(.a(\a[11] ), .b(\b[10] ), .c(new_n138), .o1(new_n139));
  xorb03aa1n02x5               g044(.a(new_n139), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nona23aa1n02x4               g045(.a(new_n132), .b(new_n129), .c(new_n97), .d(new_n133), .out0(new_n141));
  nor002aa1n02x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  inv000aa1d42x5               g049(.a(\a[12] ), .o1(new_n145));
  inv000aa1d42x5               g050(.a(\b[11] ), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(new_n146), .b(new_n145), .o1(new_n147));
  nanp02aa1n02x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  norp03aa1n02x5               g054(.a(new_n141), .b(new_n144), .c(new_n149), .o1(new_n150));
  nanb03aa1n02x5               g055(.a(new_n142), .b(new_n143), .c(new_n132), .out0(new_n151));
  nanp03aa1n02x5               g056(.a(new_n135), .b(new_n147), .c(new_n148), .o1(new_n152));
  oaoi03aa1n02x5               g057(.a(new_n145), .b(new_n146), .c(new_n142), .o1(new_n153));
  tech160nm_fioai012aa1n03p5x5 g058(.a(new_n153), .b(new_n152), .c(new_n151), .o1(new_n154));
  nor042aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n154), .c(new_n128), .d(new_n150), .o1(new_n158));
  aoi112aa1n02x5               g063(.a(new_n157), .b(new_n154), .c(new_n128), .d(new_n150), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(\s[13] ));
  tech160nm_fioai012aa1n03p5x5 g065(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1n09x5               g069(.a(new_n155), .b(new_n163), .c(new_n164), .d(new_n156), .out0(new_n165));
  oa0012aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n155), .o(new_n166));
  aoi012aa1n02x5               g071(.a(new_n166), .b(new_n154), .c(new_n165), .o1(new_n167));
  nona22aa1n02x4               g072(.a(new_n134), .b(new_n144), .c(new_n149), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n165), .o1(new_n169));
  nona22aa1n02x4               g074(.a(new_n128), .b(new_n168), .c(new_n169), .out0(new_n170));
  nanp02aa1n02x5               g075(.a(new_n170), .b(new_n167), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  aoi012aa1n02x5               g079(.a(new_n173), .b(new_n171), .c(new_n174), .o1(new_n175));
  xnrb03aa1n02x5               g080(.a(new_n175), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  oaoi03aa1n02x5               g081(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n177));
  nona23aa1n02x4               g082(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n178));
  oabi12aa1n02x5               g083(.a(new_n107), .b(new_n177), .c(new_n178), .out0(new_n179));
  oai013aa1n03x4               g084(.a(new_n126), .b(new_n111), .c(new_n112), .d(new_n122), .o1(new_n180));
  norp02aa1n02x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nanp02aa1n02x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nano23aa1n02x4               g087(.a(new_n173), .b(new_n181), .c(new_n182), .d(new_n174), .out0(new_n183));
  nano22aa1n02x4               g088(.a(new_n168), .b(new_n165), .c(new_n183), .out0(new_n184));
  aoai13aa1n04x5               g089(.a(new_n184), .b(new_n180), .c(new_n179), .d(new_n118), .o1(new_n185));
  aoai13aa1n04x5               g090(.a(new_n183), .b(new_n166), .c(new_n154), .d(new_n165), .o1(new_n186));
  oai012aa1n02x5               g091(.a(new_n182), .b(new_n181), .c(new_n173), .o1(new_n187));
  nand23aa1n04x5               g092(.a(new_n185), .b(new_n186), .c(new_n187), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nanp03aa1n02x5               g094(.a(new_n150), .b(new_n165), .c(new_n183), .o1(new_n190));
  tech160nm_fiaoi012aa1n02p5x5 g095(.a(new_n190), .b(new_n119), .c(new_n127), .o1(new_n191));
  nano22aa1n03x7               g096(.a(new_n191), .b(new_n186), .c(new_n187), .out0(new_n192));
  oaoi03aa1n02x5               g097(.a(\a[17] ), .b(\b[16] ), .c(new_n192), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv000aa1d42x5               g099(.a(\a[17] ), .o1(new_n195));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  xroi22aa1d06x4               g101(.a(new_n195), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n197));
  inv000aa1d42x5               g102(.a(\b[17] ), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  oao003aa1n02x5               g104(.a(new_n196), .b(new_n198), .c(new_n199), .carry(new_n200));
  tech160nm_fiaoi012aa1n05x5   g105(.a(new_n200), .b(new_n188), .c(new_n197), .o1(new_n201));
  inv000aa1d42x5               g106(.a(\a[19] ), .o1(new_n202));
  nanb02aa1n03x5               g107(.a(\b[18] ), .b(new_n202), .out0(new_n203));
  nand02aa1d10x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n201), .b(new_n204), .c(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g111(.a(new_n197), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n200), .o1(new_n208));
  oaih12aa1n02x5               g113(.a(new_n208), .b(new_n192), .c(new_n207), .o1(new_n209));
  norp02aa1n04x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  tech160nm_fixorc02aa1n05x5   g115(.a(\a[20] ), .b(\b[19] ), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n212), .b(new_n210), .c(new_n209), .d(new_n204), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n204), .o1(new_n214));
  oai112aa1n02x5               g119(.a(new_n211), .b(new_n203), .c(new_n201), .d(new_n214), .o1(new_n215));
  nanp02aa1n03x5               g120(.a(new_n213), .b(new_n215), .o1(\s[20] ));
  nona23aa1d16x5               g121(.a(new_n197), .b(new_n211), .c(new_n214), .d(new_n210), .out0(new_n217));
  oai112aa1n04x5               g122(.a(new_n203), .b(new_n204), .c(new_n198), .d(new_n196), .o1(new_n218));
  oai022aa1n02x5               g123(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(\a[20] ), .o1(new_n220));
  inv000aa1d42x5               g125(.a(\b[19] ), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(new_n221), .b(new_n220), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nanp03aa1n02x5               g128(.a(new_n219), .b(new_n222), .c(new_n223), .o1(new_n224));
  oaoi03aa1n03x5               g129(.a(new_n220), .b(new_n221), .c(new_n210), .o1(new_n225));
  oai012aa1n12x5               g130(.a(new_n225), .b(new_n224), .c(new_n218), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  tech160nm_fioai012aa1n05x5   g132(.a(new_n227), .b(new_n192), .c(new_n217), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n02x5               g138(.a(new_n233), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n217), .o1(new_n235));
  aoai13aa1n02x5               g140(.a(new_n231), .b(new_n226), .c(new_n188), .d(new_n235), .o1(new_n236));
  nona22aa1n02x4               g141(.a(new_n236), .b(new_n233), .c(new_n230), .out0(new_n237));
  nanp02aa1n02x5               g142(.a(new_n234), .b(new_n237), .o1(\s[22] ));
  inv000aa1d42x5               g143(.a(\a[21] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\a[22] ), .o1(new_n240));
  xroi22aa1d04x5               g145(.a(new_n239), .b(\b[20] ), .c(new_n240), .d(\b[21] ), .out0(new_n241));
  norb02aa1n03x5               g146(.a(new_n241), .b(new_n217), .out0(new_n242));
  inv000aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(\b[20] ), .b(new_n239), .out0(new_n244));
  oaoi03aa1n02x5               g149(.a(\a[22] ), .b(\b[21] ), .c(new_n244), .o1(new_n245));
  tech160nm_fiaoi012aa1n03p5x5 g150(.a(new_n245), .b(new_n226), .c(new_n241), .o1(new_n246));
  oai012aa1n04x7               g151(.a(new_n246), .b(new_n192), .c(new_n243), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  tech160nm_fixorc02aa1n04x5   g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n249), .c(new_n247), .d(new_n250), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n246), .o1(new_n254));
  aoai13aa1n02x5               g159(.a(new_n250), .b(new_n254), .c(new_n188), .d(new_n242), .o1(new_n255));
  nona22aa1n02x4               g160(.a(new_n255), .b(new_n252), .c(new_n249), .out0(new_n256));
  nanp02aa1n02x5               g161(.a(new_n253), .b(new_n256), .o1(\s[24] ));
  and002aa1n02x5               g162(.a(new_n251), .b(new_n250), .o(new_n258));
  nano22aa1n03x7               g163(.a(new_n217), .b(new_n258), .c(new_n241), .out0(new_n259));
  inv020aa1n03x5               g164(.a(new_n259), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n258), .b(new_n245), .c(new_n226), .d(new_n241), .o1(new_n261));
  oai022aa1n02x5               g166(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n262));
  aob012aa1n02x5               g167(.a(new_n262), .b(\b[23] ), .c(\a[24] ), .out0(new_n263));
  nand02aa1n06x5               g168(.a(new_n261), .b(new_n263), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  oai012aa1n04x7               g170(.a(new_n265), .b(new_n192), .c(new_n260), .o1(new_n266));
  xorb03aa1n02x5               g171(.a(new_n266), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g172(.a(\b[24] ), .b(\a[25] ), .o1(new_n268));
  xorc02aa1n02x5               g173(.a(\a[25] ), .b(\b[24] ), .out0(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[25] ), .b(\a[26] ), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n268), .c(new_n266), .d(new_n269), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n269), .b(new_n264), .c(new_n188), .d(new_n259), .o1(new_n272));
  nona22aa1n02x4               g177(.a(new_n272), .b(new_n270), .c(new_n268), .out0(new_n273));
  nanp02aa1n03x5               g178(.a(new_n271), .b(new_n273), .o1(\s[26] ));
  norb02aa1n03x5               g179(.a(new_n269), .b(new_n270), .out0(new_n275));
  nano32aa1d12x5               g180(.a(new_n217), .b(new_n275), .c(new_n241), .d(new_n258), .out0(new_n276));
  inv020aa1n03x5               g181(.a(new_n276), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(\b[25] ), .b(\a[26] ), .o1(new_n278));
  oai022aa1n02x5               g183(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n279));
  aoi022aa1n03x5               g184(.a(new_n264), .b(new_n275), .c(new_n278), .d(new_n279), .o1(new_n280));
  tech160nm_fioai012aa1n03p5x5 g185(.a(new_n280), .b(new_n192), .c(new_n277), .o1(new_n281));
  xorb03aa1n02x5               g186(.a(new_n281), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n04x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  xorc02aa1n02x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  tech160nm_fixorc02aa1n02p5x5 g189(.a(\a[28] ), .b(\b[27] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n281), .d(new_n284), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n275), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(new_n279), .b(new_n278), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n288), .c(new_n261), .d(new_n263), .o1(new_n290));
  aoai13aa1n02x5               g195(.a(new_n284), .b(new_n290), .c(new_n188), .d(new_n276), .o1(new_n291));
  nona22aa1n02x5               g196(.a(new_n291), .b(new_n286), .c(new_n283), .out0(new_n292));
  nanp02aa1n03x5               g197(.a(new_n287), .b(new_n292), .o1(\s[28] ));
  and002aa1n02x5               g198(.a(new_n285), .b(new_n284), .o(new_n294));
  aoai13aa1n06x5               g199(.a(new_n294), .b(new_n290), .c(new_n188), .d(new_n276), .o1(new_n295));
  inv000aa1d42x5               g200(.a(\a[28] ), .o1(new_n296));
  inv000aa1d42x5               g201(.a(\b[27] ), .o1(new_n297));
  oaoi03aa1n09x5               g202(.a(new_n296), .b(new_n297), .c(new_n283), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n295), .c(new_n298), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n298), .o1(new_n302));
  nona22aa1n02x5               g207(.a(new_n295), .b(new_n302), .c(new_n299), .out0(new_n303));
  norb02aa1n03x4               g208(.a(new_n303), .b(new_n301), .out0(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g210(.a(new_n300), .b(new_n284), .c(new_n285), .out0(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n290), .c(new_n188), .d(new_n276), .o1(new_n307));
  tech160nm_fioaoi03aa1n03p5x5 g212(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .o1(new_n308));
  inv000aa1n03x5               g213(.a(new_n308), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .out0(new_n310));
  inv000aa1d42x5               g215(.a(new_n310), .o1(new_n311));
  tech160nm_fiaoi012aa1n03p5x5 g216(.a(new_n311), .b(new_n307), .c(new_n309), .o1(new_n312));
  nona22aa1n02x5               g217(.a(new_n307), .b(new_n308), .c(new_n310), .out0(new_n313));
  norb02aa1n03x4               g218(.a(new_n313), .b(new_n312), .out0(\s[30] ));
  nano32aa1n02x4               g219(.a(new_n311), .b(new_n299), .c(new_n285), .d(new_n284), .out0(new_n315));
  aoai13aa1n06x5               g220(.a(new_n315), .b(new_n290), .c(new_n188), .d(new_n276), .o1(new_n316));
  tech160nm_fioaoi03aa1n03p5x5 g221(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n317), .o1(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[30] ), .b(\a[31] ), .out0(new_n319));
  tech160nm_fiaoi012aa1n03p5x5 g224(.a(new_n319), .b(new_n316), .c(new_n318), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n319), .o1(new_n321));
  nona22aa1n02x5               g226(.a(new_n316), .b(new_n317), .c(new_n321), .out0(new_n322));
  norb02aa1n03x4               g227(.a(new_n322), .b(new_n320), .out0(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n177), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g229(.a(\a[3] ), .b(\b[2] ), .c(new_n177), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n179), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g232(.a(\b[5] ), .b(new_n121), .out0(new_n328));
  oaoi03aa1n02x5               g233(.a(new_n113), .b(new_n114), .c(new_n179), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n329), .b(new_n108), .c(new_n328), .out0(\s[6] ));
  nano22aa1n02x4               g235(.a(new_n329), .b(new_n108), .c(new_n328), .out0(new_n331));
  inv000aa1d42x5               g236(.a(new_n122), .o1(new_n332));
  aoi013aa1n02x4               g237(.a(new_n332), .b(new_n179), .c(new_n115), .d(new_n116), .o1(new_n333));
  oaib12aa1n02x5               g238(.a(new_n328), .b(new_n109), .c(new_n110), .out0(new_n334));
  oa0022aa1n02x5               g239(.a(new_n331), .b(new_n334), .c(new_n111), .d(new_n333), .o(\s[7] ));
  oai022aa1n02x5               g240(.a(new_n333), .b(new_n111), .c(\b[6] ), .d(\a[7] ), .o1(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g242(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


