// Benchmark "adder" written by ABC on Wed Jul 17 16:35:06 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n309, new_n312,
    new_n314, new_n316;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nand02aa1d06x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  aoi012aa1n12x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n101));
  inv000aa1n02x5               g006(.a(new_n101), .o1(new_n102));
  nor042aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano23aa1n03x5               g011(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n107));
  nand42aa1n02x5               g012(.a(new_n107), .b(new_n102), .o1(new_n108));
  aoi012aa1n02x7               g013(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n109));
  norp02aa1n04x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nanp02aa1n03x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor022aa1n04x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nano23aa1n06x5               g018(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n114));
  nand42aa1n06x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor042aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor042aa1n03x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nand42aa1n03x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nano23aa1n03x7               g023(.a(new_n117), .b(new_n116), .c(new_n118), .d(new_n115), .out0(new_n119));
  nand02aa1n02x5               g024(.a(new_n119), .b(new_n114), .o1(new_n120));
  aoi012aa1n09x5               g025(.a(new_n116), .b(new_n117), .c(new_n115), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n121), .o1(new_n122));
  tech160nm_fiao0012aa1n02p5x5 g027(.a(new_n110), .b(new_n112), .c(new_n111), .o(new_n123));
  aoi012aa1n06x5               g028(.a(new_n123), .b(new_n114), .c(new_n122), .o1(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n120), .c(new_n108), .d(new_n109), .o1(new_n125));
  nand42aa1n03x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  aoi012aa1n02x5               g031(.a(new_n97), .b(new_n125), .c(new_n126), .o1(new_n127));
  xnrb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1n08x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nano23aa1n06x5               g035(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n126), .out0(new_n131));
  aoi012aa1d18x5               g036(.a(new_n129), .b(new_n97), .c(new_n130), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  tech160nm_fixorc02aa1n02p5x5 g038(.a(\a[11] ), .b(\b[10] ), .out0(new_n134));
  aoai13aa1n03x5               g039(.a(new_n134), .b(new_n133), .c(new_n125), .d(new_n131), .o1(new_n135));
  aoi112aa1n02x5               g040(.a(new_n134), .b(new_n133), .c(new_n125), .d(new_n131), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(\s[11] ));
  orn002aa1n02x5               g042(.a(\a[11] ), .b(\b[10] ), .o(new_n138));
  tech160nm_fixorc02aa1n02p5x5 g043(.a(\a[12] ), .b(\b[11] ), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n135), .c(new_n138), .out0(\s[12] ));
  xnrc02aa1n02x5               g045(.a(\b[10] ), .b(\a[11] ), .out0(new_n141));
  xnrc02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .out0(new_n142));
  oao003aa1n02x5               g047(.a(\a[12] ), .b(\b[11] ), .c(new_n138), .carry(new_n143));
  oai013aa1n06x5               g048(.a(new_n143), .b(new_n141), .c(new_n142), .d(new_n132), .o1(new_n144));
  and003aa1n02x5               g049(.a(new_n131), .b(new_n139), .c(new_n134), .o(new_n145));
  tech160nm_fiaoi012aa1n05x5   g050(.a(new_n144), .b(new_n125), .c(new_n145), .o1(new_n146));
  tech160nm_fixorc02aa1n03p5x5 g051(.a(\a[13] ), .b(\b[12] ), .out0(new_n147));
  xnrc02aa1n02x5               g052(.a(new_n146), .b(new_n147), .out0(\s[13] ));
  oaoi03aa1n03x5               g053(.a(\a[13] ), .b(\b[12] ), .c(new_n146), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n04x5               g055(.a(\b[14] ), .b(\a[15] ), .o1(new_n151));
  nand42aa1n08x5               g056(.a(\b[14] ), .b(\a[15] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  tech160nm_fixorc02aa1n03p5x5 g058(.a(\a[14] ), .b(\b[13] ), .out0(new_n154));
  and002aa1n02x5               g059(.a(new_n154), .b(new_n147), .o(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n144), .c(new_n125), .d(new_n145), .o1(new_n156));
  inv000aa1d42x5               g061(.a(\a[14] ), .o1(new_n157));
  inv000aa1d42x5               g062(.a(\b[13] ), .o1(new_n158));
  norp02aa1n02x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  oaoi03aa1n02x5               g064(.a(new_n157), .b(new_n158), .c(new_n159), .o1(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n153), .b(new_n156), .c(new_n160), .out0(\s[15] ));
  nand42aa1n03x5               g066(.a(new_n156), .b(new_n160), .o1(new_n162));
  nor042aa1n02x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nand42aa1n03x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n151), .c(new_n162), .d(new_n152), .o1(new_n166));
  aob012aa1n03x5               g071(.a(new_n153), .b(new_n156), .c(new_n160), .out0(new_n167));
  nona22aa1n02x5               g072(.a(new_n167), .b(new_n165), .c(new_n151), .out0(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n166), .o1(\s[16] ));
  nona23aa1n02x4               g074(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n170));
  tech160nm_fioai012aa1n05x5   g075(.a(new_n109), .b(new_n170), .c(new_n101), .o1(new_n171));
  nona23aa1n02x4               g076(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n172));
  norb02aa1n02x7               g077(.a(new_n119), .b(new_n172), .out0(new_n173));
  oabi12aa1n02x5               g078(.a(new_n123), .b(new_n172), .c(new_n121), .out0(new_n174));
  nano23aa1n06x5               g079(.a(new_n151), .b(new_n163), .c(new_n164), .d(new_n152), .out0(new_n175));
  nand43aa1n03x5               g080(.a(new_n175), .b(new_n147), .c(new_n154), .o1(new_n176));
  nano32aa1n03x7               g081(.a(new_n176), .b(new_n139), .c(new_n131), .d(new_n134), .out0(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n174), .c(new_n171), .d(new_n173), .o1(new_n178));
  oao003aa1n02x5               g083(.a(new_n157), .b(new_n158), .c(new_n159), .carry(new_n179));
  tech160nm_fiao0012aa1n02p5x5 g084(.a(new_n163), .b(new_n151), .c(new_n164), .o(new_n180));
  tech160nm_fiaoi012aa1n03p5x5 g085(.a(new_n180), .b(new_n175), .c(new_n179), .o1(new_n181));
  inv000aa1n02x5               g086(.a(new_n181), .o1(new_n182));
  aoib12aa1n12x5               g087(.a(new_n182), .b(new_n144), .c(new_n176), .out0(new_n183));
  nanp02aa1n06x5               g088(.a(new_n178), .b(new_n183), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g090(.a(\a[18] ), .o1(new_n186));
  inv040aa1d30x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  oaoi03aa1n03x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n186), .out0(\s[18] ));
  xroi22aa1d06x4               g095(.a(new_n187), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  nor002aa1n03x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  aoi112aa1n09x5               g098(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n194));
  nor042aa1n04x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  aoai13aa1n06x5               g100(.a(new_n195), .b(new_n192), .c(new_n178), .d(new_n183), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n12x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nand02aa1d06x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nor002aa1d32x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand02aa1d28x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n15x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n204), .b(new_n199), .c(new_n196), .d(new_n200), .o1(new_n205));
  norb02aa1n12x5               g110(.a(new_n200), .b(new_n199), .out0(new_n206));
  nanp02aa1n02x5               g111(.a(new_n196), .b(new_n206), .o1(new_n207));
  nona22aa1n02x5               g112(.a(new_n207), .b(new_n204), .c(new_n199), .out0(new_n208));
  nanp02aa1n03x5               g113(.a(new_n208), .b(new_n205), .o1(\s[20] ));
  nona23aa1d18x5               g114(.a(new_n202), .b(new_n200), .c(new_n199), .d(new_n201), .out0(new_n210));
  aoi012aa1n06x5               g115(.a(new_n201), .b(new_n199), .c(new_n202), .o1(new_n211));
  oai012aa1n12x5               g116(.a(new_n211), .b(new_n210), .c(new_n195), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  nanb02aa1n06x5               g118(.a(new_n210), .b(new_n191), .out0(new_n214));
  aoai13aa1n04x5               g119(.a(new_n213), .b(new_n214), .c(new_n178), .d(new_n183), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  xorc02aa1n12x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[21] ), .b(\a[22] ), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n215), .d(new_n218), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(new_n215), .b(new_n218), .o1(new_n221));
  nona22aa1n02x5               g126(.a(new_n221), .b(new_n219), .c(new_n217), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n222), .b(new_n220), .o1(\s[22] ));
  oai112aa1n06x5               g128(.a(new_n206), .b(new_n203), .c(new_n194), .d(new_n193), .o1(new_n224));
  nanb02aa1n03x5               g129(.a(new_n219), .b(new_n218), .out0(new_n225));
  inv000aa1d42x5               g130(.a(\a[22] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\b[21] ), .o1(new_n227));
  oaoi03aa1n12x5               g132(.a(new_n226), .b(new_n227), .c(new_n217), .o1(new_n228));
  aoai13aa1n12x5               g133(.a(new_n228), .b(new_n225), .c(new_n224), .d(new_n211), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  nona23aa1n08x5               g135(.a(new_n191), .b(new_n218), .c(new_n219), .d(new_n210), .out0(new_n231));
  aoai13aa1n04x5               g136(.a(new_n230), .b(new_n231), .c(new_n178), .d(new_n183), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  xorc02aa1n02x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  xorc02aa1n12x5               g140(.a(\a[24] ), .b(\b[23] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n234), .c(new_n232), .d(new_n235), .o1(new_n238));
  nanp02aa1n02x5               g143(.a(new_n232), .b(new_n235), .o1(new_n239));
  nona22aa1n02x5               g144(.a(new_n239), .b(new_n237), .c(new_n234), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[24] ));
  nanb03aa1n02x5               g146(.a(new_n132), .b(new_n139), .c(new_n134), .out0(new_n242));
  aoai13aa1n03x5               g147(.a(new_n181), .b(new_n176), .c(new_n242), .d(new_n143), .o1(new_n243));
  norb02aa1n06x4               g148(.a(new_n218), .b(new_n219), .out0(new_n244));
  and002aa1n02x5               g149(.a(new_n236), .b(new_n235), .o(new_n245));
  nano22aa1n03x7               g150(.a(new_n214), .b(new_n245), .c(new_n244), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n243), .c(new_n125), .d(new_n177), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n228), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n245), .b(new_n248), .c(new_n212), .d(new_n244), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\a[24] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[23] ), .o1(new_n251));
  tech160nm_fioaoi03aa1n03p5x5 g156(.a(new_n250), .b(new_n251), .c(new_n234), .o1(new_n252));
  nanp02aa1n02x5               g157(.a(new_n249), .b(new_n252), .o1(new_n253));
  nanb02aa1n03x5               g158(.a(new_n253), .b(new_n247), .out0(new_n254));
  xorb03aa1n02x5               g159(.a(new_n254), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g160(.a(\b[24] ), .b(\a[25] ), .o1(new_n256));
  tech160nm_fixorc02aa1n03p5x5 g161(.a(\a[25] ), .b(\b[24] ), .out0(new_n257));
  xorc02aa1n12x5               g162(.a(\a[26] ), .b(\b[25] ), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n256), .c(new_n254), .d(new_n257), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n257), .b(new_n253), .c(new_n184), .d(new_n246), .o1(new_n261));
  nona22aa1n02x5               g166(.a(new_n261), .b(new_n259), .c(new_n256), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n260), .b(new_n262), .o1(\s[26] ));
  and002aa1n06x5               g168(.a(new_n258), .b(new_n257), .o(new_n264));
  nano22aa1n03x7               g169(.a(new_n231), .b(new_n245), .c(new_n264), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n243), .c(new_n125), .d(new_n177), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n252), .o1(new_n267));
  aoai13aa1n04x5               g172(.a(new_n264), .b(new_n267), .c(new_n229), .d(new_n245), .o1(new_n268));
  aoi112aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n269));
  oab012aa1n02x4               g174(.a(new_n269), .b(\a[26] ), .c(\b[25] ), .out0(new_n270));
  nand43aa1n03x5               g175(.a(new_n266), .b(new_n268), .c(new_n270), .o1(new_n271));
  xorb03aa1n03x5               g176(.a(new_n271), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[27] ), .b(\a[28] ), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n276));
  aobi12aa1n06x5               g181(.a(new_n265), .b(new_n178), .c(new_n183), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n264), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n270), .b(new_n278), .c(new_n249), .d(new_n252), .o1(new_n279));
  oaih12aa1n02x5               g184(.a(new_n274), .b(new_n279), .c(new_n277), .o1(new_n280));
  nona22aa1n02x5               g185(.a(new_n280), .b(new_n275), .c(new_n273), .out0(new_n281));
  nanp02aa1n03x5               g186(.a(new_n276), .b(new_n281), .o1(\s[28] ));
  norb02aa1n02x5               g187(.a(new_n274), .b(new_n275), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n283), .b(new_n279), .c(new_n277), .o1(new_n284));
  aob012aa1n03x5               g189(.a(new_n273), .b(\b[27] ), .c(\a[28] ), .out0(new_n285));
  oa0012aa1n12x5               g190(.a(new_n285), .b(\b[27] ), .c(\a[28] ), .o(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  nona22aa1n02x5               g193(.a(new_n284), .b(new_n287), .c(new_n288), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n288), .b(new_n287), .c(new_n271), .d(new_n283), .o1(new_n290));
  nanp02aa1n03x5               g195(.a(new_n290), .b(new_n289), .o1(\s[29] ));
  xorb03aa1n02x5               g196(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g197(.a(new_n274), .b(new_n288), .c(new_n275), .out0(new_n293));
  oaoi03aa1n09x5               g198(.a(\a[29] ), .b(\b[28] ), .c(new_n286), .o1(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n271), .d(new_n293), .o1(new_n296));
  oaih12aa1n02x5               g201(.a(new_n293), .b(new_n279), .c(new_n277), .o1(new_n297));
  nona22aa1n02x5               g202(.a(new_n297), .b(new_n294), .c(new_n295), .out0(new_n298));
  nanp02aa1n03x5               g203(.a(new_n296), .b(new_n298), .o1(\s[30] ));
  norb02aa1n02x5               g204(.a(new_n293), .b(new_n295), .out0(new_n300));
  oaih12aa1n02x5               g205(.a(new_n300), .b(new_n279), .c(new_n277), .o1(new_n301));
  nanb02aa1n02x5               g206(.a(new_n295), .b(new_n294), .out0(new_n302));
  oai012aa1n02x5               g207(.a(new_n302), .b(\b[29] ), .c(\a[30] ), .o1(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  nona22aa1n02x5               g209(.a(new_n301), .b(new_n303), .c(new_n304), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n304), .b(new_n303), .c(new_n271), .d(new_n300), .o1(new_n306));
  nanp02aa1n03x5               g211(.a(new_n306), .b(new_n305), .o1(\s[31] ));
  xnrb03aa1n02x5               g212(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g213(.a(\a[3] ), .b(\b[2] ), .c(new_n101), .o1(new_n309));
  xorb03aa1n02x5               g214(.a(new_n309), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g215(.a(new_n171), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g216(.a(new_n117), .b(new_n171), .c(new_n118), .o1(new_n312));
  xnrb03aa1n02x5               g217(.a(new_n312), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aob012aa1n02x5               g218(.a(new_n121), .b(new_n171), .c(new_n119), .out0(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g220(.a(new_n112), .b(new_n314), .c(new_n113), .o1(new_n316));
  xnrb03aa1n02x5               g221(.a(new_n316), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g222(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


