// Benchmark "adder" written by ABC on Thu Jul 18 05:13:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n330,
    new_n331, new_n333, new_n334, new_n335, new_n337, new_n338, new_n339,
    new_n341, new_n342, new_n343, new_n344, new_n346, new_n347, new_n348,
    new_n349, new_n351, new_n352, new_n354, new_n355, new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixnrc02aa1n04x5   g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\a[9] ), .b(new_n98), .out0(new_n99));
  and002aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o(new_n100));
  oaoi03aa1n12x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  xorc02aa1n12x5               g006(.a(\a[3] ), .b(\b[2] ), .out0(new_n102));
  oaih22aa1d12x5               g007(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  aoi012aa1d24x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .o1(new_n104));
  nor042aa1n09x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nand42aa1n10x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand42aa1n08x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nano22aa1d15x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .out0(new_n108));
  nand42aa1n16x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  oai012aa1n12x5               g014(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .o1(new_n110));
  aoi022aa1n06x5               g015(.a(\b[5] ), .b(\a[6] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n111));
  oai022aa1n02x5               g016(.a(\a[6] ), .b(\b[5] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n112));
  nona23aa1n12x5               g017(.a(new_n108), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n113));
  nor042aa1n09x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  inv040aa1n04x5               g019(.a(new_n114), .o1(new_n115));
  tech160nm_fioaoi03aa1n03p5x5 g020(.a(\a[6] ), .b(\b[5] ), .c(new_n115), .o1(new_n116));
  nor042aa1n03x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nano23aa1n09x5               g022(.a(new_n117), .b(new_n105), .c(new_n106), .d(new_n107), .out0(new_n118));
  tech160nm_fioai012aa1n05x5   g023(.a(new_n106), .b(new_n117), .c(new_n105), .o1(new_n119));
  aobi12aa1n09x5               g024(.a(new_n119), .b(new_n118), .c(new_n116), .out0(new_n120));
  oai012aa1d24x5               g025(.a(new_n120), .b(new_n104), .c(new_n113), .o1(new_n121));
  oaib12aa1n09x5               g026(.a(new_n121), .b(new_n98), .c(\a[9] ), .out0(new_n122));
  xobna2aa1n03x5               g027(.a(new_n97), .b(new_n122), .c(new_n99), .out0(\s[10] ));
  nand42aa1d28x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  nor002aa1n20x5               g029(.a(\b[10] ), .b(\a[11] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n124), .b(new_n125), .out0(new_n126));
  oai022aa1n04x7               g031(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  aboi22aa1n03x5               g032(.a(new_n127), .b(new_n122), .c(\b[9] ), .d(\a[10] ), .out0(new_n128));
  aoi022aa1n06x5               g033(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n125), .out0(new_n130));
  oaib12aa1n02x5               g035(.a(new_n130), .b(new_n127), .c(new_n122), .out0(new_n131));
  oa0012aa1n02x5               g036(.a(new_n131), .b(new_n128), .c(new_n126), .o(\s[11] ));
  inv000aa1d42x5               g037(.a(new_n125), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  nand42aa1d28x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  nor002aa1n03x5               g041(.a(new_n134), .b(new_n125), .o1(new_n137));
  nanp03aa1n02x5               g042(.a(new_n131), .b(new_n135), .c(new_n137), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n136), .c(new_n133), .d(new_n131), .o1(\s[12] ));
  nano23aa1d15x5               g044(.a(new_n134), .b(new_n125), .c(new_n135), .d(new_n124), .out0(new_n140));
  xorc02aa1n12x5               g045(.a(\a[9] ), .b(\b[8] ), .out0(new_n141));
  nanb03aa1d24x5               g046(.a(new_n97), .b(new_n140), .c(new_n141), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  nanp02aa1n03x5               g048(.a(new_n121), .b(new_n143), .o1(new_n144));
  aob012aa1n03x5               g049(.a(new_n137), .b(new_n127), .c(new_n129), .out0(new_n145));
  nanp02aa1n02x5               g050(.a(new_n145), .b(new_n135), .o1(new_n146));
  tech160nm_fixorc02aa1n03p5x5 g051(.a(\a[13] ), .b(\b[12] ), .out0(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n146), .out0(\s[13] ));
  inv040aa1d32x5               g053(.a(\a[13] ), .o1(new_n149));
  inv000aa1d42x5               g054(.a(\b[12] ), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n150), .b(new_n149), .o1(new_n151));
  nanp02aa1n03x5               g056(.a(new_n144), .b(new_n146), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(new_n152), .b(new_n147), .o1(new_n153));
  xorc02aa1n02x5               g058(.a(\a[14] ), .b(\b[13] ), .out0(new_n154));
  nand02aa1d04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  oai022aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n156));
  nanb03aa1n02x5               g061(.a(new_n156), .b(new_n153), .c(new_n155), .out0(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n154), .c(new_n151), .d(new_n153), .o1(\s[14] ));
  and002aa1n02x5               g063(.a(new_n154), .b(new_n147), .o(new_n159));
  oaoi03aa1n02x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n151), .o1(new_n160));
  nor042aa1n06x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(new_n161), .b(new_n162), .out0(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n160), .c(new_n152), .d(new_n159), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n164), .b(new_n160), .c(new_n152), .d(new_n159), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(\s[15] ));
  inv000aa1d42x5               g072(.a(new_n161), .o1(new_n168));
  nor042aa1n06x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n169), .o1(new_n172));
  oai112aa1n02x5               g077(.a(new_n172), .b(new_n170), .c(\b[14] ), .d(\a[15] ), .o1(new_n173));
  nanb02aa1n03x5               g078(.a(new_n173), .b(new_n165), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n171), .c(new_n168), .d(new_n165), .o1(\s[16] ));
  nano23aa1n06x5               g080(.a(new_n161), .b(new_n169), .c(new_n170), .d(new_n162), .out0(new_n176));
  nano32aa1d12x5               g081(.a(new_n142), .b(new_n176), .c(new_n147), .d(new_n154), .out0(new_n177));
  nanp02aa1n06x5               g082(.a(new_n121), .b(new_n177), .o1(new_n178));
  nano22aa1n03x5               g083(.a(new_n169), .b(new_n162), .c(new_n170), .out0(new_n179));
  oai022aa1n02x5               g084(.a(new_n149), .b(new_n150), .c(\b[13] ), .d(\a[14] ), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n155), .b(\b[14] ), .c(\a[15] ), .o1(new_n181));
  nano23aa1n02x5               g086(.a(new_n180), .b(new_n181), .c(new_n151), .d(new_n135), .out0(new_n182));
  nand23aa1n02x5               g087(.a(new_n182), .b(new_n145), .c(new_n179), .o1(new_n183));
  aoi022aa1n02x5               g088(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n184));
  aoai13aa1n03x5               g089(.a(new_n184), .b(new_n161), .c(new_n156), .d(new_n155), .o1(new_n185));
  nand23aa1n06x5               g090(.a(new_n183), .b(new_n172), .c(new_n185), .o1(new_n186));
  nanb02aa1n09x5               g091(.a(new_n186), .b(new_n178), .out0(new_n187));
  xorc02aa1n12x5               g092(.a(\a[17] ), .b(\b[16] ), .out0(new_n188));
  nano32aa1n02x4               g093(.a(new_n188), .b(new_n183), .c(new_n185), .d(new_n172), .out0(new_n189));
  aoi022aa1n02x5               g094(.a(new_n187), .b(new_n188), .c(new_n178), .d(new_n189), .o1(\s[17] ));
  inv000aa1d42x5               g095(.a(\a[17] ), .o1(new_n191));
  nanb02aa1d36x5               g096(.a(\b[16] ), .b(new_n191), .out0(new_n192));
  aoai13aa1n02x5               g097(.a(new_n188), .b(new_n186), .c(new_n121), .d(new_n177), .o1(new_n193));
  nor042aa1n03x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  nanp02aa1n04x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  norb02aa1n06x4               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  nano22aa1n02x4               g101(.a(new_n194), .b(new_n192), .c(new_n195), .out0(new_n197));
  nanp02aa1n02x5               g102(.a(new_n193), .b(new_n197), .o1(new_n198));
  aoai13aa1n02x5               g103(.a(new_n198), .b(new_n196), .c(new_n192), .d(new_n193), .o1(\s[18] ));
  and002aa1n02x5               g104(.a(new_n188), .b(new_n196), .o(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n186), .c(new_n121), .d(new_n177), .o1(new_n201));
  oaoi03aa1n12x5               g106(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  nor002aa1d32x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nand02aa1d16x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  norb02aa1n06x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n201), .c(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n08x5               g113(.a(new_n204), .o1(new_n209));
  aob012aa1n03x5               g114(.a(new_n206), .b(new_n201), .c(new_n203), .out0(new_n210));
  nor042aa1n06x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nand02aa1d08x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  norb02aa1n06x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  norb03aa1n02x5               g118(.a(new_n212), .b(new_n204), .c(new_n211), .out0(new_n214));
  nand42aa1n02x5               g119(.a(new_n210), .b(new_n214), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n213), .c(new_n209), .d(new_n210), .o1(\s[20] ));
  nano23aa1n06x5               g121(.a(new_n204), .b(new_n211), .c(new_n212), .d(new_n205), .out0(new_n217));
  nand23aa1n06x5               g122(.a(new_n217), .b(new_n188), .c(new_n196), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoi112aa1n09x5               g124(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n220));
  oai112aa1n06x5               g125(.a(new_n206), .b(new_n213), .c(new_n220), .d(new_n194), .o1(new_n221));
  oaoi03aa1n06x5               g126(.a(\a[20] ), .b(\b[19] ), .c(new_n209), .o1(new_n222));
  inv040aa1n02x5               g127(.a(new_n222), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(new_n221), .b(new_n223), .o1(new_n224));
  nor002aa1n16x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  nand42aa1n03x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  norb02aa1n15x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n187), .d(new_n219), .o1(new_n228));
  nona22aa1n02x4               g133(.a(new_n221), .b(new_n222), .c(new_n227), .out0(new_n229));
  aoi012aa1n02x5               g134(.a(new_n229), .b(new_n187), .c(new_n219), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n228), .b(new_n230), .out0(\s[21] ));
  inv000aa1d42x5               g136(.a(new_n225), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[21] ), .b(\a[22] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  oai022aa1n02x5               g139(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(\a[22] ), .c(\b[21] ), .o1(new_n236));
  nanp02aa1n03x5               g141(.a(new_n228), .b(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n234), .c(new_n232), .d(new_n228), .o1(\s[22] ));
  nanb02aa1n12x5               g143(.a(new_n233), .b(new_n227), .out0(new_n239));
  nano32aa1n02x4               g144(.a(new_n239), .b(new_n217), .c(new_n196), .d(new_n188), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n186), .c(new_n121), .d(new_n177), .o1(new_n241));
  aob012aa1n03x5               g146(.a(new_n235), .b(\b[21] ), .c(\a[22] ), .out0(new_n242));
  aoai13aa1n12x5               g147(.a(new_n242), .b(new_n239), .c(new_n221), .d(new_n223), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  aob012aa1n03x5               g150(.a(new_n245), .b(new_n241), .c(new_n244), .out0(new_n246));
  nano22aa1n03x7               g151(.a(new_n233), .b(new_n232), .c(new_n226), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n222), .c(new_n217), .d(new_n202), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n245), .o1(new_n249));
  and003aa1n02x5               g154(.a(new_n248), .b(new_n249), .c(new_n242), .o(new_n250));
  aobi12aa1n02x7               g155(.a(new_n246), .b(new_n250), .c(new_n241), .out0(\s[23] ));
  nor002aa1d24x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  inv030aa1n06x5               g157(.a(new_n252), .o1(new_n253));
  xorc02aa1n02x5               g158(.a(\a[24] ), .b(\b[23] ), .out0(new_n254));
  oai022aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n255));
  aoi012aa1n02x5               g160(.a(new_n255), .b(\a[24] ), .c(\b[23] ), .o1(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n249), .c(new_n241), .d(new_n244), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n254), .c(new_n246), .d(new_n253), .o1(\s[24] ));
  nand42aa1n03x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  tech160nm_fixnrc02aa1n05x5   g164(.a(\b[23] ), .b(\a[24] ), .out0(new_n260));
  nano22aa1n09x5               g165(.a(new_n260), .b(new_n253), .c(new_n259), .out0(new_n261));
  nano22aa1n02x4               g166(.a(new_n218), .b(new_n247), .c(new_n261), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n261), .o1(new_n263));
  oaoi03aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .c(new_n253), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n263), .c(new_n248), .d(new_n242), .o1(new_n266));
  tech160nm_fixorc02aa1n03p5x5 g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n266), .c(new_n187), .d(new_n262), .o1(new_n268));
  aoi112aa1n02x5               g173(.a(new_n267), .b(new_n264), .c(new_n243), .d(new_n261), .o1(new_n269));
  aobi12aa1n02x5               g174(.a(new_n269), .b(new_n187), .c(new_n262), .out0(new_n270));
  norb02aa1n02x5               g175(.a(new_n268), .b(new_n270), .out0(\s[25] ));
  norp02aa1n02x5               g176(.a(\b[24] ), .b(\a[25] ), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .out0(new_n274));
  nanp02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .o1(new_n275));
  oai022aa1n02x5               g180(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n276));
  norb02aa1n02x5               g181(.a(new_n275), .b(new_n276), .out0(new_n277));
  nand42aa1n02x5               g182(.a(new_n268), .b(new_n277), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n278), .b(new_n274), .c(new_n273), .d(new_n268), .o1(\s[26] ));
  and002aa1n02x5               g184(.a(new_n274), .b(new_n267), .o(new_n280));
  nano32aa1n03x7               g185(.a(new_n218), .b(new_n280), .c(new_n247), .d(new_n261), .out0(new_n281));
  aoai13aa1n12x5               g186(.a(new_n281), .b(new_n186), .c(new_n121), .d(new_n177), .o1(new_n282));
  aoai13aa1n09x5               g187(.a(new_n280), .b(new_n264), .c(new_n243), .d(new_n261), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n276), .b(new_n275), .o1(new_n284));
  nanp03aa1n06x5               g189(.a(new_n282), .b(new_n283), .c(new_n284), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  aoi122aa1n02x5               g191(.a(new_n286), .b(new_n275), .c(new_n276), .d(new_n266), .e(new_n280), .o1(new_n287));
  aoi022aa1n02x5               g192(.a(new_n287), .b(new_n282), .c(new_n285), .d(new_n286), .o1(\s[27] ));
  nor002aa1n12x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  nor002aa1n02x5               g194(.a(\b[27] ), .b(\a[28] ), .o1(new_n290));
  and002aa1n12x5               g195(.a(\b[27] ), .b(\a[28] ), .o(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n290), .o1(new_n292));
  inv000aa1n03x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n285), .d(new_n286), .o1(new_n294));
  aoi022aa1n03x5               g199(.a(new_n266), .b(new_n280), .c(new_n275), .d(new_n276), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n286), .o1(new_n296));
  norp03aa1n02x5               g201(.a(new_n291), .b(new_n290), .c(new_n289), .o1(new_n297));
  aoai13aa1n02x5               g202(.a(new_n297), .b(new_n296), .c(new_n295), .d(new_n282), .o1(new_n298));
  nanp02aa1n03x5               g203(.a(new_n294), .b(new_n298), .o1(\s[28] ));
  norb02aa1n03x5               g204(.a(new_n286), .b(new_n293), .out0(new_n300));
  nanp02aa1n03x5               g205(.a(new_n285), .b(new_n300), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n300), .o1(new_n302));
  aoib12aa1n06x5               g207(.a(new_n290), .b(new_n289), .c(new_n291), .out0(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n302), .c(new_n295), .d(new_n282), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n303), .b(new_n305), .out0(new_n306));
  aoi022aa1n03x5               g211(.a(new_n304), .b(new_n305), .c(new_n301), .d(new_n306), .o1(\s[29] ));
  xnrb03aa1n02x5               g212(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g213(.a(new_n305), .b(new_n286), .c(new_n292), .o1(new_n309));
  nanb02aa1n03x5               g214(.a(new_n309), .b(new_n285), .out0(new_n310));
  tech160nm_fioaoi03aa1n04x5   g215(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n311), .o1(new_n312));
  aoai13aa1n02x7               g217(.a(new_n312), .b(new_n309), .c(new_n295), .d(new_n282), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  aoi012aa1n02x5               g219(.a(new_n303), .b(\a[29] ), .c(\b[28] ), .o1(new_n315));
  oabi12aa1n02x5               g220(.a(new_n314), .b(\a[29] ), .c(\b[28] ), .out0(new_n316));
  norp02aa1n02x5               g221(.a(new_n315), .b(new_n316), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n313), .b(new_n314), .c(new_n310), .d(new_n317), .o1(\s[30] ));
  nanp03aa1n02x5               g223(.a(new_n300), .b(new_n305), .c(new_n314), .o1(new_n319));
  nanb02aa1n03x5               g224(.a(new_n319), .b(new_n285), .out0(new_n320));
  inv000aa1d42x5               g225(.a(\a[30] ), .o1(new_n321));
  inv000aa1d42x5               g226(.a(\b[29] ), .o1(new_n322));
  oaoi03aa1n02x5               g227(.a(new_n321), .b(new_n322), .c(new_n311), .o1(new_n323));
  aoai13aa1n02x7               g228(.a(new_n323), .b(new_n319), .c(new_n295), .d(new_n282), .o1(new_n324));
  xorc02aa1n02x5               g229(.a(\a[31] ), .b(\b[30] ), .out0(new_n325));
  oabi12aa1n02x5               g230(.a(new_n325), .b(\a[30] ), .c(\b[29] ), .out0(new_n326));
  oaoi13aa1n03x5               g231(.a(new_n326), .b(new_n311), .c(new_n321), .d(new_n322), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n324), .b(new_n325), .c(new_n320), .d(new_n327), .o1(\s[31] ));
  orn002aa1n02x5               g233(.a(\a[2] ), .b(\b[1] ), .o(new_n329));
  nanp02aa1n02x5               g234(.a(\b[1] ), .b(\a[2] ), .o1(new_n330));
  nanb03aa1n02x5               g235(.a(new_n100), .b(new_n329), .c(new_n330), .out0(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n102), .b(new_n331), .c(new_n329), .out0(\s[3] ));
  nanp02aa1n02x5               g237(.a(new_n101), .b(new_n102), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[4] ), .b(\b[3] ), .out0(new_n334));
  oab012aa1n02x4               g239(.a(new_n334), .b(\a[3] ), .c(\b[2] ), .out0(new_n335));
  aboi22aa1n03x5               g240(.a(new_n104), .b(new_n334), .c(new_n335), .d(new_n333), .out0(\s[4] ));
  and002aa1n02x5               g241(.a(\b[4] ), .b(\a[5] ), .o(new_n337));
  orn003aa1d24x5               g242(.a(new_n104), .b(new_n337), .c(new_n110), .o(new_n338));
  obai22aa1n02x7               g243(.a(new_n109), .b(new_n104), .c(new_n114), .d(new_n337), .out0(new_n339));
  and002aa1n02x5               g244(.a(new_n338), .b(new_n339), .o(\s[5] ));
  and002aa1n02x5               g245(.a(\b[5] ), .b(\a[6] ), .o(new_n341));
  norp02aa1n02x5               g246(.a(\b[5] ), .b(\a[6] ), .o1(new_n342));
  norp02aa1n02x5               g247(.a(new_n341), .b(new_n342), .o1(new_n343));
  nona32aa1n03x5               g248(.a(new_n338), .b(new_n342), .c(new_n341), .d(new_n114), .out0(new_n344));
  aoai13aa1n02x5               g249(.a(new_n344), .b(new_n343), .c(new_n115), .d(new_n338), .o1(\s[6] ));
  norb02aa1n02x5               g250(.a(new_n107), .b(new_n105), .out0(new_n346));
  aoib12aa1n02x5               g251(.a(new_n346), .b(new_n344), .c(new_n341), .out0(new_n347));
  aoi022aa1n02x5               g252(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n348));
  nano22aa1n03x7               g253(.a(new_n105), .b(new_n344), .c(new_n348), .out0(new_n349));
  norp02aa1n02x5               g254(.a(new_n349), .b(new_n347), .o1(\s[7] ));
  obai22aa1n03x5               g255(.a(new_n106), .b(new_n117), .c(new_n349), .d(new_n105), .out0(new_n351));
  norb03aa1n02x5               g256(.a(new_n106), .b(new_n105), .c(new_n117), .out0(new_n352));
  oaib12aa1n03x5               g257(.a(new_n351), .b(new_n349), .c(new_n352), .out0(\s[8] ));
  nanp02aa1n02x5               g258(.a(new_n118), .b(new_n116), .o1(new_n354));
  and002aa1n02x5               g259(.a(new_n141), .b(new_n119), .o(new_n355));
  oai112aa1n02x5               g260(.a(new_n354), .b(new_n355), .c(new_n104), .d(new_n113), .o1(new_n356));
  oaib12aa1n02x5               g261(.a(new_n356), .b(new_n141), .c(new_n121), .out0(\s[9] ));
endmodule


