// Benchmark "adder" written by ABC on Wed Jul 17 14:06:38 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n332, new_n333, new_n335, new_n336, new_n338, new_n339, new_n340,
    new_n341, new_n343, new_n344, new_n347, new_n348, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n20x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1n20x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nand42aa1n03x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  orn002aa1n02x5               g006(.a(\a[2] ), .b(\b[1] ), .o(new_n102));
  nanp02aa1n04x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  aob012aa1n12x5               g008(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(new_n104));
  inv040aa1d32x5               g009(.a(\a[3] ), .o1(new_n105));
  inv000aa1d42x5               g010(.a(\b[2] ), .o1(new_n106));
  nand22aa1n03x5               g011(.a(new_n106), .b(new_n105), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand42aa1n02x5               g013(.a(new_n107), .b(new_n108), .o1(new_n109));
  oa0022aa1n02x5               g014(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n110));
  aoai13aa1n04x5               g015(.a(new_n110), .b(new_n109), .c(new_n104), .d(new_n102), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  norp02aa1n04x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  tech160nm_fiaoi012aa1n03p5x5 g018(.a(new_n113), .b(\a[6] ), .c(\b[5] ), .o1(new_n114));
  norp02aa1n04x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  aoi012aa1n02x7               g020(.a(new_n115), .b(\a[4] ), .c(\b[3] ), .o1(new_n116));
  nand42aa1n06x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor002aa1d32x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand42aa1d28x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  norp02aa1n02x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n119), .b(new_n117), .c(new_n120), .d(new_n118), .out0(new_n121));
  nano32aa1n02x4               g026(.a(new_n121), .b(new_n116), .c(new_n114), .d(new_n112), .out0(new_n122));
  tech160nm_finand02aa1n05x5   g027(.a(new_n122), .b(new_n111), .o1(new_n123));
  nand42aa1n08x5               g028(.a(\b[5] ), .b(\a[6] ), .o1(new_n124));
  nano22aa1n02x5               g029(.a(new_n118), .b(new_n124), .c(new_n119), .out0(new_n125));
  oai022aa1n02x5               g030(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n126));
  norb02aa1n03x5               g031(.a(new_n117), .b(new_n115), .out0(new_n127));
  inv000aa1d42x5               g032(.a(new_n118), .o1(new_n128));
  oaoi03aa1n02x5               g033(.a(\a[8] ), .b(\b[7] ), .c(new_n128), .o1(new_n129));
  aoi013aa1n06x5               g034(.a(new_n129), .b(new_n125), .c(new_n127), .d(new_n126), .o1(new_n130));
  nanp02aa1n06x5               g035(.a(new_n123), .b(new_n130), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(new_n131), .b(new_n101), .o1(new_n132));
  obai22aa1n02x7               g037(.a(new_n132), .b(new_n100), .c(new_n97), .d(new_n99), .out0(new_n133));
  nona32aa1n02x4               g038(.a(new_n132), .b(new_n100), .c(new_n99), .d(new_n97), .out0(new_n134));
  nanp02aa1n02x5               g039(.a(new_n133), .b(new_n134), .o1(\s[10] ));
  nand42aa1n06x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n137), .b(\a[10] ), .c(\b[9] ), .o1(new_n138));
  inv000aa1n06x5               g043(.a(new_n137), .o1(new_n139));
  aoi022aa1n02x5               g044(.a(new_n134), .b(new_n98), .c(new_n139), .d(new_n136), .o1(new_n140));
  aoi013aa1n02x4               g045(.a(new_n140), .b(new_n138), .c(new_n136), .d(new_n134), .o1(\s[11] ));
  nanp03aa1n02x5               g046(.a(new_n134), .b(new_n136), .c(new_n138), .o1(new_n142));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1d28x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n03x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  norp02aa1n02x5               g050(.a(new_n145), .b(new_n137), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(new_n142), .b(new_n139), .o1(new_n147));
  aoi022aa1n02x5               g052(.a(new_n147), .b(new_n145), .c(new_n142), .d(new_n146), .o1(\s[12] ));
  nona23aa1n02x5               g053(.a(new_n101), .b(new_n98), .c(new_n97), .d(new_n100), .out0(new_n149));
  nano32aa1n06x5               g054(.a(new_n149), .b(new_n145), .c(new_n139), .d(new_n136), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n131), .b(new_n150), .o1(new_n151));
  nanb03aa1n06x5               g056(.a(new_n143), .b(new_n144), .c(new_n136), .out0(new_n152));
  oai112aa1n06x5               g057(.a(new_n139), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n153));
  aoi012aa1n12x5               g058(.a(new_n143), .b(new_n137), .c(new_n144), .o1(new_n154));
  oai012aa1n18x5               g059(.a(new_n154), .b(new_n153), .c(new_n152), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n155), .b(new_n151), .out0(new_n156));
  nor002aa1d32x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nand02aa1n04x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n157), .b(new_n158), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  oai112aa1n02x5               g065(.a(new_n154), .b(new_n159), .c(new_n153), .d(new_n152), .o1(new_n161));
  aboi22aa1n03x5               g066(.a(new_n161), .b(new_n151), .c(new_n156), .d(new_n160), .out0(\s[13] ));
  inv000aa1d42x5               g067(.a(new_n157), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n160), .b(new_n155), .c(new_n131), .d(new_n150), .o1(new_n164));
  nor002aa1n16x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand22aa1n12x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  xobna2aa1n03x5               g072(.a(new_n167), .b(new_n164), .c(new_n163), .out0(\s[14] ));
  nona23aa1d18x5               g073(.a(new_n166), .b(new_n158), .c(new_n157), .d(new_n165), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n155), .c(new_n131), .d(new_n150), .o1(new_n171));
  aoi012aa1n06x5               g076(.a(new_n165), .b(new_n157), .c(new_n166), .o1(new_n172));
  nor002aa1d32x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n171), .c(new_n172), .out0(\s[15] ));
  aob012aa1n03x5               g081(.a(new_n175), .b(new_n171), .c(new_n172), .out0(new_n177));
  nor002aa1d32x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanp02aa1n09x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  aoib12aa1n02x5               g085(.a(new_n173), .b(new_n179), .c(new_n178), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n173), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n175), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n171), .d(new_n172), .o1(new_n184));
  aoi022aa1n03x5               g089(.a(new_n184), .b(new_n180), .c(new_n177), .d(new_n181), .o1(\s[16] ));
  nona23aa1d18x5               g090(.a(new_n179), .b(new_n174), .c(new_n173), .d(new_n178), .out0(new_n186));
  nor042aa1d18x5               g091(.a(new_n186), .b(new_n169), .o1(new_n187));
  nand22aa1n12x5               g092(.a(new_n150), .b(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  tech160nm_fiaoi012aa1n03p5x5 g094(.a(new_n178), .b(new_n173), .c(new_n179), .o1(new_n190));
  tech160nm_fioai012aa1n05x5   g095(.a(new_n190), .b(new_n186), .c(new_n172), .o1(new_n191));
  aoi012aa1d24x5               g096(.a(new_n191), .b(new_n155), .c(new_n187), .o1(new_n192));
  aoai13aa1n12x5               g097(.a(new_n192), .b(new_n188), .c(new_n123), .d(new_n130), .o1(new_n193));
  nor042aa1d18x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  nanp02aa1n03x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  oaib12aa1n02x5               g100(.a(new_n193), .b(new_n194), .c(new_n195), .out0(new_n196));
  oai022aa1n02x5               g101(.a(\a[16] ), .b(\b[15] ), .c(\b[16] ), .d(\a[17] ), .o1(new_n197));
  aoi122aa1n02x5               g102(.a(new_n197), .b(\b[16] ), .c(\a[17] ), .d(new_n173), .e(new_n179), .o1(new_n198));
  oai012aa1n02x5               g103(.a(new_n198), .b(new_n186), .c(new_n172), .o1(new_n199));
  tech160nm_fiao0012aa1n02p5x5 g104(.a(new_n199), .b(new_n155), .c(new_n187), .o(new_n200));
  aoai13aa1n02x5               g105(.a(new_n196), .b(new_n200), .c(new_n189), .d(new_n131), .o1(\s[17] ));
  inv040aa1n08x5               g106(.a(new_n194), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(new_n193), .b(new_n195), .o1(new_n203));
  xorc02aa1n12x5               g108(.a(\a[18] ), .b(\b[17] ), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n203), .c(new_n202), .out0(\s[18] ));
  and003aa1n12x5               g110(.a(new_n204), .b(new_n195), .c(new_n202), .o(new_n206));
  oaoi03aa1n12x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n207));
  xorc02aa1n12x5               g112(.a(\a[19] ), .b(\b[18] ), .out0(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n207), .c(new_n193), .d(new_n206), .o1(new_n209));
  aoi112aa1n02x5               g114(.a(new_n208), .b(new_n207), .c(new_n193), .d(new_n206), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n209), .b(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  xorc02aa1n12x5               g117(.a(\a[20] ), .b(\b[19] ), .out0(new_n213));
  norp02aa1n02x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norp02aa1n02x5               g119(.a(new_n213), .b(new_n214), .o1(new_n215));
  inv000aa1d42x5               g120(.a(\a[19] ), .o1(new_n216));
  oaib12aa1n06x5               g121(.a(new_n209), .b(\b[18] ), .c(new_n216), .out0(new_n217));
  aoi022aa1n02x5               g122(.a(new_n217), .b(new_n213), .c(new_n209), .d(new_n215), .o1(\s[20] ));
  inv000aa1d42x5               g123(.a(\a[20] ), .o1(new_n219));
  xroi22aa1d04x5               g124(.a(new_n216), .b(\b[18] ), .c(new_n219), .d(\b[19] ), .out0(new_n220));
  nand22aa1n03x5               g125(.a(new_n206), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  nanp03aa1d12x5               g127(.a(new_n207), .b(new_n208), .c(new_n213), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[19] ), .o1(new_n224));
  oaoi03aa1n03x5               g129(.a(new_n219), .b(new_n224), .c(new_n214), .o1(new_n225));
  nanp02aa1n02x5               g130(.a(new_n223), .b(new_n225), .o1(new_n226));
  xorc02aa1n02x5               g131(.a(\a[21] ), .b(\b[20] ), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n226), .c(new_n193), .d(new_n222), .o1(new_n228));
  nano22aa1n02x4               g133(.a(new_n227), .b(new_n223), .c(new_n225), .out0(new_n229));
  aobi12aa1n02x5               g134(.a(new_n229), .b(new_n193), .c(new_n222), .out0(new_n230));
  norb02aa1n02x5               g135(.a(new_n228), .b(new_n230), .out0(\s[21] ));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  inv040aa1d30x5               g137(.a(\a[21] ), .o1(new_n233));
  aoib12aa1n02x5               g138(.a(new_n232), .b(new_n233), .c(\b[20] ), .out0(new_n234));
  oaib12aa1n06x5               g139(.a(new_n228), .b(\b[20] ), .c(new_n233), .out0(new_n235));
  aoi022aa1n02x5               g140(.a(new_n235), .b(new_n232), .c(new_n228), .d(new_n234), .o1(\s[22] ));
  inv040aa1d32x5               g141(.a(\a[22] ), .o1(new_n237));
  xroi22aa1d06x4               g142(.a(new_n233), .b(\b[20] ), .c(new_n237), .d(\b[21] ), .out0(new_n238));
  and003aa1n02x5               g143(.a(new_n206), .b(new_n238), .c(new_n220), .o(new_n239));
  inv020aa1n03x5               g144(.a(new_n238), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(\b[20] ), .b(\a[21] ), .c(\a[22] ), .d(\b[21] ), .o1(new_n241));
  aoib12aa1n02x5               g146(.a(new_n241), .b(new_n237), .c(\b[21] ), .out0(new_n242));
  aoai13aa1n09x5               g147(.a(new_n242), .b(new_n240), .c(new_n223), .d(new_n225), .o1(new_n243));
  tech160nm_fixorc02aa1n03p5x5 g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n243), .c(new_n193), .d(new_n239), .o1(new_n245));
  nanb02aa1n02x5               g150(.a(new_n244), .b(new_n242), .out0(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(new_n226), .c(new_n238), .o1(new_n247));
  aobi12aa1n02x5               g152(.a(new_n247), .b(new_n193), .c(new_n239), .out0(new_n248));
  norb02aa1n02x5               g153(.a(new_n245), .b(new_n248), .out0(\s[23] ));
  tech160nm_fixorc02aa1n03p5x5 g154(.a(\a[24] ), .b(\b[23] ), .out0(new_n250));
  norp02aa1n02x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  norp02aa1n02x5               g156(.a(new_n250), .b(new_n251), .o1(new_n252));
  oai012aa1n06x5               g157(.a(new_n245), .b(\b[22] ), .c(\a[23] ), .o1(new_n253));
  aoi022aa1n02x7               g158(.a(new_n253), .b(new_n250), .c(new_n245), .d(new_n252), .o1(\s[24] ));
  and002aa1n06x5               g159(.a(new_n250), .b(new_n244), .o(new_n255));
  nona23aa1n06x5               g160(.a(new_n193), .b(new_n255), .c(new_n240), .d(new_n221), .out0(new_n256));
  inv000aa1d42x5               g161(.a(\a[24] ), .o1(new_n257));
  inv000aa1d42x5               g162(.a(\b[23] ), .o1(new_n258));
  tech160nm_fioaoi03aa1n02p5x5 g163(.a(new_n257), .b(new_n258), .c(new_n251), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  aoi012aa1d18x5               g165(.a(new_n260), .b(new_n243), .c(new_n255), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n192), .o1(new_n263));
  aoi012aa1n02x5               g168(.a(new_n263), .b(new_n131), .c(new_n189), .o1(new_n264));
  nano32aa1n03x7               g169(.a(new_n264), .b(new_n255), .c(new_n222), .d(new_n238), .out0(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  oai012aa1n02x5               g171(.a(new_n266), .b(new_n265), .c(new_n262), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n266), .b(new_n260), .c(new_n243), .d(new_n255), .o1(new_n268));
  aobi12aa1n03x7               g173(.a(new_n267), .b(new_n268), .c(new_n256), .out0(\s[25] ));
  xorc02aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .out0(new_n270));
  nor042aa1n06x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  norp02aa1n02x5               g176(.a(new_n270), .b(new_n271), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n266), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n273), .b(new_n274), .c(new_n256), .d(new_n261), .o1(new_n275));
  aoi022aa1n03x5               g180(.a(new_n275), .b(new_n270), .c(new_n267), .d(new_n272), .o1(\s[26] ));
  and002aa1n02x5               g181(.a(new_n270), .b(new_n266), .o(new_n277));
  aoai13aa1n04x5               g182(.a(new_n277), .b(new_n260), .c(new_n243), .d(new_n255), .o1(new_n278));
  nano32aa1n03x7               g183(.a(new_n221), .b(new_n277), .c(new_n238), .d(new_n255), .out0(new_n279));
  norp02aa1n02x5               g184(.a(\b[25] ), .b(\a[26] ), .o1(new_n280));
  aob012aa1n02x5               g185(.a(new_n271), .b(\b[25] ), .c(\a[26] ), .out0(new_n281));
  norb02aa1n02x5               g186(.a(new_n281), .b(new_n280), .out0(new_n282));
  inv000aa1n02x5               g187(.a(new_n282), .o1(new_n283));
  tech160nm_fiaoi012aa1n05x5   g188(.a(new_n283), .b(new_n193), .c(new_n279), .o1(new_n284));
  nor042aa1n03x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  and002aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o(new_n286));
  norp02aa1n02x5               g191(.a(new_n286), .b(new_n285), .o1(new_n287));
  nanp02aa1n06x5               g192(.a(new_n193), .b(new_n279), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n285), .o1(new_n289));
  nano23aa1n02x4               g194(.a(new_n286), .b(new_n280), .c(new_n281), .d(new_n289), .out0(new_n290));
  nanp03aa1n02x5               g195(.a(new_n278), .b(new_n288), .c(new_n290), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n291), .b(new_n287), .c(new_n284), .d(new_n278), .o1(\s[27] ));
  inv000aa1d42x5               g197(.a(\b[26] ), .o1(new_n293));
  nand23aa1n03x5               g198(.a(new_n278), .b(new_n288), .c(new_n282), .o1(new_n294));
  oaib12aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(\a[27] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n289), .b(new_n286), .c(new_n284), .d(new_n278), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .out0(new_n297));
  norp02aa1n02x5               g202(.a(new_n297), .b(new_n285), .o1(new_n298));
  aoi022aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n295), .d(new_n298), .o1(\s[28] ));
  inv000aa1d42x5               g204(.a(\a[28] ), .o1(new_n300));
  xroi22aa1d04x5               g205(.a(\a[27] ), .b(new_n293), .c(new_n300), .d(\b[27] ), .out0(new_n301));
  nand42aa1n02x5               g206(.a(new_n294), .b(new_n301), .o1(new_n302));
  inv000aa1n03x5               g207(.a(new_n301), .o1(new_n303));
  oaoi03aa1n12x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n303), .c(new_n284), .d(new_n278), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norp02aa1n02x5               g212(.a(new_n304), .b(new_n307), .o1(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n302), .d(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g215(.a(new_n297), .b(new_n307), .c(new_n287), .o(new_n311));
  nanp02aa1n03x5               g216(.a(new_n294), .b(new_n311), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  inv000aa1d42x5               g218(.a(\b[28] ), .o1(new_n314));
  oaib12aa1n02x5               g219(.a(new_n304), .b(new_n314), .c(\a[29] ), .out0(new_n315));
  oa0012aa1n02x5               g220(.a(new_n315), .b(\b[28] ), .c(\a[29] ), .o(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n313), .c(new_n284), .d(new_n278), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .out0(new_n318));
  oabi12aa1n02x5               g223(.a(new_n318), .b(\a[29] ), .c(\b[28] ), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n315), .b(new_n319), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n317), .b(new_n318), .c(new_n312), .d(new_n320), .o1(\s[30] ));
  nano22aa1n02x4               g226(.a(new_n303), .b(new_n307), .c(new_n318), .out0(new_n322));
  nand42aa1n02x5               g227(.a(new_n294), .b(new_n322), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[31] ), .b(\b[30] ), .out0(new_n324));
  oai122aa1n02x7               g229(.a(new_n315), .b(\a[30] ), .c(\b[29] ), .d(\a[29] ), .e(\b[28] ), .o1(new_n325));
  aob012aa1n02x5               g230(.a(new_n325), .b(\b[29] ), .c(\a[30] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n326), .b(new_n324), .out0(new_n327));
  inv000aa1n02x5               g232(.a(new_n322), .o1(new_n328));
  aoai13aa1n03x5               g233(.a(new_n326), .b(new_n328), .c(new_n284), .d(new_n278), .o1(new_n329));
  aoi022aa1n03x5               g234(.a(new_n329), .b(new_n324), .c(new_n323), .d(new_n327), .o1(\s[31] ));
  xobna2aa1n03x5               g235(.a(new_n109), .b(new_n104), .c(new_n102), .out0(\s[3] ));
  tech160nm_fiao0012aa1n02p5x5 g236(.a(new_n109), .b(new_n102), .c(new_n104), .o(new_n332));
  xorc02aa1n02x5               g237(.a(\a[4] ), .b(\b[3] ), .out0(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n332), .c(new_n107), .out0(\s[4] ));
  nanp02aa1n02x5               g239(.a(\b[3] ), .b(\a[4] ), .o1(new_n335));
  nanb02aa1n02x5               g240(.a(new_n113), .b(new_n112), .out0(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n336), .b(new_n111), .c(new_n335), .out0(\s[5] ));
  norb02aa1n02x5               g242(.a(new_n124), .b(new_n120), .out0(new_n338));
  aoi013aa1n02x4               g243(.a(new_n113), .b(new_n111), .c(new_n112), .d(new_n335), .o1(new_n339));
  nanp03aa1n02x5               g244(.a(new_n111), .b(new_n112), .c(new_n335), .o1(new_n340));
  oai112aa1n02x5               g245(.a(new_n340), .b(new_n338), .c(\b[4] ), .d(\a[5] ), .o1(new_n341));
  oai012aa1n02x5               g246(.a(new_n341), .b(new_n339), .c(new_n338), .o1(\s[6] ));
  nanp02aa1n02x5               g247(.a(new_n341), .b(new_n125), .o1(new_n343));
  aoi022aa1n02x5               g248(.a(new_n341), .b(new_n124), .c(new_n128), .d(new_n119), .o1(new_n344));
  norb02aa1n02x5               g249(.a(new_n343), .b(new_n344), .out0(\s[7] ));
  xnbna2aa1n03x5               g250(.a(new_n127), .b(new_n343), .c(new_n128), .out0(\s[8] ));
  nanb02aa1n02x5               g251(.a(new_n100), .b(new_n101), .out0(new_n347));
  inv000aa1d42x5               g252(.a(new_n347), .o1(new_n348));
  aoi113aa1n02x5               g253(.a(new_n129), .b(new_n348), .c(new_n125), .d(new_n127), .e(new_n126), .o1(new_n349));
  aoi022aa1n02x5               g254(.a(new_n131), .b(new_n348), .c(new_n349), .d(new_n123), .o1(\s[9] ));
endmodule


