// Benchmark "adder" written by ABC on Thu Jul 18 12:31:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n155, new_n156, new_n157, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n342, new_n343, new_n344,
    new_n346, new_n349, new_n350, new_n351, new_n353, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[1] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\b[0] ), .o1(new_n98));
  nor022aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oaoi13aa1n04x5               g005(.a(new_n99), .b(new_n100), .c(new_n97), .d(new_n98), .o1(new_n101));
  nor022aa1n16x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n106));
  tech160nm_fioai012aa1n05x5   g011(.a(new_n103), .b(new_n104), .c(new_n102), .o1(new_n107));
  oai012aa1n06x5               g012(.a(new_n107), .b(new_n106), .c(new_n101), .o1(new_n108));
  nor022aa1n08x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor002aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nona23aa1n02x4               g017(.a(new_n111), .b(new_n110), .c(new_n112), .d(new_n109), .out0(new_n113));
  nor002aa1n16x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  norb02aa1n03x5               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  nor042aa1n06x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand42aa1n08x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  norb02aa1n03x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  nano22aa1n03x7               g024(.a(new_n113), .b(new_n116), .c(new_n119), .out0(new_n120));
  aoi022aa1d24x5               g025(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n121));
  oaoi13aa1n02x7               g026(.a(new_n109), .b(new_n121), .c(new_n117), .d(new_n114), .o1(new_n122));
  oaoi03aa1n03x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  nor042aa1n02x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nand42aa1n10x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n127));
  oai012aa1n02x5               g032(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nor002aa1n12x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nand42aa1n10x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor002aa1n02x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nona22aa1n02x4               g039(.a(new_n127), .b(new_n124), .c(new_n134), .out0(new_n135));
  aoi022aa1n02x5               g040(.a(new_n135), .b(new_n130), .c(new_n132), .d(new_n133), .o1(new_n136));
  and002aa1n06x5               g041(.a(\b[0] ), .b(\a[1] ), .o(new_n137));
  oaoi03aa1n03x5               g042(.a(\a[2] ), .b(\b[1] ), .c(new_n137), .o1(new_n138));
  norb02aa1n06x5               g043(.a(new_n103), .b(new_n102), .out0(new_n139));
  norb02aa1n02x7               g044(.a(new_n105), .b(new_n104), .out0(new_n140));
  nand03aa1n02x5               g045(.a(new_n138), .b(new_n139), .c(new_n140), .o1(new_n141));
  nano23aa1n03x7               g046(.a(new_n112), .b(new_n109), .c(new_n110), .d(new_n111), .out0(new_n142));
  nanp03aa1n02x5               g047(.a(new_n142), .b(new_n116), .c(new_n119), .o1(new_n143));
  inv000aa1d42x5               g048(.a(\a[7] ), .o1(new_n144));
  inv000aa1d42x5               g049(.a(\b[6] ), .o1(new_n145));
  nanp02aa1n02x5               g050(.a(new_n145), .b(new_n144), .o1(new_n146));
  oai012aa1n06x5               g051(.a(new_n121), .b(new_n117), .c(new_n114), .o1(new_n147));
  nanp02aa1n03x5               g052(.a(new_n147), .b(new_n146), .o1(new_n148));
  tech160nm_fiaoi012aa1n02p5x5 g053(.a(new_n112), .b(new_n148), .c(new_n111), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n143), .c(new_n141), .d(new_n107), .o1(new_n150));
  oai022aa1n04x7               g055(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n151));
  nano22aa1n02x4               g056(.a(new_n131), .b(new_n130), .c(new_n133), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n151), .c(new_n150), .d(new_n126), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n153), .b(new_n136), .out0(\s[11] ));
  nor042aa1n02x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand42aa1n16x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  norb02aa1n06x4               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n153), .c(new_n132), .out0(\s[12] ));
  nanp02aa1n03x5               g063(.a(new_n108), .b(new_n120), .o1(new_n159));
  nano23aa1n03x5               g064(.a(new_n134), .b(new_n155), .c(new_n156), .d(new_n130), .out0(new_n160));
  nano23aa1n03x5               g065(.a(new_n124), .b(new_n131), .c(new_n133), .d(new_n125), .out0(new_n161));
  nand22aa1n03x5               g066(.a(new_n161), .b(new_n160), .o1(new_n162));
  nanp03aa1n02x5               g067(.a(new_n151), .b(new_n130), .c(new_n133), .o1(new_n163));
  nand23aa1n03x5               g068(.a(new_n163), .b(new_n132), .c(new_n157), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(new_n164), .b(new_n156), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n162), .c(new_n159), .d(new_n149), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  nand42aa1d28x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  nor002aa1d32x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1d28x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nanb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n174));
  nona22aa1n02x4               g079(.a(new_n172), .b(new_n171), .c(new_n168), .out0(new_n175));
  aoai13aa1n02x5               g080(.a(new_n174), .b(new_n175), .c(new_n170), .d(new_n166), .o1(\s[14] ));
  nano23aa1n06x5               g081(.a(new_n168), .b(new_n171), .c(new_n172), .d(new_n169), .out0(new_n177));
  inv000aa1d42x5               g082(.a(new_n168), .o1(new_n178));
  oaoi03aa1n02x5               g083(.a(\a[14] ), .b(\b[13] ), .c(new_n178), .o1(new_n179));
  tech160nm_fixorc02aa1n05x5   g084(.a(\a[15] ), .b(\b[14] ), .out0(new_n180));
  aoai13aa1n06x5               g085(.a(new_n180), .b(new_n179), .c(new_n166), .d(new_n177), .o1(new_n181));
  aoi112aa1n02x5               g086(.a(new_n180), .b(new_n179), .c(new_n166), .d(new_n177), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n181), .b(new_n182), .out0(\s[15] ));
  inv000aa1d42x5               g088(.a(\a[15] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\b[14] ), .o1(new_n185));
  nanp02aa1n02x5               g090(.a(new_n185), .b(new_n184), .o1(new_n186));
  nor002aa1n10x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  and002aa1n12x5               g092(.a(\b[15] ), .b(\a[16] ), .o(new_n188));
  nor042aa1n02x5               g093(.a(new_n188), .b(new_n187), .o1(new_n189));
  oai022aa1n02x5               g094(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n190));
  nona22aa1n03x5               g095(.a(new_n181), .b(new_n188), .c(new_n190), .out0(new_n191));
  aoai13aa1n03x5               g096(.a(new_n191), .b(new_n189), .c(new_n186), .d(new_n181), .o1(\s[16] ));
  nano32aa1n03x7               g097(.a(new_n162), .b(new_n189), .c(new_n177), .d(new_n180), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n194));
  aoi112aa1n03x5               g099(.a(new_n188), .b(new_n187), .c(\a[15] ), .d(\b[14] ), .o1(new_n195));
  oai012aa1n02x5               g100(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .o1(new_n196));
  nano23aa1n03x7               g101(.a(new_n173), .b(new_n196), .c(new_n178), .d(new_n156), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n187), .o1(new_n198));
  oai122aa1n06x5               g103(.a(new_n172), .b(new_n171), .c(new_n168), .d(new_n185), .e(new_n184), .o1(new_n199));
  aoai13aa1n03x5               g104(.a(new_n198), .b(new_n188), .c(new_n199), .d(new_n186), .o1(new_n200));
  aoi013aa1n06x5               g105(.a(new_n200), .b(new_n164), .c(new_n197), .d(new_n195), .o1(new_n201));
  xnrc02aa1n12x5               g106(.a(\b[16] ), .b(\a[17] ), .out0(new_n202));
  xobna2aa1n03x5               g107(.a(new_n202), .b(new_n194), .c(new_n201), .out0(\s[17] ));
  nor002aa1n03x5               g108(.a(\b[16] ), .b(\a[17] ), .o1(new_n204));
  inv040aa1n03x5               g109(.a(new_n204), .o1(new_n205));
  nanp02aa1n12x5               g110(.a(new_n194), .b(new_n201), .o1(new_n206));
  nanb02aa1n06x5               g111(.a(new_n202), .b(new_n206), .out0(new_n207));
  nor042aa1n06x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand22aa1n12x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  norb02aa1n06x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  oai022aa1n04x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  nanb03aa1n03x5               g116(.a(new_n211), .b(new_n207), .c(new_n209), .out0(new_n212));
  aoai13aa1n02x5               g117(.a(new_n212), .b(new_n210), .c(new_n205), .d(new_n207), .o1(\s[18] ));
  norb02aa1d21x5               g118(.a(new_n210), .b(new_n202), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  oaoi03aa1n02x5               g120(.a(\a[18] ), .b(\b[17] ), .c(new_n205), .o1(new_n216));
  inv000aa1n02x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n03x5               g122(.a(new_n217), .b(new_n215), .c(new_n194), .d(new_n201), .o1(new_n218));
  xorc02aa1n02x5               g123(.a(\a[19] ), .b(\b[18] ), .out0(new_n219));
  aoi112aa1n02x5               g124(.a(new_n219), .b(new_n216), .c(new_n206), .d(new_n214), .o1(new_n220));
  aoi012aa1n02x5               g125(.a(new_n220), .b(new_n218), .c(new_n219), .o1(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nand42aa1n06x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  inv040aa1d32x5               g130(.a(\a[19] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[18] ), .o1(new_n227));
  oaoi03aa1n02x5               g132(.a(new_n226), .b(new_n227), .c(new_n218), .o1(new_n228));
  nand02aa1n02x5               g133(.a(new_n218), .b(new_n219), .o1(new_n229));
  aoi012aa1n02x5               g134(.a(new_n223), .b(new_n226), .c(new_n227), .o1(new_n230));
  nanp03aa1n02x5               g135(.a(new_n229), .b(new_n224), .c(new_n230), .o1(new_n231));
  oaih12aa1n02x5               g136(.a(new_n231), .b(new_n228), .c(new_n225), .o1(\s[20] ));
  nand42aa1n03x5               g137(.a(new_n227), .b(new_n226), .o1(new_n233));
  nand42aa1n04x5               g138(.a(\b[18] ), .b(\a[19] ), .o1(new_n234));
  nano32aa1n03x7               g139(.a(new_n223), .b(new_n233), .c(new_n224), .d(new_n234), .out0(new_n235));
  nand22aa1n12x5               g140(.a(new_n214), .b(new_n235), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nanb03aa1n02x5               g142(.a(new_n223), .b(new_n224), .c(new_n234), .out0(new_n238));
  nand03aa1n02x5               g143(.a(new_n211), .b(new_n233), .c(new_n209), .o1(new_n239));
  aoai13aa1n04x5               g144(.a(new_n224), .b(new_n223), .c(new_n226), .d(new_n227), .o1(new_n240));
  oai012aa1n06x5               g145(.a(new_n240), .b(new_n239), .c(new_n238), .o1(new_n241));
  nor002aa1d32x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  nanp02aa1n06x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n243), .b(new_n242), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n241), .c(new_n206), .d(new_n237), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n244), .b(new_n241), .c(new_n206), .d(new_n237), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n245), .b(new_n246), .out0(\s[21] ));
  inv000aa1d42x5               g152(.a(new_n242), .o1(new_n248));
  nor042aa1n02x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  nand02aa1d06x5               g154(.a(\b[21] ), .b(\a[22] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n250), .b(new_n249), .out0(new_n251));
  norb03aa1n02x5               g156(.a(new_n250), .b(new_n242), .c(new_n249), .out0(new_n252));
  nand42aa1n02x5               g157(.a(new_n245), .b(new_n252), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n251), .c(new_n248), .d(new_n245), .o1(\s[22] ));
  nano23aa1n06x5               g159(.a(new_n242), .b(new_n249), .c(new_n250), .d(new_n243), .out0(new_n255));
  nano22aa1n02x4               g160(.a(new_n215), .b(new_n235), .c(new_n255), .out0(new_n256));
  nano22aa1n03x5               g161(.a(new_n223), .b(new_n234), .c(new_n224), .out0(new_n257));
  oai012aa1n02x5               g162(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .o1(new_n258));
  oab012aa1n02x5               g163(.a(new_n258), .b(new_n204), .c(new_n208), .out0(new_n259));
  inv000aa1n02x5               g164(.a(new_n240), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n255), .b(new_n260), .c(new_n259), .d(new_n257), .o1(new_n261));
  oaoi03aa1n09x5               g166(.a(\a[22] ), .b(\b[21] ), .c(new_n248), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(new_n261), .b(new_n263), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[23] ), .b(\b[22] ), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n264), .c(new_n206), .d(new_n256), .o1(new_n266));
  aoi112aa1n02x5               g171(.a(new_n265), .b(new_n264), .c(new_n206), .d(new_n256), .o1(new_n267));
  norb02aa1n03x4               g172(.a(new_n266), .b(new_n267), .out0(\s[23] ));
  norp02aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[24] ), .b(\b[23] ), .out0(new_n271));
  nanp02aa1n02x5               g176(.a(\b[23] ), .b(\a[24] ), .o1(new_n272));
  oai022aa1n02x5               g177(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n273));
  norb02aa1n02x5               g178(.a(new_n272), .b(new_n273), .out0(new_n274));
  nanp02aa1n03x5               g179(.a(new_n266), .b(new_n274), .o1(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n271), .c(new_n270), .d(new_n266), .o1(\s[24] ));
  nano32aa1n02x5               g181(.a(new_n236), .b(new_n271), .c(new_n255), .d(new_n265), .out0(new_n277));
  and002aa1n18x5               g182(.a(new_n271), .b(new_n265), .o(new_n278));
  inv040aa1n03x5               g183(.a(new_n278), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(new_n273), .b(new_n272), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n279), .c(new_n261), .d(new_n263), .o1(new_n281));
  xnrc02aa1n12x5               g186(.a(\b[24] ), .b(\a[25] ), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n281), .c(new_n206), .d(new_n277), .o1(new_n284));
  aoi112aa1n02x5               g189(.a(new_n283), .b(new_n281), .c(new_n206), .d(new_n277), .o1(new_n285));
  norb02aa1n03x4               g190(.a(new_n284), .b(new_n285), .out0(\s[25] ));
  norp02aa1n02x5               g191(.a(\b[24] ), .b(\a[25] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  xorc02aa1n03x5               g193(.a(\a[26] ), .b(\b[25] ), .out0(new_n289));
  nanp02aa1n02x5               g194(.a(\b[25] ), .b(\a[26] ), .o1(new_n290));
  oai022aa1n02x5               g195(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n291));
  norb02aa1n02x5               g196(.a(new_n290), .b(new_n291), .out0(new_n292));
  nanp02aa1n03x5               g197(.a(new_n284), .b(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n288), .d(new_n284), .o1(\s[26] ));
  nanp03aa1n02x5               g199(.a(new_n164), .b(new_n197), .c(new_n195), .o1(new_n295));
  nanb02aa1n02x5               g200(.a(new_n200), .b(new_n295), .out0(new_n296));
  norb02aa1n06x4               g201(.a(new_n289), .b(new_n282), .out0(new_n297));
  inv000aa1n02x5               g202(.a(new_n297), .o1(new_n298));
  nano23aa1n06x5               g203(.a(new_n236), .b(new_n298), .c(new_n278), .d(new_n255), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n296), .c(new_n150), .d(new_n193), .o1(new_n300));
  aoi022aa1n06x5               g205(.a(new_n281), .b(new_n297), .c(new_n290), .d(new_n291), .o1(new_n301));
  xorc02aa1n12x5               g206(.a(\a[27] ), .b(\b[26] ), .out0(new_n302));
  xnbna2aa1n06x5               g207(.a(new_n302), .b(new_n301), .c(new_n300), .out0(\s[27] ));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n278), .b(new_n262), .c(new_n241), .d(new_n255), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(new_n291), .b(new_n290), .o1(new_n307));
  aoai13aa1n04x5               g212(.a(new_n307), .b(new_n298), .c(new_n306), .d(new_n280), .o1(new_n308));
  aoai13aa1n02x5               g213(.a(new_n302), .b(new_n308), .c(new_n206), .d(new_n299), .o1(new_n309));
  tech160nm_fixorc02aa1n03p5x5 g214(.a(\a[28] ), .b(\b[27] ), .out0(new_n310));
  inv000aa1d42x5               g215(.a(new_n302), .o1(new_n311));
  oai022aa1n02x5               g216(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n312));
  aoi012aa1n02x5               g217(.a(new_n312), .b(\a[28] ), .c(\b[27] ), .o1(new_n313));
  aoai13aa1n04x5               g218(.a(new_n313), .b(new_n311), .c(new_n301), .d(new_n300), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n310), .c(new_n309), .d(new_n305), .o1(\s[28] ));
  and002aa1n02x5               g220(.a(new_n310), .b(new_n302), .o(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n308), .c(new_n206), .d(new_n299), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n316), .o1(new_n318));
  aob012aa1n02x5               g223(.a(new_n312), .b(\b[27] ), .c(\a[28] ), .out0(new_n319));
  aoai13aa1n02x7               g224(.a(new_n319), .b(new_n318), .c(new_n301), .d(new_n300), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .out0(new_n321));
  norb02aa1n02x5               g226(.a(new_n319), .b(new_n321), .out0(new_n322));
  aoi022aa1n03x5               g227(.a(new_n320), .b(new_n321), .c(new_n317), .d(new_n322), .o1(\s[29] ));
  xnrb03aa1n02x5               g228(.a(new_n137), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g229(.a(new_n311), .b(new_n310), .c(new_n321), .out0(new_n325));
  aoai13aa1n02x5               g230(.a(new_n325), .b(new_n308), .c(new_n206), .d(new_n299), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n325), .o1(new_n327));
  oaoi03aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .c(new_n319), .o1(new_n328));
  inv000aa1n03x5               g233(.a(new_n328), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n327), .c(new_n301), .d(new_n300), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .out0(new_n331));
  norp02aa1n02x5               g236(.a(new_n328), .b(new_n331), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n326), .d(new_n332), .o1(\s[30] ));
  nano32aa1d15x5               g238(.a(new_n311), .b(new_n331), .c(new_n310), .d(new_n321), .out0(new_n334));
  aoai13aa1n02x5               g239(.a(new_n334), .b(new_n308), .c(new_n206), .d(new_n299), .o1(new_n335));
  inv000aa1d42x5               g240(.a(new_n334), .o1(new_n336));
  oao003aa1n02x5               g241(.a(\a[30] ), .b(\b[29] ), .c(new_n329), .carry(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n336), .c(new_n301), .d(new_n300), .o1(new_n338));
  xorc02aa1n02x5               g243(.a(\a[31] ), .b(\b[30] ), .out0(new_n339));
  norb02aa1n02x5               g244(.a(new_n337), .b(new_n339), .out0(new_n340));
  aoi022aa1n03x5               g245(.a(new_n338), .b(new_n339), .c(new_n335), .d(new_n340), .o1(\s[31] ));
  norb03aa1n02x5               g246(.a(new_n100), .b(new_n137), .c(new_n99), .out0(new_n342));
  inv000aa1d42x5               g247(.a(new_n104), .o1(new_n343));
  aoi012aa1n02x5               g248(.a(new_n99), .b(new_n343), .c(new_n105), .o1(new_n344));
  aboi22aa1n03x5               g249(.a(new_n342), .b(new_n344), .c(new_n138), .d(new_n140), .out0(\s[3] ));
  nanp02aa1n02x5               g250(.a(new_n138), .b(new_n140), .o1(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n139), .b(new_n346), .c(new_n343), .out0(\s[4] ));
  xnbna2aa1n03x5               g252(.a(new_n116), .b(new_n141), .c(new_n107), .out0(\s[5] ));
  aoi012aa1n02x5               g253(.a(new_n114), .b(new_n108), .c(new_n115), .o1(new_n349));
  norb03aa1n02x5               g254(.a(new_n118), .b(new_n114), .c(new_n117), .out0(new_n350));
  aob012aa1n02x5               g255(.a(new_n350), .b(new_n108), .c(new_n116), .out0(new_n351));
  oai012aa1n02x5               g256(.a(new_n351), .b(new_n349), .c(new_n119), .o1(\s[6] ));
  aoi022aa1n02x5               g257(.a(new_n351), .b(new_n118), .c(new_n146), .d(new_n110), .o1(new_n353));
  aoi013aa1n02x4               g258(.a(new_n353), .b(new_n351), .c(new_n121), .d(new_n146), .o1(\s[7] ));
  aoi022aa1n02x5               g259(.a(new_n351), .b(new_n121), .c(new_n144), .d(new_n145), .o1(new_n355));
  xnrb03aa1n02x5               g260(.a(new_n355), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g261(.a(new_n126), .b(new_n159), .c(new_n149), .out0(\s[9] ));
endmodule


