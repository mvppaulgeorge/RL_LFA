// Benchmark "adder" written by ABC on Wed Jul 17 20:37:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n321, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n339, new_n340, new_n342, new_n343, new_n345, new_n346,
    new_n348, new_n349, new_n350, new_n352, new_n353, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor022aa1n06x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  aoi022aa1d24x5               g003(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n99));
  norp02aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  norb02aa1n09x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  oai022aa1n12x5               g007(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  oaoi13aa1n12x5               g008(.a(new_n103), .b(new_n102), .c(new_n99), .d(new_n98), .o1(new_n104));
  nand02aa1n03x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  oai112aa1n02x5               g011(.a(new_n105), .b(new_n106), .c(\b[7] ), .d(\a[8] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[5] ), .o1(new_n108));
  nanb02aa1d24x5               g013(.a(\a[6] ), .b(new_n108), .out0(new_n109));
  nand02aa1d08x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nand02aa1d04x5               g015(.a(new_n109), .b(new_n110), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  oai012aa1n02x5               g017(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .o1(new_n113));
  nor042aa1n06x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  and002aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o(new_n115));
  nor043aa1n02x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nona22aa1n09x5               g021(.a(new_n116), .b(new_n111), .c(new_n107), .out0(new_n117));
  oai022aa1n02x5               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  oaih12aa1n02x5               g023(.a(new_n110), .b(\b[6] ), .c(\a[7] ), .o1(new_n119));
  oaih12aa1n02x5               g024(.a(new_n105), .b(\b[7] ), .c(\a[8] ), .o1(new_n120));
  nor042aa1n02x5               g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  oai022aa1n02x5               g026(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n122));
  aoai13aa1n04x5               g027(.a(new_n112), .b(new_n122), .c(new_n121), .d(new_n118), .o1(new_n123));
  oai012aa1d24x5               g028(.a(new_n123), .b(new_n117), .c(new_n104), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  xorc02aa1n12x5               g030(.a(\a[10] ), .b(\b[9] ), .out0(new_n126));
  aoai13aa1n09x5               g031(.a(new_n126), .b(new_n97), .c(new_n124), .d(new_n125), .o1(new_n127));
  aoi112aa1n02x7               g032(.a(new_n126), .b(new_n97), .c(new_n124), .d(new_n125), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n127), .b(new_n128), .out0(\s[10] ));
  inv000aa1n03x5               g034(.a(new_n97), .o1(new_n130));
  oaoi03aa1n02x5               g035(.a(\a[10] ), .b(\b[9] ), .c(new_n130), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nor002aa1n20x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  tech160nm_finand02aa1n05x5   g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n127), .c(new_n132), .out0(\s[11] ));
  nand02aa1n02x5               g041(.a(new_n127), .b(new_n132), .o1(new_n137));
  nand42aa1n02x5               g042(.a(new_n137), .b(new_n135), .o1(new_n138));
  nor022aa1n08x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand42aa1n06x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  aoib12aa1n02x5               g046(.a(new_n133), .b(new_n140), .c(new_n139), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n133), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n135), .o1(new_n144));
  aoai13aa1n03x5               g049(.a(new_n143), .b(new_n144), .c(new_n127), .d(new_n132), .o1(new_n145));
  aoi022aa1n03x5               g050(.a(new_n145), .b(new_n141), .c(new_n138), .d(new_n142), .o1(\s[12] ));
  nano23aa1n06x5               g051(.a(new_n133), .b(new_n139), .c(new_n140), .d(new_n134), .out0(new_n147));
  nand23aa1n06x5               g052(.a(new_n147), .b(new_n125), .c(new_n126), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  oai022aa1n02x5               g054(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n150));
  aoi022aa1n02x7               g055(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n151));
  aoi112aa1n06x5               g056(.a(new_n139), .b(new_n133), .c(new_n150), .d(new_n151), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n140), .b(new_n152), .out0(new_n153));
  tech160nm_fixorc02aa1n03p5x5 g058(.a(\a[13] ), .b(\b[12] ), .out0(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n153), .c(new_n124), .d(new_n149), .o1(new_n155));
  aoi112aa1n02x7               g060(.a(new_n154), .b(new_n153), .c(new_n124), .d(new_n149), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n155), .b(new_n156), .out0(\s[13] ));
  norp02aa1n24x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  tech160nm_fixorc02aa1n03p5x5 g064(.a(\a[14] ), .b(\b[13] ), .out0(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n155), .c(new_n159), .out0(\s[14] ));
  oaoi03aa1n02x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n159), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  and002aa1n02x5               g068(.a(new_n160), .b(new_n154), .o(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n153), .c(new_n124), .d(new_n149), .o1(new_n165));
  nor002aa1n20x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nand02aa1n08x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n165), .c(new_n163), .out0(\s[15] ));
  nand02aa1n02x5               g074(.a(new_n165), .b(new_n163), .o1(new_n170));
  nand42aa1n02x5               g075(.a(new_n170), .b(new_n168), .o1(new_n171));
  nor002aa1n03x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  norp02aa1n02x5               g079(.a(new_n174), .b(new_n166), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n166), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n167), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n176), .b(new_n177), .c(new_n165), .d(new_n163), .o1(new_n178));
  aoi022aa1n03x5               g083(.a(new_n178), .b(new_n174), .c(new_n171), .d(new_n175), .o1(\s[16] ));
  nano23aa1n06x5               g084(.a(new_n166), .b(new_n172), .c(new_n173), .d(new_n167), .out0(new_n180));
  nano32aa1d12x5               g085(.a(new_n148), .b(new_n180), .c(new_n154), .d(new_n160), .out0(new_n181));
  nanp02aa1n09x5               g086(.a(new_n124), .b(new_n181), .o1(new_n182));
  nanb03aa1n06x5               g087(.a(new_n172), .b(new_n173), .c(new_n167), .out0(new_n183));
  aoi012aa1n02x7               g088(.a(new_n158), .b(\a[12] ), .c(\b[11] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\a[14] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\b[13] ), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(new_n186), .b(new_n185), .c(\a[13] ), .d(\b[12] ), .o1(new_n187));
  aoi012aa1n02x7               g092(.a(new_n166), .b(\a[14] ), .c(\b[13] ), .o1(new_n188));
  nand03aa1n04x5               g093(.a(new_n187), .b(new_n184), .c(new_n188), .o1(new_n189));
  norp03aa1n02x5               g094(.a(new_n152), .b(new_n189), .c(new_n183), .o1(new_n190));
  aoi022aa1d24x5               g095(.a(\b[14] ), .b(\a[15] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n158), .c(new_n185), .d(new_n186), .o1(new_n192));
  norp02aa1n02x5               g097(.a(new_n172), .b(new_n166), .o1(new_n193));
  aoi022aa1n03x5               g098(.a(new_n192), .b(new_n193), .c(\b[15] ), .d(\a[16] ), .o1(new_n194));
  tech160nm_finor002aa1n03p5x5 g099(.a(new_n190), .b(new_n194), .o1(new_n195));
  nand02aa1d04x5               g100(.a(new_n182), .b(new_n195), .o1(new_n196));
  xorc02aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  norp03aa1n02x5               g102(.a(new_n190), .b(new_n194), .c(new_n197), .o1(new_n198));
  aoi022aa1n02x5               g103(.a(new_n196), .b(new_n197), .c(new_n182), .d(new_n198), .o1(\s[17] ));
  nor022aa1n08x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  inv000aa1n03x5               g105(.a(new_n200), .o1(new_n201));
  inv020aa1n02x5               g106(.a(new_n194), .o1(new_n202));
  oai013aa1n09x5               g107(.a(new_n202), .b(new_n152), .c(new_n189), .d(new_n183), .o1(new_n203));
  aoai13aa1n06x5               g108(.a(new_n197), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n204));
  xorc02aa1n02x5               g109(.a(\a[18] ), .b(\b[17] ), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n204), .c(new_n201), .out0(\s[18] ));
  oaoi03aa1n02x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n201), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  xnrc02aa1n02x5               g114(.a(\b[17] ), .b(\a[18] ), .out0(new_n210));
  nano22aa1n06x5               g115(.a(new_n210), .b(new_n201), .c(new_n209), .out0(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n212));
  xorc02aa1n12x5               g117(.a(\a[19] ), .b(\b[18] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n212), .c(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n04x5               g120(.a(new_n213), .b(new_n207), .c(new_n196), .d(new_n211), .o1(new_n216));
  nor002aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  tech160nm_finand02aa1n03p5x5 g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n06x4               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  norp02aa1n02x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  aoib12aa1n02x5               g125(.a(new_n220), .b(new_n218), .c(new_n217), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n220), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n213), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n222), .b(new_n223), .c(new_n212), .d(new_n208), .o1(new_n224));
  aoi022aa1n03x5               g129(.a(new_n224), .b(new_n219), .c(new_n216), .d(new_n221), .o1(\s[20] ));
  nand23aa1n06x5               g130(.a(new_n211), .b(new_n213), .c(new_n219), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n228));
  oaih22aa1d12x5               g133(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n229));
  aoi022aa1n06x5               g134(.a(\b[18] ), .b(\a[19] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n230));
  oai022aa1n02x7               g135(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n231));
  aoi012aa1n06x5               g136(.a(new_n231), .b(new_n229), .c(new_n230), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n218), .b(new_n232), .out0(new_n233));
  inv000aa1n02x5               g138(.a(new_n233), .o1(new_n234));
  xorc02aa1n12x5               g139(.a(\a[21] ), .b(\b[20] ), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n228), .c(new_n234), .out0(\s[21] ));
  aoai13aa1n04x5               g141(.a(new_n235), .b(new_n233), .c(new_n196), .d(new_n227), .o1(new_n237));
  xorc02aa1n02x5               g142(.a(\a[22] ), .b(\b[21] ), .out0(new_n238));
  nor002aa1d32x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  norp02aa1n02x5               g144(.a(new_n238), .b(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n239), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n235), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n241), .b(new_n242), .c(new_n228), .d(new_n234), .o1(new_n243));
  aoi022aa1n03x5               g148(.a(new_n243), .b(new_n238), .c(new_n237), .d(new_n240), .o1(\s[22] ));
  inv000aa1d42x5               g149(.a(\a[21] ), .o1(new_n245));
  inv040aa1d32x5               g150(.a(\a[22] ), .o1(new_n246));
  xroi22aa1d04x5               g151(.a(new_n245), .b(\b[20] ), .c(new_n246), .d(\b[21] ), .out0(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n226), .out0(new_n248));
  aoai13aa1n04x5               g153(.a(new_n248), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[21] ), .b(\a[22] ), .o1(new_n250));
  tech160nm_fiaoi012aa1n04x5   g155(.a(new_n239), .b(\a[20] ), .c(\b[19] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\b[21] ), .o1(new_n252));
  aoi022aa1n02x7               g157(.a(new_n252), .b(new_n246), .c(\a[21] ), .d(\b[20] ), .o1(new_n253));
  nand23aa1n03x5               g158(.a(new_n253), .b(new_n251), .c(new_n250), .o1(new_n254));
  oaoi03aa1n03x5               g159(.a(new_n246), .b(new_n252), .c(new_n239), .o1(new_n255));
  oai012aa1n12x5               g160(.a(new_n255), .b(new_n254), .c(new_n232), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  nand02aa1n02x5               g162(.a(new_n249), .b(new_n257), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  oai112aa1n02x5               g165(.a(new_n255), .b(new_n260), .c(new_n254), .d(new_n232), .o1(new_n261));
  aboi22aa1n03x5               g166(.a(new_n261), .b(new_n249), .c(new_n258), .d(new_n259), .out0(\s[23] ));
  tech160nm_finand02aa1n03p5x5 g167(.a(new_n258), .b(new_n259), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .out0(new_n264));
  nor042aa1n12x5               g169(.a(\b[22] ), .b(\a[23] ), .o1(new_n265));
  norp02aa1n02x5               g170(.a(new_n264), .b(new_n265), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n265), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n260), .c(new_n249), .d(new_n257), .o1(new_n268));
  aoi022aa1n03x5               g173(.a(new_n268), .b(new_n264), .c(new_n263), .d(new_n266), .o1(\s[24] ));
  nanp02aa1n02x5               g174(.a(\b[22] ), .b(\a[23] ), .o1(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[23] ), .b(\a[24] ), .out0(new_n271));
  nano22aa1n06x5               g176(.a(new_n271), .b(new_n267), .c(new_n270), .out0(new_n272));
  nano22aa1n03x7               g177(.a(new_n226), .b(new_n247), .c(new_n272), .out0(new_n273));
  aoai13aa1n04x5               g178(.a(new_n273), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n274));
  oaoi03aa1n12x5               g179(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .o1(new_n275));
  aoi012aa1n02x5               g180(.a(new_n275), .b(new_n256), .c(new_n272), .o1(new_n276));
  nand02aa1d04x5               g181(.a(new_n274), .b(new_n276), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  nanp02aa1n02x5               g183(.a(new_n264), .b(new_n259), .o1(new_n279));
  oaoi13aa1n02x5               g184(.a(new_n279), .b(new_n255), .c(new_n254), .d(new_n232), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n275), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n278), .o1(new_n282));
  nano22aa1n02x4               g187(.a(new_n280), .b(new_n281), .c(new_n282), .out0(new_n283));
  aoi022aa1n02x5               g188(.a(new_n277), .b(new_n278), .c(new_n274), .d(new_n283), .o1(\s[25] ));
  tech160nm_finand02aa1n03p5x5 g189(.a(new_n277), .b(new_n278), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .out0(new_n286));
  nor042aa1d18x5               g191(.a(\b[24] ), .b(\a[25] ), .o1(new_n287));
  norp02aa1n02x5               g192(.a(new_n286), .b(new_n287), .o1(new_n288));
  inv040aa1n08x5               g193(.a(new_n287), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n282), .c(new_n274), .d(new_n276), .o1(new_n290));
  aoi022aa1n03x5               g195(.a(new_n290), .b(new_n286), .c(new_n285), .d(new_n288), .o1(\s[26] ));
  nanp02aa1n02x5               g196(.a(\b[24] ), .b(\a[25] ), .o1(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[25] ), .b(\a[26] ), .out0(new_n293));
  nano22aa1n02x4               g198(.a(new_n293), .b(new_n289), .c(new_n292), .out0(new_n294));
  nano32aa1n03x7               g199(.a(new_n226), .b(new_n294), .c(new_n247), .d(new_n272), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n294), .b(new_n275), .c(new_n256), .d(new_n272), .o1(new_n296));
  oaoi03aa1n02x5               g201(.a(\a[26] ), .b(\b[25] ), .c(new_n289), .o1(new_n297));
  inv000aa1n02x5               g202(.a(new_n297), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n296), .b(new_n298), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  aoai13aa1n04x5               g205(.a(new_n300), .b(new_n299), .c(new_n196), .d(new_n295), .o1(new_n301));
  aoai13aa1n12x5               g206(.a(new_n295), .b(new_n203), .c(new_n124), .d(new_n181), .o1(new_n302));
  nano32aa1n03x7               g207(.a(new_n300), .b(new_n302), .c(new_n296), .d(new_n298), .out0(new_n303));
  norb02aa1n03x4               g208(.a(new_n301), .b(new_n303), .out0(\s[27] ));
  xorc02aa1n02x5               g209(.a(\a[28] ), .b(\b[27] ), .out0(new_n305));
  norp02aa1n02x5               g210(.a(\b[26] ), .b(\a[27] ), .o1(new_n306));
  norp02aa1n02x5               g211(.a(new_n305), .b(new_n306), .o1(new_n307));
  oaoi13aa1n02x7               g212(.a(new_n297), .b(new_n294), .c(new_n280), .d(new_n275), .o1(new_n308));
  inv000aa1n03x5               g213(.a(new_n306), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n300), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n309), .b(new_n310), .c(new_n308), .d(new_n302), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n311), .b(new_n305), .c(new_n301), .d(new_n307), .o1(\s[28] ));
  and002aa1n02x5               g217(.a(new_n305), .b(new_n300), .o(new_n313));
  aoai13aa1n02x7               g218(.a(new_n313), .b(new_n299), .c(new_n196), .d(new_n295), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .c(new_n309), .carry(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n308), .d(new_n302), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n316), .b(new_n318), .out0(new_n319));
  aoi022aa1n03x5               g224(.a(new_n317), .b(new_n318), .c(new_n314), .d(new_n319), .o1(\s[29] ));
  nanp02aa1n02x5               g225(.a(\b[0] ), .b(\a[1] ), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g227(.a(new_n310), .b(new_n305), .c(new_n318), .out0(new_n323));
  aoai13aa1n02x7               g228(.a(new_n323), .b(new_n299), .c(new_n196), .d(new_n295), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .carry(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n325), .c(new_n308), .d(new_n302), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .out0(new_n328));
  norb02aa1n02x5               g233(.a(new_n326), .b(new_n328), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n324), .d(new_n329), .o1(\s[30] ));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  nano32aa1n03x7               g236(.a(new_n310), .b(new_n328), .c(new_n305), .d(new_n318), .out0(new_n332));
  aoai13aa1n02x7               g237(.a(new_n332), .b(new_n299), .c(new_n196), .d(new_n295), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n332), .o1(new_n334));
  oao003aa1n02x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n334), .c(new_n308), .d(new_n302), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n335), .b(new_n331), .out0(new_n337));
  aoi022aa1n03x5               g242(.a(new_n336), .b(new_n331), .c(new_n333), .d(new_n337), .o1(\s[31] ));
  oai012aa1n02x5               g243(.a(new_n102), .b(new_n99), .c(new_n98), .o1(new_n339));
  norp03aa1n02x5               g244(.a(new_n102), .b(new_n99), .c(new_n98), .o1(new_n340));
  norb02aa1n02x5               g245(.a(new_n339), .b(new_n340), .out0(\s[3] ));
  xorc02aa1n02x5               g246(.a(\a[4] ), .b(\b[3] ), .out0(new_n342));
  norp02aa1n02x5               g247(.a(new_n342), .b(new_n100), .o1(new_n343));
  aboi22aa1n03x5               g248(.a(new_n104), .b(new_n342), .c(new_n343), .d(new_n339), .out0(\s[4] ));
  inv000aa1d42x5               g249(.a(new_n104), .o1(new_n345));
  norp02aa1n02x5               g250(.a(new_n115), .b(new_n114), .o1(new_n346));
  xobna2aa1n03x5               g251(.a(new_n346), .b(new_n345), .c(new_n106), .out0(\s[5] ));
  inv000aa1d42x5               g252(.a(new_n111), .o1(new_n348));
  inv000aa1d42x5               g253(.a(new_n114), .o1(new_n349));
  nanb03aa1n03x5               g254(.a(new_n104), .b(new_n346), .c(new_n106), .out0(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n348), .b(new_n350), .c(new_n349), .out0(\s[6] ));
  aob012aa1n02x5               g256(.a(new_n348), .b(new_n350), .c(new_n349), .out0(new_n352));
  xorc02aa1n02x5               g257(.a(\a[7] ), .b(\b[6] ), .out0(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n353), .b(new_n352), .c(new_n109), .out0(\s[7] ));
  aoai13aa1n02x5               g259(.a(new_n109), .b(new_n111), .c(new_n350), .d(new_n349), .o1(new_n355));
  nanp02aa1n03x5               g260(.a(new_n355), .b(new_n353), .o1(new_n356));
  inv000aa1d42x5               g261(.a(\a[7] ), .o1(new_n357));
  oaib12aa1n02x5               g262(.a(new_n356), .b(\b[6] ), .c(new_n357), .out0(new_n358));
  xorc02aa1n02x5               g263(.a(\a[8] ), .b(\b[7] ), .out0(new_n359));
  aoib12aa1n02x5               g264(.a(new_n359), .b(new_n357), .c(\b[6] ), .out0(new_n360));
  aoi022aa1n02x5               g265(.a(new_n358), .b(new_n359), .c(new_n356), .d(new_n360), .o1(\s[8] ));
  oab012aa1n02x4               g266(.a(new_n125), .b(new_n117), .c(new_n104), .out0(new_n362));
  aoi022aa1n02x5               g267(.a(new_n362), .b(new_n123), .c(new_n124), .d(new_n125), .o1(\s[9] ));
endmodule


