// Benchmark "adder" written by ABC on Thu Jul 18 11:40:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n344,
    new_n345, new_n347, new_n350, new_n351, new_n353, new_n355, new_n357;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n03x5               g001(.a(\a[3] ), .b(\b[2] ), .o(new_n97));
  oao003aa1n09x5               g002(.a(\a[4] ), .b(\b[3] ), .c(new_n97), .carry(new_n98));
  nor022aa1n16x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nand42aa1n08x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand02aa1d28x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nanb03aa1n12x5               g006(.a(new_n99), .b(new_n101), .c(new_n100), .out0(new_n102));
  nand02aa1d06x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor042aa1n03x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nona22aa1n03x5               g009(.a(new_n101), .b(new_n104), .c(new_n103), .out0(new_n105));
  tech160nm_fixorc02aa1n03p5x5 g010(.a(\a[4] ), .b(\b[3] ), .out0(new_n106));
  nanb03aa1n06x5               g011(.a(new_n102), .b(new_n106), .c(new_n105), .out0(new_n107));
  xnrc02aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .out0(new_n108));
  tech160nm_fixorc02aa1n05x5   g013(.a(\a[5] ), .b(\b[4] ), .out0(new_n109));
  xorc02aa1n12x5               g014(.a(\a[8] ), .b(\b[7] ), .out0(new_n110));
  nor022aa1n16x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n06x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanb02aa1n02x5               g017(.a(new_n111), .b(new_n112), .out0(new_n113));
  nona23aa1n08x5               g018(.a(new_n109), .b(new_n110), .c(new_n108), .d(new_n113), .out0(new_n114));
  nand42aa1n03x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nano22aa1n03x5               g020(.a(new_n111), .b(new_n115), .c(new_n112), .out0(new_n116));
  oai022aa1n03x5               g021(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\a[7] ), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(\b[6] ), .b(new_n118), .out0(new_n119));
  oaoi03aa1n03x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  aoi013aa1n06x4               g025(.a(new_n120), .b(new_n116), .c(new_n110), .d(new_n117), .o1(new_n121));
  aoai13aa1n12x5               g026(.a(new_n121), .b(new_n114), .c(new_n107), .d(new_n98), .o1(new_n122));
  nor042aa1n09x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  xorc02aa1n12x5               g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  nor042aa1n09x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nanp02aa1n12x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  norb02aa1n06x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  aoi112aa1n02x5               g032(.a(new_n123), .b(new_n127), .c(new_n122), .d(new_n124), .o1(new_n128));
  aoai13aa1n06x5               g033(.a(new_n127), .b(new_n123), .c(new_n122), .d(new_n124), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(\s[10] ));
  oai012aa1n02x5               g035(.a(new_n126), .b(new_n125), .c(new_n123), .o1(new_n131));
  nor002aa1d32x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1d28x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n129), .c(new_n131), .out0(\s[11] ));
  nanp02aa1n06x5               g040(.a(new_n129), .b(new_n131), .o1(new_n136));
  nanp02aa1n03x5               g041(.a(new_n136), .b(new_n134), .o1(new_n137));
  nor002aa1n20x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand42aa1d28x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  inv000aa1d42x5               g045(.a(new_n138), .o1(new_n141));
  aoi012aa1n02x5               g046(.a(new_n132), .b(new_n141), .c(new_n139), .o1(new_n142));
  inv040aa1n03x5               g047(.a(new_n132), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n134), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n143), .b(new_n144), .c(new_n129), .d(new_n131), .o1(new_n145));
  aoi022aa1n03x5               g050(.a(new_n145), .b(new_n140), .c(new_n137), .d(new_n142), .o1(\s[12] ));
  norb03aa1n02x7               g051(.a(new_n101), .b(new_n104), .c(new_n103), .out0(new_n147));
  xnrc02aa1n02x5               g052(.a(\b[3] ), .b(\a[4] ), .out0(new_n148));
  oai013aa1n03x5               g053(.a(new_n98), .b(new_n147), .c(new_n102), .d(new_n148), .o1(new_n149));
  xorc02aa1n02x5               g054(.a(\a[6] ), .b(\b[5] ), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n109), .b(new_n150), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n112), .b(new_n111), .out0(new_n152));
  nano22aa1n03x7               g057(.a(new_n151), .b(new_n110), .c(new_n152), .out0(new_n153));
  nanp03aa1n02x5               g058(.a(new_n116), .b(new_n110), .c(new_n117), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n120), .b(new_n154), .out0(new_n155));
  nano23aa1d12x5               g060(.a(new_n132), .b(new_n138), .c(new_n139), .d(new_n133), .out0(new_n156));
  nand23aa1n09x5               g061(.a(new_n156), .b(new_n124), .c(new_n127), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n155), .c(new_n149), .d(new_n153), .o1(new_n159));
  nanb03aa1d24x5               g064(.a(new_n138), .b(new_n139), .c(new_n133), .out0(new_n160));
  oai112aa1n06x5               g065(.a(new_n143), .b(new_n126), .c(new_n125), .d(new_n123), .o1(new_n161));
  aoi012aa1d24x5               g066(.a(new_n138), .b(new_n132), .c(new_n139), .o1(new_n162));
  oai012aa1d24x5               g067(.a(new_n162), .b(new_n161), .c(new_n160), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  nor042aa1n04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand42aa1n06x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n159), .c(new_n164), .out0(\s[13] ));
  orn002aa1n02x5               g073(.a(\a[13] ), .b(\b[12] ), .o(new_n169));
  aoai13aa1n02x5               g074(.a(new_n167), .b(new_n163), .c(new_n122), .d(new_n158), .o1(new_n170));
  nor042aa1n04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1n16x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n170), .c(new_n169), .out0(\s[14] ));
  nano23aa1d15x5               g079(.a(new_n165), .b(new_n171), .c(new_n172), .d(new_n166), .out0(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n163), .c(new_n122), .d(new_n158), .o1(new_n176));
  aoi012aa1d18x5               g081(.a(new_n171), .b(new_n165), .c(new_n172), .o1(new_n177));
  xorc02aa1n12x5               g082(.a(\a[15] ), .b(\b[14] ), .out0(new_n178));
  xnbna2aa1n03x5               g083(.a(new_n178), .b(new_n176), .c(new_n177), .out0(\s[15] ));
  nand42aa1n03x5               g084(.a(new_n159), .b(new_n164), .o1(new_n180));
  inv000aa1d42x5               g085(.a(new_n177), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n178), .b(new_n181), .c(new_n180), .d(new_n175), .o1(new_n182));
  tech160nm_fixorc02aa1n04x5   g087(.a(\a[16] ), .b(\b[15] ), .out0(new_n183));
  nor042aa1n06x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norp02aa1n02x5               g089(.a(new_n183), .b(new_n184), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n184), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n178), .o1(new_n187));
  aoai13aa1n03x5               g092(.a(new_n186), .b(new_n187), .c(new_n176), .d(new_n177), .o1(new_n188));
  aoi022aa1n02x5               g093(.a(new_n188), .b(new_n183), .c(new_n182), .d(new_n185), .o1(\s[16] ));
  nano32aa1d12x5               g094(.a(new_n157), .b(new_n183), .c(new_n175), .d(new_n178), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n155), .c(new_n149), .d(new_n153), .o1(new_n191));
  and002aa1n03x5               g096(.a(new_n183), .b(new_n178), .o(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n181), .c(new_n163), .d(new_n175), .o1(new_n193));
  oao003aa1n02x5               g098(.a(\a[16] ), .b(\b[15] ), .c(new_n186), .carry(new_n194));
  nand23aa1n06x5               g099(.a(new_n191), .b(new_n193), .c(new_n194), .o1(new_n195));
  xorc02aa1n12x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  nano22aa1n02x4               g101(.a(new_n196), .b(new_n193), .c(new_n194), .out0(new_n197));
  aoi022aa1n02x5               g102(.a(new_n195), .b(new_n196), .c(new_n197), .d(new_n191), .o1(\s[17] ));
  inv000aa1d42x5               g103(.a(\a[17] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(\b[16] ), .b(new_n199), .out0(new_n200));
  inv020aa1n04x5               g105(.a(new_n192), .o1(new_n201));
  nano22aa1n02x4               g106(.a(new_n138), .b(new_n133), .c(new_n139), .out0(new_n202));
  oai012aa1n02x5               g107(.a(new_n126), .b(\b[10] ), .c(\a[11] ), .o1(new_n203));
  oab012aa1n04x5               g108(.a(new_n203), .b(new_n123), .c(new_n125), .out0(new_n204));
  inv000aa1n02x5               g109(.a(new_n162), .o1(new_n205));
  aoai13aa1n04x5               g110(.a(new_n175), .b(new_n205), .c(new_n204), .d(new_n202), .o1(new_n206));
  aoai13aa1n12x5               g111(.a(new_n194), .b(new_n201), .c(new_n206), .d(new_n177), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n196), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n208));
  nor042aa1d18x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nand42aa1n10x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  norb02aa1n09x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n208), .c(new_n200), .out0(\s[18] ));
  and002aa1n02x5               g117(.a(new_n196), .b(new_n211), .o(new_n213));
  aoai13aa1n06x5               g118(.a(new_n213), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n214));
  oaoi03aa1n02x5               g119(.a(\a[18] ), .b(\b[17] ), .c(new_n200), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  nor042aa1d18x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nand42aa1n06x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  norb02aa1n12x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n214), .c(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g125(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g126(.a(new_n219), .b(new_n215), .c(new_n195), .d(new_n213), .o1(new_n222));
  nor002aa1d32x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nand42aa1n20x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  inv000aa1d42x5               g130(.a(\a[19] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[18] ), .o1(new_n227));
  aboi22aa1n03x5               g132(.a(new_n223), .b(new_n224), .c(new_n226), .d(new_n227), .out0(new_n228));
  inv040aa1n03x5               g133(.a(new_n217), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n219), .o1(new_n230));
  aoai13aa1n02x5               g135(.a(new_n229), .b(new_n230), .c(new_n214), .d(new_n216), .o1(new_n231));
  aoi022aa1n03x5               g136(.a(new_n231), .b(new_n225), .c(new_n222), .d(new_n228), .o1(\s[20] ));
  nano32aa1n03x7               g137(.a(new_n230), .b(new_n196), .c(new_n225), .d(new_n211), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n234));
  nanb03aa1n09x5               g139(.a(new_n223), .b(new_n224), .c(new_n218), .out0(new_n235));
  nor042aa1n04x5               g140(.a(\b[16] ), .b(\a[17] ), .o1(new_n236));
  oai112aa1n06x5               g141(.a(new_n229), .b(new_n210), .c(new_n209), .d(new_n236), .o1(new_n237));
  aoi012aa1d24x5               g142(.a(new_n223), .b(new_n217), .c(new_n224), .o1(new_n238));
  oaih12aa1n12x5               g143(.a(new_n238), .b(new_n237), .c(new_n235), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nor002aa1n20x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  nand42aa1n06x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  norb02aa1n06x4               g147(.a(new_n242), .b(new_n241), .out0(new_n243));
  xnbna2aa1n03x5               g148(.a(new_n243), .b(new_n234), .c(new_n240), .out0(\s[21] ));
  aoai13aa1n03x5               g149(.a(new_n243), .b(new_n239), .c(new_n195), .d(new_n233), .o1(new_n245));
  nor042aa1n06x5               g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  nand42aa1n20x5               g151(.a(\b[21] ), .b(\a[22] ), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  aoib12aa1n02x5               g153(.a(new_n241), .b(new_n247), .c(new_n246), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n241), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n243), .o1(new_n251));
  aoai13aa1n02x5               g156(.a(new_n250), .b(new_n251), .c(new_n234), .d(new_n240), .o1(new_n252));
  aoi022aa1n03x5               g157(.a(new_n252), .b(new_n248), .c(new_n245), .d(new_n249), .o1(\s[22] ));
  inv020aa1n02x5               g158(.a(new_n233), .o1(new_n254));
  nano22aa1n02x4               g159(.a(new_n254), .b(new_n243), .c(new_n248), .out0(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n256));
  nano23aa1d12x5               g161(.a(new_n241), .b(new_n246), .c(new_n247), .d(new_n242), .out0(new_n257));
  aoi012aa1d18x5               g162(.a(new_n246), .b(new_n241), .c(new_n247), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  tech160nm_fiaoi012aa1n03p5x5 g164(.a(new_n259), .b(new_n239), .c(new_n257), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(new_n256), .b(new_n260), .o1(new_n261));
  xorc02aa1n12x5               g166(.a(\a[23] ), .b(\b[22] ), .out0(new_n262));
  aoi112aa1n02x5               g167(.a(new_n262), .b(new_n259), .c(new_n239), .d(new_n257), .o1(new_n263));
  aoi022aa1n02x5               g168(.a(new_n261), .b(new_n262), .c(new_n256), .d(new_n263), .o1(\s[23] ));
  inv000aa1n02x5               g169(.a(new_n260), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n262), .b(new_n265), .c(new_n195), .d(new_n255), .o1(new_n266));
  tech160nm_fixorc02aa1n02p5x5 g171(.a(\a[24] ), .b(\b[23] ), .out0(new_n267));
  nor042aa1n06x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n267), .b(new_n268), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n268), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n262), .o1(new_n271));
  aoai13aa1n02x7               g176(.a(new_n270), .b(new_n271), .c(new_n256), .d(new_n260), .o1(new_n272));
  aoi022aa1n02x7               g177(.a(new_n272), .b(new_n267), .c(new_n266), .d(new_n269), .o1(\s[24] ));
  and002aa1n12x5               g178(.a(new_n267), .b(new_n262), .o(new_n274));
  nano22aa1n02x4               g179(.a(new_n254), .b(new_n274), .c(new_n257), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n276));
  nano22aa1n02x4               g181(.a(new_n223), .b(new_n218), .c(new_n224), .out0(new_n277));
  oaih12aa1n02x5               g182(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .o1(new_n278));
  oab012aa1n02x4               g183(.a(new_n278), .b(new_n236), .c(new_n209), .out0(new_n279));
  inv000aa1n02x5               g184(.a(new_n238), .o1(new_n280));
  aoai13aa1n04x5               g185(.a(new_n257), .b(new_n280), .c(new_n279), .d(new_n277), .o1(new_n281));
  inv000aa1n06x5               g186(.a(new_n274), .o1(new_n282));
  oao003aa1n02x5               g187(.a(\a[24] ), .b(\b[23] ), .c(new_n270), .carry(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n282), .c(new_n281), .d(new_n258), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n276), .b(new_n285), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[25] ), .b(\b[24] ), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n274), .b(new_n259), .c(new_n239), .d(new_n257), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n287), .o1(new_n289));
  and003aa1n02x5               g194(.a(new_n288), .b(new_n289), .c(new_n283), .o(new_n290));
  aoi022aa1n02x5               g195(.a(new_n286), .b(new_n287), .c(new_n276), .d(new_n290), .o1(\s[25] ));
  aoai13aa1n03x5               g196(.a(new_n287), .b(new_n284), .c(new_n195), .d(new_n275), .o1(new_n292));
  xorc02aa1n03x5               g197(.a(\a[26] ), .b(\b[25] ), .out0(new_n293));
  nor042aa1n03x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  norp02aa1n02x5               g199(.a(new_n293), .b(new_n294), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n294), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n289), .c(new_n276), .d(new_n285), .o1(new_n297));
  aoi022aa1n02x7               g202(.a(new_n297), .b(new_n293), .c(new_n292), .d(new_n295), .o1(\s[26] ));
  and002aa1n12x5               g203(.a(new_n293), .b(new_n287), .o(new_n299));
  nano32aa1n03x7               g204(.a(new_n254), .b(new_n299), .c(new_n257), .d(new_n274), .out0(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n207), .c(new_n122), .d(new_n190), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[26] ), .b(\b[25] ), .c(new_n296), .carry(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  aoi012aa1d18x5               g208(.a(new_n303), .b(new_n284), .c(new_n299), .o1(new_n304));
  nanp02aa1n02x5               g209(.a(new_n301), .b(new_n304), .o1(new_n305));
  xorc02aa1n12x5               g210(.a(\a[27] ), .b(\b[26] ), .out0(new_n306));
  aoi112aa1n02x5               g211(.a(new_n306), .b(new_n303), .c(new_n284), .d(new_n299), .o1(new_n307));
  aoi022aa1n02x5               g212(.a(new_n305), .b(new_n306), .c(new_n301), .d(new_n307), .o1(\s[27] ));
  inv000aa1d42x5               g213(.a(new_n299), .o1(new_n309));
  aoai13aa1n04x5               g214(.a(new_n302), .b(new_n309), .c(new_n288), .d(new_n283), .o1(new_n310));
  aoai13aa1n02x5               g215(.a(new_n306), .b(new_n310), .c(new_n195), .d(new_n300), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[28] ), .b(\b[27] ), .out0(new_n312));
  norp02aa1n02x5               g217(.a(\b[26] ), .b(\a[27] ), .o1(new_n313));
  norp02aa1n02x5               g218(.a(new_n312), .b(new_n313), .o1(new_n314));
  inv000aa1n03x5               g219(.a(new_n313), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n306), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n315), .b(new_n316), .c(new_n301), .d(new_n304), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n312), .c(new_n311), .d(new_n314), .o1(\s[28] ));
  and002aa1n02x5               g223(.a(new_n312), .b(new_n306), .o(new_n319));
  aoai13aa1n02x5               g224(.a(new_n319), .b(new_n310), .c(new_n195), .d(new_n300), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n319), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[28] ), .b(\b[27] ), .c(new_n315), .carry(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n321), .c(new_n301), .d(new_n304), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[29] ), .b(\b[28] ), .out0(new_n324));
  norb02aa1n02x5               g229(.a(new_n322), .b(new_n324), .out0(new_n325));
  aoi022aa1n03x5               g230(.a(new_n323), .b(new_n324), .c(new_n320), .d(new_n325), .o1(\s[29] ));
  xorb03aa1n02x5               g231(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g232(.a(new_n316), .b(new_n312), .c(new_n324), .out0(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n310), .c(new_n195), .d(new_n300), .o1(new_n329));
  inv000aa1n02x5               g234(.a(new_n328), .o1(new_n330));
  oao003aa1n02x5               g235(.a(\a[29] ), .b(\b[28] ), .c(new_n322), .carry(new_n331));
  aoai13aa1n03x5               g236(.a(new_n331), .b(new_n330), .c(new_n301), .d(new_n304), .o1(new_n332));
  xorc02aa1n02x5               g237(.a(\a[30] ), .b(\b[29] ), .out0(new_n333));
  norb02aa1n02x5               g238(.a(new_n331), .b(new_n333), .out0(new_n334));
  aoi022aa1n03x5               g239(.a(new_n332), .b(new_n333), .c(new_n329), .d(new_n334), .o1(\s[30] ));
  nano32aa1n06x5               g240(.a(new_n316), .b(new_n333), .c(new_n312), .d(new_n324), .out0(new_n336));
  aoai13aa1n02x5               g241(.a(new_n336), .b(new_n310), .c(new_n195), .d(new_n300), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[31] ), .b(\b[30] ), .out0(new_n338));
  oao003aa1n02x5               g243(.a(\a[30] ), .b(\b[29] ), .c(new_n331), .carry(new_n339));
  norb02aa1n02x5               g244(.a(new_n339), .b(new_n338), .out0(new_n340));
  inv000aa1d42x5               g245(.a(new_n336), .o1(new_n341));
  aoai13aa1n03x5               g246(.a(new_n339), .b(new_n341), .c(new_n301), .d(new_n304), .o1(new_n342));
  aoi022aa1n03x5               g247(.a(new_n342), .b(new_n338), .c(new_n337), .d(new_n340), .o1(\s[31] ));
  oai012aa1n02x5               g248(.a(new_n101), .b(new_n104), .c(new_n103), .o1(new_n344));
  nanb02aa1n02x5               g249(.a(new_n99), .b(new_n100), .out0(new_n345));
  aboi22aa1n03x5               g250(.a(new_n102), .b(new_n105), .c(new_n344), .d(new_n345), .out0(\s[3] ));
  aoi113aa1n02x5               g251(.a(new_n99), .b(new_n106), .c(new_n105), .d(new_n101), .e(new_n100), .o1(new_n347));
  oaoi13aa1n02x5               g252(.a(new_n347), .b(new_n149), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g253(.a(new_n109), .b(new_n107), .c(new_n98), .out0(\s[5] ));
  orn002aa1n02x5               g254(.a(\a[5] ), .b(\b[4] ), .o(new_n350));
  nanp02aa1n02x5               g255(.a(new_n149), .b(new_n109), .o1(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n150), .b(new_n351), .c(new_n350), .out0(\s[6] ));
  aboi22aa1n03x5               g257(.a(new_n151), .b(new_n149), .c(new_n117), .d(new_n115), .out0(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n353), .b(new_n119), .c(new_n112), .out0(\s[7] ));
  nanb02aa1n02x5               g259(.a(new_n353), .b(new_n152), .out0(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n110), .b(new_n355), .c(new_n119), .out0(\s[8] ));
  aoi112aa1n02x5               g261(.a(new_n124), .b(new_n155), .c(new_n149), .d(new_n153), .o1(new_n357));
  aoi012aa1n02x5               g262(.a(new_n357), .b(new_n122), .c(new_n124), .o1(\s[9] ));
endmodule


