// Benchmark "adder" written by ABC on Wed Jul 17 13:02:28 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n216, new_n217, new_n218, new_n219, new_n220, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n309,
    new_n311, new_n312, new_n315, new_n317, new_n318, new_n319, new_n321,
    new_n322, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  nor042aa1n04x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nand42aa1n02x5               g003(.a(\b[8] ), .b(\a[9] ), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norb02aa1n06x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  nanp02aa1n04x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nor042aa1n12x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano22aa1n03x7               g010(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n106));
  nand22aa1n09x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  nor002aa1n03x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nona22aa1n09x5               g013(.a(new_n103), .b(new_n108), .c(new_n107), .out0(new_n109));
  nand23aa1n06x5               g014(.a(new_n106), .b(new_n109), .c(new_n102), .o1(new_n110));
  tech160nm_fioai012aa1n03p5x5 g015(.a(new_n101), .b(new_n104), .c(new_n100), .o1(new_n111));
  nor002aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1d28x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor042aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n10x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n09x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  tech160nm_fixorc02aa1n04x5   g021(.a(\a[6] ), .b(\b[5] ), .out0(new_n117));
  tech160nm_fixorc02aa1n05x5   g022(.a(\a[5] ), .b(\b[4] ), .out0(new_n118));
  nand23aa1n03x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .o1(new_n119));
  orn002aa1n24x5               g024(.a(\a[5] ), .b(\b[4] ), .o(new_n120));
  oaoi03aa1n09x5               g025(.a(\a[6] ), .b(\b[5] ), .c(new_n120), .o1(new_n121));
  nona22aa1n09x5               g026(.a(new_n113), .b(new_n114), .c(new_n112), .out0(new_n122));
  aoi022aa1n09x5               g027(.a(new_n116), .b(new_n121), .c(new_n113), .d(new_n122), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n123), .b(new_n119), .c(new_n110), .d(new_n111), .o1(new_n124));
  aoai13aa1n02x5               g029(.a(new_n97), .b(new_n98), .c(new_n124), .d(new_n99), .o1(new_n125));
  nor042aa1n02x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  and002aa1n06x5               g031(.a(\b[9] ), .b(\a[10] ), .o(new_n127));
  norp03aa1n02x5               g032(.a(new_n127), .b(new_n98), .c(new_n126), .o1(new_n128));
  aob012aa1n06x5               g033(.a(new_n128), .b(new_n124), .c(new_n99), .out0(new_n129));
  nanp02aa1n02x5               g034(.a(new_n125), .b(new_n129), .o1(\s[10] ));
  nand42aa1n20x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor002aa1n16x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb03aa1n02x5               g037(.a(new_n131), .b(new_n127), .c(new_n132), .out0(new_n133));
  norb02aa1n02x5               g038(.a(new_n131), .b(new_n132), .out0(new_n134));
  aoib12aa1n02x5               g039(.a(new_n134), .b(new_n129), .c(new_n127), .out0(new_n135));
  aoi012aa1n02x5               g040(.a(new_n135), .b(new_n129), .c(new_n133), .o1(\s[11] ));
  aoi012aa1n02x5               g041(.a(new_n132), .b(new_n129), .c(new_n133), .o1(new_n137));
  nor042aa1n06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand42aa1d28x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  nona22aa1n09x5               g045(.a(new_n139), .b(new_n138), .c(new_n132), .out0(new_n141));
  tech160nm_fiao0012aa1n02p5x5 g046(.a(new_n141), .b(new_n129), .c(new_n133), .o(new_n142));
  oai012aa1n02x5               g047(.a(new_n142), .b(new_n137), .c(new_n140), .o1(\s[12] ));
  nano23aa1d15x5               g048(.a(new_n138), .b(new_n132), .c(new_n139), .d(new_n131), .out0(new_n144));
  nanb02aa1n02x5               g049(.a(new_n98), .b(new_n99), .out0(new_n145));
  nona22aa1d18x5               g050(.a(new_n144), .b(new_n97), .c(new_n145), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  oab012aa1n09x5               g052(.a(new_n127), .b(new_n126), .c(new_n98), .out0(new_n148));
  aoi022aa1d24x5               g053(.a(new_n144), .b(new_n148), .c(new_n141), .d(new_n139), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  xnrc02aa1n12x5               g055(.a(\b[12] ), .b(\a[13] ), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n150), .c(new_n124), .d(new_n147), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n152), .b(new_n150), .c(new_n124), .d(new_n147), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(\s[13] ));
  nor042aa1d18x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  inv040aa1n08x5               g061(.a(new_n156), .o1(new_n157));
  tech160nm_fixnrc02aa1n02p5x5 g062(.a(\b[13] ), .b(\a[14] ), .out0(new_n158));
  xobna2aa1n03x5               g063(.a(new_n158), .b(new_n153), .c(new_n157), .out0(\s[14] ));
  norp02aa1n02x5               g064(.a(new_n158), .b(new_n151), .o1(new_n160));
  aoai13aa1n06x5               g065(.a(new_n160), .b(new_n150), .c(new_n124), .d(new_n147), .o1(new_n161));
  oaoi03aa1n12x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nor042aa1n03x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n161), .c(new_n163), .out0(\s[15] ));
  aobi12aa1n06x5               g072(.a(new_n166), .b(new_n161), .c(new_n163), .out0(new_n168));
  nor042aa1n03x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nand42aa1n06x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nanb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(new_n171));
  oai012aa1n02x5               g076(.a(new_n171), .b(new_n168), .c(new_n164), .o1(new_n172));
  norb03aa1n03x5               g077(.a(new_n170), .b(new_n164), .c(new_n169), .out0(new_n173));
  oaib12aa1n02x5               g078(.a(new_n172), .b(new_n168), .c(new_n173), .out0(\s[16] ));
  nano23aa1d15x5               g079(.a(new_n164), .b(new_n169), .c(new_n170), .d(new_n165), .out0(new_n175));
  nona22aa1n09x5               g080(.a(new_n175), .b(new_n158), .c(new_n151), .out0(new_n176));
  nor042aa1n06x5               g081(.a(new_n176), .b(new_n146), .o1(new_n177));
  nanp02aa1n06x5               g082(.a(new_n124), .b(new_n177), .o1(new_n178));
  aboi22aa1n12x5               g083(.a(new_n173), .b(new_n170), .c(new_n175), .d(new_n162), .out0(new_n179));
  oai012aa1d24x5               g084(.a(new_n179), .b(new_n149), .c(new_n176), .o1(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  xorc02aa1n12x5               g086(.a(\a[17] ), .b(\b[16] ), .out0(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n178), .c(new_n181), .out0(\s[17] ));
  nor042aa1d18x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  inv040aa1n08x5               g089(.a(new_n184), .o1(new_n185));
  aoai13aa1n02x5               g090(.a(new_n182), .b(new_n180), .c(new_n124), .d(new_n177), .o1(new_n186));
  xnrc02aa1n12x5               g091(.a(\b[17] ), .b(\a[18] ), .out0(new_n187));
  xobna2aa1n03x5               g092(.a(new_n187), .b(new_n186), .c(new_n185), .out0(\s[18] ));
  norb02aa1n02x5               g093(.a(new_n182), .b(new_n187), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n180), .c(new_n124), .d(new_n177), .o1(new_n190));
  oaoi03aa1n12x5               g095(.a(\a[18] ), .b(\b[17] ), .c(new_n185), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  nor002aa1n12x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nand02aa1d16x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  norb02aa1n06x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n190), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aobi12aa1n06x5               g102(.a(new_n195), .b(new_n190), .c(new_n192), .out0(new_n198));
  nor042aa1n06x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1d28x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1n03x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  oabi12aa1n02x5               g106(.a(new_n201), .b(new_n198), .c(new_n193), .out0(new_n202));
  norb03aa1n02x5               g107(.a(new_n200), .b(new_n193), .c(new_n199), .out0(new_n203));
  oaib12aa1n02x5               g108(.a(new_n202), .b(new_n198), .c(new_n203), .out0(\s[20] ));
  nano23aa1d15x5               g109(.a(new_n193), .b(new_n199), .c(new_n200), .d(new_n194), .out0(new_n205));
  nanb03aa1d18x5               g110(.a(new_n187), .b(new_n205), .c(new_n182), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n180), .c(new_n124), .d(new_n177), .o1(new_n208));
  nor002aa1n02x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  aoi112aa1n06x5               g114(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n210));
  oai112aa1n06x5               g115(.a(new_n195), .b(new_n201), .c(new_n210), .d(new_n209), .o1(new_n211));
  oaib12aa1n02x5               g116(.a(new_n211), .b(new_n203), .c(new_n200), .out0(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  tech160nm_fixorc02aa1n04x5   g118(.a(\a[21] ), .b(\b[20] ), .out0(new_n214));
  xnbna2aa1n03x5               g119(.a(new_n214), .b(new_n208), .c(new_n213), .out0(\s[21] ));
  aobi12aa1n06x5               g120(.a(new_n214), .b(new_n208), .c(new_n213), .out0(new_n216));
  nor042aa1n02x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  xnrc02aa1n02x5               g122(.a(\b[21] ), .b(\a[22] ), .out0(new_n218));
  tech160nm_fioai012aa1n05x5   g123(.a(new_n218), .b(new_n216), .c(new_n217), .o1(new_n219));
  norp02aa1n02x5               g124(.a(new_n218), .b(new_n217), .o1(new_n220));
  oaib12aa1n02x5               g125(.a(new_n219), .b(new_n216), .c(new_n220), .out0(\s[22] ));
  inv000aa1d42x5               g126(.a(\a[21] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\a[22] ), .o1(new_n223));
  xroi22aa1d04x5               g128(.a(new_n222), .b(\b[20] ), .c(new_n223), .d(\b[21] ), .out0(new_n224));
  nanp03aa1n02x5               g129(.a(new_n189), .b(new_n205), .c(new_n224), .o1(new_n225));
  tech160nm_fiao0012aa1n02p5x5 g130(.a(new_n225), .b(new_n178), .c(new_n181), .o(new_n226));
  oa0012aa1n06x5               g131(.a(new_n200), .b(new_n199), .c(new_n193), .o(new_n227));
  inv040aa1n02x5               g132(.a(new_n227), .o1(new_n228));
  nanb02aa1n03x5               g133(.a(new_n218), .b(new_n214), .out0(new_n229));
  inv000aa1d42x5               g134(.a(\b[21] ), .o1(new_n230));
  oaoi03aa1n09x5               g135(.a(new_n223), .b(new_n230), .c(new_n217), .o1(new_n231));
  aoai13aa1n12x5               g136(.a(new_n231), .b(new_n229), .c(new_n228), .d(new_n211), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n225), .c(new_n178), .d(new_n181), .o1(new_n234));
  xorc02aa1n12x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n224), .b(new_n227), .c(new_n205), .d(new_n191), .o1(new_n236));
  nano22aa1n02x4               g141(.a(new_n235), .b(new_n236), .c(new_n231), .out0(new_n237));
  aoi022aa1n02x5               g142(.a(new_n226), .b(new_n237), .c(new_n234), .d(new_n235), .o1(\s[23] ));
  nor002aa1n02x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[23] ), .b(\a[24] ), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n239), .c(new_n234), .d(new_n235), .o1(new_n241));
  norp02aa1n02x5               g146(.a(new_n240), .b(new_n239), .o1(new_n242));
  aob012aa1n03x5               g147(.a(new_n242), .b(new_n234), .c(new_n235), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n241), .b(new_n243), .o1(\s[24] ));
  norb02aa1n06x4               g149(.a(new_n235), .b(new_n240), .out0(new_n245));
  nanb03aa1n02x5               g150(.a(new_n206), .b(new_n245), .c(new_n224), .out0(new_n246));
  inv030aa1n02x5               g151(.a(new_n245), .o1(new_n247));
  inv000aa1d42x5               g152(.a(\a[24] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(\b[23] ), .o1(new_n249));
  oao003aa1n02x5               g154(.a(new_n248), .b(new_n249), .c(new_n239), .carry(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n12x5               g156(.a(new_n251), .b(new_n247), .c(new_n236), .d(new_n231), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n246), .c(new_n178), .d(new_n181), .o1(new_n254));
  xorb03aa1n02x5               g159(.a(new_n254), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g160(.a(\b[24] ), .b(\a[25] ), .o1(new_n256));
  tech160nm_fixorc02aa1n03p5x5 g161(.a(\a[25] ), .b(\b[24] ), .out0(new_n257));
  xnrc02aa1n02x5               g162(.a(\b[25] ), .b(\a[26] ), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n256), .c(new_n254), .d(new_n257), .o1(new_n259));
  oabi12aa1n02x5               g164(.a(new_n258), .b(\a[25] ), .c(\b[24] ), .out0(new_n260));
  ao0012aa1n03x7               g165(.a(new_n260), .b(new_n254), .c(new_n257), .o(new_n261));
  nanp02aa1n03x5               g166(.a(new_n261), .b(new_n259), .o1(\s[26] ));
  norb02aa1n02x5               g167(.a(new_n257), .b(new_n258), .out0(new_n263));
  nano23aa1n06x5               g168(.a(new_n247), .b(new_n206), .c(new_n263), .d(new_n224), .out0(new_n264));
  aoai13aa1n12x5               g169(.a(new_n264), .b(new_n180), .c(new_n124), .d(new_n177), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n263), .b(new_n250), .c(new_n232), .d(new_n245), .o1(new_n266));
  aob012aa1n02x5               g171(.a(new_n260), .b(\b[25] ), .c(\a[26] ), .out0(new_n267));
  nand23aa1n06x5               g172(.a(new_n265), .b(new_n266), .c(new_n267), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[27] ), .b(\b[26] ), .out0(new_n271));
  xnrc02aa1n12x5               g176(.a(\b[27] ), .b(\a[28] ), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n270), .c(new_n268), .d(new_n271), .o1(new_n273));
  aobi12aa1n06x5               g178(.a(new_n267), .b(new_n252), .c(new_n263), .out0(new_n274));
  inv000aa1d42x5               g179(.a(new_n271), .o1(new_n275));
  nor042aa1n03x5               g180(.a(new_n272), .b(new_n270), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .d(new_n265), .o1(new_n277));
  nanp02aa1n03x5               g182(.a(new_n273), .b(new_n277), .o1(\s[28] ));
  norb02aa1n03x5               g183(.a(new_n271), .b(new_n272), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  xnrc02aa1n12x5               g185(.a(\b[28] ), .b(\a[29] ), .out0(new_n281));
  tech160nm_fiaoi012aa1n05x5   g186(.a(new_n276), .b(\a[28] ), .c(\b[27] ), .o1(new_n282));
  norp02aa1n02x5               g187(.a(new_n282), .b(new_n281), .o1(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n280), .c(new_n274), .d(new_n265), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n281), .b(new_n282), .c(new_n268), .d(new_n279), .o1(new_n285));
  nanp02aa1n03x5               g190(.a(new_n285), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g191(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g192(.a(new_n271), .b(new_n281), .c(new_n272), .out0(new_n288));
  nanp02aa1n03x5               g193(.a(new_n268), .b(new_n288), .o1(new_n289));
  inv000aa1d42x5               g194(.a(\b[28] ), .o1(new_n290));
  oaib12aa1n06x5               g195(.a(new_n282), .b(new_n290), .c(\a[29] ), .out0(new_n291));
  oa0012aa1n02x5               g196(.a(new_n291), .b(\b[28] ), .c(\a[29] ), .o(new_n292));
  xorc02aa1n02x5               g197(.a(\a[30] ), .b(\b[29] ), .out0(new_n293));
  inv000aa1n02x5               g198(.a(new_n288), .o1(new_n294));
  oai112aa1n06x5               g199(.a(new_n291), .b(new_n293), .c(\b[28] ), .d(\a[29] ), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n294), .c(new_n274), .d(new_n265), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n293), .c(new_n289), .d(new_n292), .o1(\s[30] ));
  nano23aa1d12x5               g203(.a(new_n281), .b(new_n272), .c(new_n293), .d(new_n271), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(\a[30] ), .o1(new_n301));
  inv000aa1d42x5               g206(.a(\b[29] ), .o1(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[30] ), .b(\a[31] ), .out0(new_n303));
  oaoi13aa1n02x5               g208(.a(new_n303), .b(new_n295), .c(new_n301), .d(new_n302), .o1(new_n304));
  aoai13aa1n02x5               g209(.a(new_n304), .b(new_n300), .c(new_n274), .d(new_n265), .o1(new_n305));
  oa0012aa1n02x5               g210(.a(new_n295), .b(new_n302), .c(new_n301), .o(new_n306));
  aoai13aa1n03x5               g211(.a(new_n303), .b(new_n306), .c(new_n268), .d(new_n299), .o1(new_n307));
  nanp02aa1n03x5               g212(.a(new_n307), .b(new_n305), .o1(\s[31] ));
  norb02aa1n02x5               g213(.a(new_n105), .b(new_n104), .out0(new_n309));
  xobna2aa1n03x5               g214(.a(new_n309), .b(new_n109), .c(new_n103), .out0(\s[3] ));
  inv000aa1d42x5               g215(.a(new_n104), .o1(new_n311));
  oai112aa1n02x5               g216(.a(new_n309), .b(new_n103), .c(new_n107), .d(new_n108), .o1(new_n312));
  xnbna2aa1n03x5               g217(.a(new_n102), .b(new_n312), .c(new_n311), .out0(\s[4] ));
  xnbna2aa1n03x5               g218(.a(new_n118), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  aob012aa1n02x5               g219(.a(new_n118), .b(new_n110), .c(new_n111), .out0(new_n315));
  xnbna2aa1n03x5               g220(.a(new_n117), .b(new_n315), .c(new_n120), .out0(\s[6] ));
  nanb02aa1n02x5               g221(.a(new_n114), .b(new_n115), .out0(new_n317));
  nanp02aa1n02x5               g222(.a(\b[5] ), .b(\a[6] ), .o1(new_n318));
  nanp03aa1n02x5               g223(.a(new_n315), .b(new_n117), .c(new_n120), .o1(new_n319));
  xnbna2aa1n03x5               g224(.a(new_n317), .b(new_n319), .c(new_n318), .out0(\s[7] ));
  norb02aa1n02x5               g225(.a(new_n113), .b(new_n112), .out0(new_n321));
  nano22aa1n02x4               g226(.a(new_n317), .b(new_n319), .c(new_n318), .out0(new_n322));
  aoi013aa1n02x4               g227(.a(new_n114), .b(new_n319), .c(new_n318), .d(new_n115), .o1(new_n323));
  oai022aa1n02x5               g228(.a(new_n321), .b(new_n323), .c(new_n322), .d(new_n122), .o1(\s[8] ));
  xorb03aa1n02x5               g229(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


