// Benchmark "adder" written by ABC on Wed Jul 17 21:07:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n315, new_n316, new_n317, new_n319,
    new_n320, new_n322, new_n323, new_n324, new_n325;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  tech160nm_fixnrc02aa1n04x5   g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  nand22aa1n04x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand42aa1n10x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor042aa1d18x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai012aa1n12x5               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  orn002aa1n24x5               g008(.a(\a[4] ), .b(\b[3] ), .o(new_n104));
  nand42aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  oai112aa1n06x5               g010(.a(new_n104), .b(new_n105), .c(\b[2] ), .d(\a[3] ), .o1(new_n106));
  oabi12aa1n18x5               g011(.a(new_n106), .b(new_n99), .c(new_n103), .out0(new_n107));
  inv020aa1d28x5               g012(.a(\a[5] ), .o1(new_n108));
  inv040aa1d32x5               g013(.a(\b[4] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  inv040aa1n08x5               g015(.a(new_n110), .o1(new_n111));
  oai122aa1n06x5               g016(.a(new_n111), .b(\a[6] ), .c(\b[5] ), .d(new_n108), .e(new_n109), .o1(new_n112));
  aoi022aa1n06x5               g017(.a(new_n109), .b(new_n108), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  nor022aa1n16x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nanb02aa1n03x5               g020(.a(new_n114), .b(new_n115), .out0(new_n116));
  aoi022aa1d24x5               g021(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n117));
  nano23aa1n06x5               g022(.a(new_n112), .b(new_n116), .c(new_n113), .d(new_n117), .out0(new_n118));
  oaoi03aa1n02x5               g023(.a(\a[8] ), .b(\b[7] ), .c(new_n111), .o1(new_n119));
  nor022aa1n08x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  and002aa1n03x5               g025(.a(\b[5] ), .b(\a[6] ), .o(new_n121));
  aoi112aa1n06x5               g026(.a(new_n121), .b(new_n120), .c(new_n108), .d(new_n109), .o1(new_n122));
  nona23aa1n03x5               g027(.a(new_n117), .b(new_n115), .c(new_n110), .d(new_n114), .out0(new_n123));
  oabi12aa1n06x5               g028(.a(new_n119), .b(new_n123), .c(new_n122), .out0(new_n124));
  tech160nm_fiao0012aa1n05x5   g029(.a(new_n124), .b(new_n118), .c(new_n107), .o(new_n125));
  nand42aa1d28x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  nand43aa1n02x5               g031(.a(new_n125), .b(new_n98), .c(new_n126), .o1(new_n127));
  nor042aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  oai022aa1d18x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  nanb03aa1n02x5               g036(.a(new_n131), .b(new_n127), .c(new_n129), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n130), .c(new_n98), .d(new_n127), .o1(\s[10] ));
  nano23aa1d15x5               g038(.a(new_n97), .b(new_n128), .c(new_n129), .d(new_n126), .out0(new_n134));
  aoi022aa1n09x5               g039(.a(new_n125), .b(new_n134), .c(new_n129), .d(new_n131), .o1(new_n135));
  nor002aa1n20x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n136), .o1(new_n137));
  nand02aa1d16x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n135), .b(new_n138), .c(new_n137), .out0(\s[11] ));
  norb02aa1n02x5               g044(.a(new_n138), .b(new_n136), .out0(new_n140));
  nanb02aa1n03x5               g045(.a(new_n135), .b(new_n140), .out0(new_n141));
  nor042aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n24x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  norb03aa1n02x5               g049(.a(new_n143), .b(new_n136), .c(new_n142), .out0(new_n145));
  oaib12aa1n03x5               g050(.a(new_n145), .b(new_n135), .c(new_n140), .out0(new_n146));
  aoai13aa1n03x5               g051(.a(new_n146), .b(new_n144), .c(new_n141), .d(new_n137), .o1(\s[12] ));
  nano23aa1d15x5               g052(.a(new_n136), .b(new_n142), .c(new_n143), .d(new_n138), .out0(new_n148));
  nand22aa1n12x5               g053(.a(new_n148), .b(new_n134), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n124), .c(new_n118), .d(new_n107), .o1(new_n151));
  oai022aa1n04x5               g056(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n152));
  aoi022aa1d24x5               g057(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  aoai13aa1n06x5               g058(.a(new_n143), .b(new_n152), .c(new_n131), .d(new_n153), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(new_n151), .b(new_n154), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nanp02aa1n12x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanp03aa1n03x5               g064(.a(new_n155), .b(new_n158), .c(new_n159), .o1(new_n160));
  nor002aa1n08x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand02aa1n06x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  nona23aa1n02x4               g068(.a(new_n160), .b(new_n162), .c(new_n161), .d(new_n157), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n163), .c(new_n158), .d(new_n160), .o1(\s[14] ));
  nona23aa1n09x5               g070(.a(new_n162), .b(new_n159), .c(new_n157), .d(new_n161), .out0(new_n166));
  oai012aa1n02x5               g071(.a(new_n162), .b(new_n161), .c(new_n157), .o1(new_n167));
  tech160nm_fioai012aa1n04x5   g072(.a(new_n167), .b(new_n154), .c(new_n166), .o1(new_n168));
  oabi12aa1n06x5               g073(.a(new_n168), .b(new_n151), .c(new_n166), .out0(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n06x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand42aa1n06x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  nor042aa1n04x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1n08x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  norb02aa1n02x5               g081(.a(new_n172), .b(new_n171), .out0(new_n177));
  oaih22aa1n04x5               g082(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n178));
  aoi122aa1n03x5               g083(.a(new_n178), .b(\b[15] ), .c(\a[16] ), .d(new_n169), .e(new_n177), .o1(new_n179));
  oabi12aa1n03x5               g084(.a(new_n179), .b(new_n173), .c(new_n176), .out0(\s[16] ));
  nano23aa1n03x7               g085(.a(new_n157), .b(new_n161), .c(new_n162), .d(new_n159), .out0(new_n181));
  nano23aa1d12x5               g086(.a(new_n171), .b(new_n174), .c(new_n175), .d(new_n172), .out0(new_n182));
  nano22aa1d15x5               g087(.a(new_n149), .b(new_n181), .c(new_n182), .out0(new_n183));
  aoai13aa1n12x5               g088(.a(new_n183), .b(new_n124), .c(new_n107), .d(new_n118), .o1(new_n184));
  aoi022aa1n12x5               g089(.a(new_n168), .b(new_n182), .c(new_n175), .d(new_n178), .o1(new_n185));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n184), .out0(\s[17] ));
  nor002aa1n16x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  nanp02aa1n12x5               g094(.a(new_n185), .b(new_n184), .o1(new_n190));
  nanp02aa1n06x5               g095(.a(new_n190), .b(new_n186), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[18] ), .b(\b[17] ), .out0(new_n192));
  nand42aa1n16x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  oai022aa1d18x5               g098(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n194));
  nanb03aa1n03x5               g099(.a(new_n194), .b(new_n191), .c(new_n193), .out0(new_n195));
  aoai13aa1n03x5               g100(.a(new_n195), .b(new_n192), .c(new_n189), .d(new_n191), .o1(\s[18] ));
  nand42aa1d28x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nor042aa1n04x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nano23aa1d15x5               g103(.a(new_n188), .b(new_n198), .c(new_n193), .d(new_n197), .out0(new_n199));
  oaoi03aa1n02x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n200));
  xorc02aa1n12x5               g105(.a(\a[19] ), .b(\b[18] ), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n202));
  aoi112aa1n02x5               g107(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n203));
  norb02aa1n03x4               g108(.a(new_n202), .b(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[18] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  xorc02aa1n12x5               g113(.a(\a[20] ), .b(\b[19] ), .out0(new_n209));
  nand02aa1n08x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  oai022aa1n02x7               g116(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n212));
  nona22aa1n03x5               g117(.a(new_n202), .b(new_n211), .c(new_n212), .out0(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n208), .d(new_n202), .o1(\s[20] ));
  nand23aa1n06x5               g119(.a(new_n199), .b(new_n201), .c(new_n209), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  oai112aa1n03x5               g121(.a(new_n194), .b(new_n193), .c(new_n207), .d(new_n206), .o1(new_n217));
  aoib12aa1n02x5               g122(.a(new_n211), .b(new_n217), .c(new_n212), .out0(new_n218));
  orn002aa1n24x5               g123(.a(\a[21] ), .b(\b[20] ), .o(new_n219));
  nand22aa1n12x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  nanp02aa1n12x5               g125(.a(new_n219), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n218), .c(new_n190), .d(new_n216), .o1(new_n223));
  aoi112aa1n02x7               g128(.a(new_n222), .b(new_n218), .c(new_n190), .d(new_n216), .o1(new_n224));
  norb02aa1n03x4               g129(.a(new_n223), .b(new_n224), .out0(\s[21] ));
  xnrc02aa1n12x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  and002aa1n02x5               g132(.a(\b[21] ), .b(\a[22] ), .o(new_n228));
  oai022aa1n02x5               g133(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n229));
  nona22aa1n03x5               g134(.a(new_n223), .b(new_n228), .c(new_n229), .out0(new_n230));
  aoai13aa1n03x5               g135(.a(new_n230), .b(new_n227), .c(new_n219), .d(new_n223), .o1(\s[22] ));
  nor002aa1n02x5               g136(.a(new_n226), .b(new_n221), .o1(new_n232));
  norb02aa1n09x5               g137(.a(new_n232), .b(new_n215), .out0(new_n233));
  nanb02aa1n06x5               g138(.a(new_n212), .b(new_n217), .out0(new_n234));
  nano32aa1n03x7               g139(.a(new_n226), .b(new_n219), .c(new_n220), .d(new_n210), .out0(new_n235));
  nanp02aa1n02x5               g140(.a(new_n234), .b(new_n235), .o1(new_n236));
  oaib12aa1n02x5               g141(.a(new_n236), .b(new_n228), .c(new_n229), .out0(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n237), .c(new_n190), .d(new_n233), .o1(new_n239));
  oaoi03aa1n03x5               g144(.a(\a[22] ), .b(\b[21] ), .c(new_n219), .o1(new_n240));
  nona22aa1n02x4               g145(.a(new_n236), .b(new_n240), .c(new_n238), .out0(new_n241));
  aoi012aa1n02x5               g146(.a(new_n241), .b(new_n190), .c(new_n233), .o1(new_n242));
  norb02aa1n03x4               g147(.a(new_n239), .b(new_n242), .out0(\s[23] ));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  tech160nm_fixorc02aa1n02p5x5 g150(.a(\a[24] ), .b(\b[23] ), .out0(new_n246));
  and002aa1n02x5               g151(.a(\b[23] ), .b(\a[24] ), .o(new_n247));
  oai022aa1n02x5               g152(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n248));
  nona22aa1n03x5               g153(.a(new_n239), .b(new_n247), .c(new_n248), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n246), .c(new_n245), .d(new_n239), .o1(\s[24] ));
  nano32aa1n02x5               g155(.a(new_n215), .b(new_n246), .c(new_n232), .d(new_n238), .out0(new_n251));
  and002aa1n06x5               g156(.a(new_n246), .b(new_n238), .o(new_n252));
  aoai13aa1n04x5               g157(.a(new_n252), .b(new_n240), .c(new_n234), .d(new_n235), .o1(new_n253));
  aob012aa1n02x5               g158(.a(new_n248), .b(\b[23] ), .c(\a[24] ), .out0(new_n254));
  nanp02aa1n02x5               g159(.a(new_n253), .b(new_n254), .o1(new_n255));
  xnrc02aa1n12x5               g160(.a(\b[24] ), .b(\a[25] ), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n255), .c(new_n190), .d(new_n251), .o1(new_n258));
  aoi112aa1n02x5               g163(.a(new_n257), .b(new_n255), .c(new_n190), .d(new_n251), .o1(new_n259));
  norb02aa1n03x4               g164(.a(new_n258), .b(new_n259), .out0(\s[25] ));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  and002aa1n02x5               g168(.a(\b[25] ), .b(\a[26] ), .o(new_n264));
  oai022aa1n02x5               g169(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n265));
  nona22aa1n03x5               g170(.a(new_n258), .b(new_n264), .c(new_n265), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n266), .b(new_n263), .c(new_n262), .d(new_n258), .o1(\s[26] ));
  norb02aa1n09x5               g172(.a(new_n263), .b(new_n256), .out0(new_n268));
  nand23aa1n02x5               g173(.a(new_n233), .b(new_n252), .c(new_n268), .o1(new_n269));
  inv040aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n268), .o1(new_n271));
  aob012aa1n02x5               g176(.a(new_n265), .b(\b[25] ), .c(\a[26] ), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n271), .c(new_n253), .d(new_n254), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n190), .d(new_n270), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(new_n274), .b(new_n273), .c(new_n190), .d(new_n270), .o1(new_n276));
  norb02aa1n03x4               g181(.a(new_n275), .b(new_n276), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  xorc02aa1n02x5               g184(.a(\a[28] ), .b(\b[27] ), .out0(new_n280));
  oai022aa1d24x5               g185(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n281));
  aoi012aa1n02x5               g186(.a(new_n281), .b(\a[28] ), .c(\b[27] ), .o1(new_n282));
  tech160nm_finand02aa1n05x5   g187(.a(new_n275), .b(new_n282), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n280), .c(new_n279), .d(new_n275), .o1(\s[28] ));
  xorc02aa1n02x5               g189(.a(\a[29] ), .b(\b[28] ), .out0(new_n285));
  and002aa1n02x5               g190(.a(new_n280), .b(new_n274), .o(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n273), .c(new_n190), .d(new_n270), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[27] ), .o1(new_n288));
  oaib12aa1n18x5               g193(.a(new_n281), .b(new_n288), .c(\a[28] ), .out0(new_n289));
  nanp03aa1n03x5               g194(.a(new_n287), .b(new_n289), .c(new_n285), .o1(new_n290));
  tech160nm_fiaoi012aa1n04x5   g195(.a(new_n269), .b(new_n185), .c(new_n184), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n289), .o1(new_n292));
  oaoi13aa1n02x5               g197(.a(new_n292), .b(new_n286), .c(new_n291), .d(new_n273), .o1(new_n293));
  oai012aa1n03x5               g198(.a(new_n290), .b(new_n293), .c(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g200(.a(new_n274), .b(new_n285), .c(new_n280), .o(new_n296));
  tech160nm_fioaoi03aa1n03p5x5 g201(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .o1(new_n297));
  oaoi13aa1n02x7               g202(.a(new_n297), .b(new_n296), .c(new_n291), .d(new_n273), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n296), .b(new_n273), .c(new_n190), .d(new_n270), .o1(new_n300));
  norb02aa1n03x5               g205(.a(new_n299), .b(new_n297), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n300), .b(new_n301), .o1(new_n302));
  oai012aa1n03x5               g207(.a(new_n302), .b(new_n298), .c(new_n299), .o1(\s[30] ));
  and003aa1n02x5               g208(.a(new_n286), .b(new_n299), .c(new_n285), .o(new_n304));
  tech160nm_fiaoi012aa1n03p5x5 g209(.a(new_n301), .b(\a[30] ), .c(\b[29] ), .o1(new_n305));
  oaoi13aa1n02x7               g210(.a(new_n305), .b(new_n304), .c(new_n291), .d(new_n273), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[31] ), .b(\b[30] ), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n304), .b(new_n273), .c(new_n190), .d(new_n270), .o1(new_n308));
  norb02aa1n02x5               g213(.a(new_n307), .b(new_n305), .out0(new_n309));
  nanp02aa1n03x5               g214(.a(new_n308), .b(new_n309), .o1(new_n310));
  oai012aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n307), .o1(\s[31] ));
  xnrb03aa1n02x5               g216(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oao003aa1n02x5               g217(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .carry(new_n313));
  aoai13aa1n02x5               g218(.a(new_n107), .b(new_n313), .c(new_n105), .d(new_n104), .o1(\s[4] ));
  nanp02aa1n02x5               g219(.a(\b[4] ), .b(\a[5] ), .o1(new_n315));
  nanp02aa1n02x5               g220(.a(new_n109), .b(new_n108), .o1(new_n316));
  aoi022aa1n02x5               g221(.a(new_n107), .b(new_n105), .c(new_n316), .d(new_n315), .o1(new_n317));
  aoi013aa1n02x4               g222(.a(new_n317), .b(new_n113), .c(new_n315), .d(new_n107), .o1(\s[5] ));
  norp02aa1n02x5               g223(.a(new_n121), .b(new_n120), .o1(new_n319));
  nanp03aa1n03x5               g224(.a(new_n107), .b(new_n315), .c(new_n113), .o1(new_n320));
  xnbna2aa1n03x5               g225(.a(new_n319), .b(new_n320), .c(new_n316), .out0(\s[6] ));
  nanp02aa1n02x5               g226(.a(new_n320), .b(new_n122), .o1(new_n322));
  nanp03aa1n03x5               g227(.a(new_n322), .b(new_n111), .c(new_n117), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[7] ), .b(\b[6] ), .out0(new_n324));
  aoib12aa1n02x5               g229(.a(new_n324), .b(new_n322), .c(new_n121), .out0(new_n325));
  norb02aa1n02x5               g230(.a(new_n323), .b(new_n325), .out0(\s[7] ));
  xobna2aa1n03x5               g231(.a(new_n116), .b(new_n323), .c(new_n111), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


