// Benchmark "adder" written by ABC on Thu Jul 18 11:49:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n325, new_n326, new_n327, new_n329, new_n330, new_n331,
    new_n333, new_n334, new_n335, new_n337, new_n338, new_n340, new_n341,
    new_n342, new_n343, new_n345, new_n346, new_n348, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n16x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n16x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norb03aa1d15x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  inv040aa1d32x5               g007(.a(\a[3] ), .o1(new_n103));
  aoi022aa1n12x5               g008(.a(\b[2] ), .b(\a[3] ), .c(\a[2] ), .d(\b[1] ), .o1(new_n104));
  oaib12aa1n06x5               g009(.a(new_n104), .b(\b[2] ), .c(new_n103), .out0(new_n105));
  inv000aa1d42x5               g010(.a(\a[4] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[3] ), .o1(new_n107));
  aboi22aa1n06x5               g012(.a(\b[2] ), .b(new_n103), .c(new_n107), .d(new_n106), .out0(new_n108));
  oai012aa1n18x5               g013(.a(new_n108), .b(new_n102), .c(new_n105), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  inv040aa1n02x5               g015(.a(new_n110), .o1(new_n111));
  nanp02aa1n12x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  oai112aa1n03x5               g017(.a(new_n111), .b(new_n112), .c(new_n107), .d(new_n106), .o1(new_n113));
  tech160nm_fixnrc02aa1n04x5   g018(.a(\b[5] ), .b(\a[6] ), .out0(new_n114));
  nor002aa1d32x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nor022aa1n08x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand02aa1d28x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nona23aa1n09x5               g023(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n119));
  nor043aa1n04x5               g024(.a(new_n119), .b(new_n114), .c(new_n113), .o1(new_n120));
  nano22aa1n02x4               g025(.a(new_n110), .b(new_n112), .c(new_n118), .out0(new_n121));
  nanp02aa1n02x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  oaih22aa1d12x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  oai112aa1n03x5               g028(.a(new_n123), .b(new_n122), .c(\b[7] ), .d(\a[8] ), .o1(new_n124));
  aoi012aa1n02x5               g029(.a(new_n117), .b(new_n110), .c(new_n118), .o1(new_n125));
  oaib12aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n121), .out0(new_n126));
  nand02aa1n08x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n97), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n126), .c(new_n120), .d(new_n109), .o1(new_n129));
  nor002aa1d32x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand02aa1n16x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  nand42aa1n02x5               g038(.a(new_n129), .b(new_n98), .o1(new_n134));
  oaoi03aa1n02x5               g039(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n135));
  nor042aa1d18x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand02aa1d28x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aoai13aa1n06x5               g043(.a(new_n138), .b(new_n135), .c(new_n134), .d(new_n132), .o1(new_n139));
  aoi112aa1n02x5               g044(.a(new_n138), .b(new_n135), .c(new_n134), .d(new_n132), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(\s[11] ));
  nor002aa1d32x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d28x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  norp02aa1n02x5               g049(.a(new_n144), .b(new_n136), .o1(new_n145));
  tech160nm_fioai012aa1n03p5x5 g050(.a(new_n139), .b(\b[10] ), .c(\a[11] ), .o1(new_n146));
  aoi022aa1n02x5               g051(.a(new_n146), .b(new_n144), .c(new_n139), .d(new_n145), .o1(\s[12] ));
  nano23aa1n09x5               g052(.a(new_n136), .b(new_n142), .c(new_n143), .d(new_n137), .out0(new_n148));
  nano23aa1n09x5               g053(.a(new_n97), .b(new_n130), .c(new_n131), .d(new_n127), .out0(new_n149));
  nand22aa1n09x5               g054(.a(new_n149), .b(new_n148), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n126), .c(new_n120), .d(new_n109), .o1(new_n152));
  nanb03aa1n03x5               g057(.a(new_n142), .b(new_n143), .c(new_n137), .out0(new_n153));
  inv030aa1n03x5               g058(.a(new_n136), .o1(new_n154));
  oai112aa1n06x5               g059(.a(new_n154), .b(new_n131), .c(new_n130), .d(new_n97), .o1(new_n155));
  norp02aa1n02x5               g060(.a(new_n155), .b(new_n153), .o1(new_n156));
  aoi012aa1d24x5               g061(.a(new_n142), .b(new_n136), .c(new_n143), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nona22aa1n03x5               g063(.a(new_n152), .b(new_n156), .c(new_n158), .out0(new_n159));
  nor042aa1d18x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand02aa1n04x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  norp03aa1n02x5               g067(.a(new_n156), .b(new_n158), .c(new_n162), .o1(new_n163));
  aoi022aa1n02x5               g068(.a(new_n159), .b(new_n162), .c(new_n152), .d(new_n163), .o1(\s[13] ));
  inv040aa1n02x5               g069(.a(new_n160), .o1(new_n165));
  nona32aa1n02x4               g070(.a(new_n109), .b(new_n119), .c(new_n114), .d(new_n113), .out0(new_n166));
  nanb02aa1n02x5               g071(.a(new_n126), .b(new_n166), .out0(new_n167));
  oai012aa1n06x5               g072(.a(new_n157), .b(new_n155), .c(new_n153), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n162), .b(new_n168), .c(new_n167), .d(new_n151), .o1(new_n169));
  nor042aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand02aa1n04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n169), .c(new_n165), .out0(\s[14] ));
  nano23aa1d15x5               g078(.a(new_n160), .b(new_n170), .c(new_n171), .d(new_n161), .out0(new_n174));
  tech160nm_fioaoi03aa1n02p5x5 g079(.a(\a[14] ), .b(\b[13] ), .c(new_n165), .o1(new_n175));
  nor042aa1n04x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nand42aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n175), .c(new_n159), .d(new_n174), .o1(new_n179));
  aoi112aa1n02x5               g084(.a(new_n178), .b(new_n175), .c(new_n159), .d(new_n174), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(\s[15] ));
  nor042aa1n04x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand02aa1d08x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  aoib12aa1n02x5               g089(.a(new_n176), .b(new_n183), .c(new_n182), .out0(new_n185));
  tech160nm_fioai012aa1n03p5x5 g090(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(new_n186), .b(new_n184), .c(new_n179), .d(new_n185), .o1(\s[16] ));
  nano23aa1n06x5               g092(.a(new_n176), .b(new_n182), .c(new_n183), .d(new_n177), .out0(new_n188));
  aoai13aa1n09x5               g093(.a(new_n188), .b(new_n175), .c(new_n168), .d(new_n174), .o1(new_n189));
  nano22aa1n12x5               g094(.a(new_n150), .b(new_n174), .c(new_n188), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n126), .c(new_n109), .d(new_n120), .o1(new_n191));
  aoi012aa1d18x5               g096(.a(new_n182), .b(new_n176), .c(new_n183), .o1(new_n192));
  nand23aa1d12x5               g097(.a(new_n191), .b(new_n189), .c(new_n192), .o1(new_n193));
  xorc02aa1n12x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  nano32aa1n02x4               g099(.a(new_n194), .b(new_n191), .c(new_n192), .d(new_n189), .out0(new_n195));
  aoi012aa1n02x5               g100(.a(new_n195), .b(new_n193), .c(new_n194), .o1(\s[17] ));
  norp02aa1n02x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[18] ), .b(\b[17] ), .out0(new_n198));
  aoi112aa1n02x5               g103(.a(new_n197), .b(new_n198), .c(new_n193), .d(new_n194), .o1(new_n199));
  aoai13aa1n03x5               g104(.a(new_n198), .b(new_n197), .c(new_n193), .d(new_n194), .o1(new_n200));
  norb02aa1n02x5               g105(.a(new_n200), .b(new_n199), .out0(\s[18] ));
  and002aa1n12x5               g106(.a(new_n198), .b(new_n194), .o(new_n202));
  nand02aa1n02x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  oai022aa1n03x5               g108(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n204));
  and002aa1n02x5               g109(.a(new_n204), .b(new_n203), .o(new_n205));
  xorc02aa1n12x5               g110(.a(\a[19] ), .b(\b[18] ), .out0(new_n206));
  aoai13aa1n09x5               g111(.a(new_n206), .b(new_n205), .c(new_n193), .d(new_n202), .o1(new_n207));
  aoi112aa1n02x5               g112(.a(new_n206), .b(new_n205), .c(new_n193), .d(new_n202), .o1(new_n208));
  norb02aa1n02x7               g113(.a(new_n207), .b(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n02x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  and002aa1n03x5               g116(.a(\b[19] ), .b(\a[20] ), .o(new_n212));
  nor042aa1n02x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  nor042aa1d18x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  oab012aa1n02x4               g119(.a(new_n214), .b(new_n212), .c(new_n211), .out0(new_n215));
  inv030aa1n02x5               g120(.a(new_n214), .o1(new_n216));
  tech160nm_finand02aa1n03p5x5 g121(.a(new_n207), .b(new_n216), .o1(new_n217));
  aoi022aa1n02x7               g122(.a(new_n217), .b(new_n213), .c(new_n207), .d(new_n215), .o1(\s[20] ));
  nand23aa1n06x5               g123(.a(new_n202), .b(new_n206), .c(new_n213), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoi112aa1n06x5               g125(.a(new_n212), .b(new_n211), .c(\a[19] ), .d(\b[18] ), .o1(new_n221));
  oai012aa1n02x7               g126(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .o1(new_n222));
  norb02aa1n03x5               g127(.a(new_n204), .b(new_n222), .out0(new_n223));
  oaoi03aa1n02x5               g128(.a(\a[20] ), .b(\b[19] ), .c(new_n216), .o1(new_n224));
  tech160nm_fiao0012aa1n02p5x5 g129(.a(new_n224), .b(new_n223), .c(new_n221), .o(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n09x5               g132(.a(new_n227), .b(new_n225), .c(new_n193), .d(new_n220), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n224), .b(new_n227), .c(new_n223), .d(new_n221), .o1(new_n229));
  aobi12aa1n02x5               g134(.a(new_n229), .b(new_n193), .c(new_n220), .out0(new_n230));
  norb02aa1n03x4               g135(.a(new_n228), .b(new_n230), .out0(\s[21] ));
  xnrc02aa1n12x5               g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  nor042aa1n06x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n232), .b(new_n234), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n234), .o1(new_n236));
  tech160nm_finand02aa1n03p5x5 g141(.a(new_n228), .b(new_n236), .o1(new_n237));
  aoi022aa1n02x7               g142(.a(new_n237), .b(new_n233), .c(new_n228), .d(new_n235), .o1(\s[22] ));
  nor042aa1n06x5               g143(.a(new_n232), .b(new_n226), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n219), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n239), .b(new_n224), .c(new_n223), .d(new_n221), .o1(new_n241));
  oao003aa1n02x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n236), .carry(new_n242));
  nanp02aa1n02x5               g147(.a(new_n241), .b(new_n242), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  aoai13aa1n09x5               g149(.a(new_n244), .b(new_n243), .c(new_n193), .d(new_n240), .o1(new_n245));
  nano22aa1n02x4               g150(.a(new_n244), .b(new_n241), .c(new_n242), .out0(new_n246));
  aobi12aa1n02x5               g151(.a(new_n246), .b(new_n193), .c(new_n240), .out0(new_n247));
  norb02aa1n03x4               g152(.a(new_n245), .b(new_n247), .out0(\s[23] ));
  tech160nm_fixorc02aa1n05x5   g153(.a(\a[24] ), .b(\b[23] ), .out0(new_n249));
  nor042aa1n03x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  norp02aa1n02x5               g155(.a(new_n249), .b(new_n250), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n250), .o1(new_n252));
  tech160nm_finand02aa1n03p5x5 g157(.a(new_n245), .b(new_n252), .o1(new_n253));
  aoi022aa1n02x7               g158(.a(new_n253), .b(new_n249), .c(new_n245), .d(new_n251), .o1(\s[24] ));
  and002aa1n02x5               g159(.a(new_n249), .b(new_n244), .o(new_n255));
  nano22aa1n02x5               g160(.a(new_n219), .b(new_n255), .c(new_n239), .out0(new_n256));
  inv000aa1n02x5               g161(.a(new_n255), .o1(new_n257));
  oao003aa1n02x5               g162(.a(\a[24] ), .b(\b[23] ), .c(new_n252), .carry(new_n258));
  aoai13aa1n12x5               g163(.a(new_n258), .b(new_n257), .c(new_n241), .d(new_n242), .o1(new_n259));
  tech160nm_fixorc02aa1n03p5x5 g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  aoai13aa1n09x5               g165(.a(new_n260), .b(new_n259), .c(new_n193), .d(new_n256), .o1(new_n261));
  nanb02aa1n02x5               g166(.a(new_n260), .b(new_n258), .out0(new_n262));
  aoi012aa1n02x5               g167(.a(new_n262), .b(new_n243), .c(new_n255), .o1(new_n263));
  aobi12aa1n02x5               g168(.a(new_n263), .b(new_n193), .c(new_n256), .out0(new_n264));
  norb02aa1n03x4               g169(.a(new_n261), .b(new_n264), .out0(\s[25] ));
  tech160nm_fixorc02aa1n03p5x5 g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  nor042aa1n03x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  norp02aa1n02x5               g172(.a(new_n266), .b(new_n267), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n267), .o1(new_n269));
  tech160nm_finand02aa1n05x5   g174(.a(new_n261), .b(new_n269), .o1(new_n270));
  aoi022aa1n02x7               g175(.a(new_n270), .b(new_n266), .c(new_n261), .d(new_n268), .o1(\s[26] ));
  and002aa1n02x5               g176(.a(new_n266), .b(new_n260), .o(new_n272));
  nano32aa1n06x5               g177(.a(new_n219), .b(new_n272), .c(new_n239), .d(new_n255), .out0(new_n273));
  nand22aa1n09x5               g178(.a(new_n193), .b(new_n273), .o1(new_n274));
  oao003aa1n02x5               g179(.a(\a[26] ), .b(\b[25] ), .c(new_n269), .carry(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoi012aa1n12x5               g181(.a(new_n276), .b(new_n259), .c(new_n272), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(new_n274), .b(new_n277), .o1(new_n278));
  xorc02aa1n12x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  aoi112aa1n02x5               g184(.a(new_n279), .b(new_n276), .c(new_n259), .d(new_n272), .o1(new_n280));
  aoi022aa1n02x5               g185(.a(new_n278), .b(new_n279), .c(new_n274), .d(new_n280), .o1(\s[27] ));
  nanp02aa1n09x5               g186(.a(new_n259), .b(new_n272), .o1(new_n282));
  nanp02aa1n12x5               g187(.a(new_n282), .b(new_n275), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n279), .b(new_n283), .c(new_n193), .d(new_n273), .o1(new_n284));
  tech160nm_fixorc02aa1n03p5x5 g189(.a(\a[28] ), .b(\b[27] ), .out0(new_n285));
  norp02aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  norp02aa1n02x5               g191(.a(new_n285), .b(new_n286), .o1(new_n287));
  inv000aa1n03x5               g192(.a(new_n286), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n279), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n288), .b(new_n289), .c(new_n274), .d(new_n277), .o1(new_n290));
  aoi022aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n284), .d(new_n287), .o1(\s[28] ));
  and002aa1n02x5               g196(.a(new_n285), .b(new_n279), .o(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n283), .c(new_n193), .d(new_n273), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n292), .o1(new_n294));
  oao003aa1n02x5               g199(.a(\a[28] ), .b(\b[27] ), .c(new_n288), .carry(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n274), .d(new_n277), .o1(new_n296));
  tech160nm_fixorc02aa1n03p5x5 g201(.a(\a[29] ), .b(\b[28] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n295), .b(new_n297), .out0(new_n298));
  aoi022aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n293), .d(new_n298), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g205(.a(new_n289), .b(new_n285), .c(new_n297), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n283), .c(new_n193), .d(new_n273), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n301), .o1(new_n303));
  inv000aa1d42x5               g208(.a(\b[28] ), .o1(new_n304));
  inv000aa1d42x5               g209(.a(\a[29] ), .o1(new_n305));
  oaib12aa1n02x5               g210(.a(new_n295), .b(\b[28] ), .c(new_n305), .out0(new_n306));
  oaib12aa1n02x5               g211(.a(new_n306), .b(new_n304), .c(\a[29] ), .out0(new_n307));
  aoai13aa1n06x5               g212(.a(new_n307), .b(new_n303), .c(new_n274), .d(new_n277), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .out0(new_n309));
  oaoi13aa1n02x5               g214(.a(new_n309), .b(new_n306), .c(new_n305), .d(new_n304), .o1(new_n310));
  aoi022aa1n02x7               g215(.a(new_n308), .b(new_n309), .c(new_n302), .d(new_n310), .o1(\s[30] ));
  nanb02aa1n02x5               g216(.a(\b[30] ), .b(\a[31] ), .out0(new_n312));
  nanb02aa1n02x5               g217(.a(\a[31] ), .b(\b[30] ), .out0(new_n313));
  nanp02aa1n02x5               g218(.a(new_n313), .b(new_n312), .o1(new_n314));
  nano32aa1n02x5               g219(.a(new_n289), .b(new_n309), .c(new_n285), .d(new_n297), .out0(new_n315));
  aoai13aa1n06x5               g220(.a(new_n315), .b(new_n283), .c(new_n193), .d(new_n273), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n315), .o1(new_n317));
  norp02aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .o1(new_n318));
  aoi022aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n318), .b(new_n306), .c(new_n319), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n317), .c(new_n274), .d(new_n277), .o1(new_n321));
  oai112aa1n02x5               g226(.a(new_n312), .b(new_n313), .c(\b[29] ), .d(\a[30] ), .o1(new_n322));
  aoi012aa1n02x5               g227(.a(new_n322), .b(new_n306), .c(new_n319), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n314), .c(new_n316), .d(new_n323), .o1(\s[31] ));
  inv000aa1d42x5               g229(.a(new_n102), .o1(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[2] ), .b(\a[3] ), .out0(new_n326));
  oai012aa1n02x5               g231(.a(new_n100), .b(new_n99), .c(new_n101), .o1(new_n327));
  aboi22aa1n03x5               g232(.a(new_n105), .b(new_n325), .c(new_n327), .d(new_n326), .out0(\s[3] ));
  nanb02aa1n02x5               g233(.a(new_n105), .b(new_n325), .out0(new_n329));
  xorc02aa1n02x5               g234(.a(\a[4] ), .b(\b[3] ), .out0(new_n330));
  aoib12aa1n02x5               g235(.a(new_n330), .b(new_n103), .c(\b[2] ), .out0(new_n331));
  aoi022aa1n02x5               g236(.a(new_n329), .b(new_n331), .c(new_n109), .d(new_n330), .o1(\s[4] ));
  and002aa1n02x5               g237(.a(\b[3] ), .b(\a[4] ), .o(new_n333));
  inv000aa1d42x5               g238(.a(new_n333), .o1(new_n334));
  nanb02aa1n02x5               g239(.a(new_n115), .b(new_n116), .out0(new_n335));
  xnbna2aa1n03x5               g240(.a(new_n335), .b(new_n109), .c(new_n334), .out0(\s[5] ));
  inv000aa1d42x5               g241(.a(new_n115), .o1(new_n337));
  nona22aa1n02x4               g242(.a(new_n109), .b(new_n333), .c(new_n335), .out0(new_n338));
  xobna2aa1n03x5               g243(.a(new_n114), .b(new_n338), .c(new_n337), .out0(\s[6] ));
  nanb02aa1n02x5               g244(.a(new_n110), .b(new_n112), .out0(new_n340));
  inv000aa1d42x5               g245(.a(new_n340), .o1(new_n341));
  nanp02aa1n02x5               g246(.a(new_n123), .b(new_n122), .o1(new_n342));
  nona32aa1n02x4               g247(.a(new_n109), .b(new_n335), .c(new_n114), .d(new_n333), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n341), .b(new_n343), .c(new_n342), .out0(\s[7] ));
  norb02aa1n02x5               g249(.a(new_n118), .b(new_n117), .out0(new_n345));
  aob012aa1n02x5               g250(.a(new_n341), .b(new_n343), .c(new_n342), .out0(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n345), .b(new_n346), .c(new_n111), .out0(\s[8] ));
  oaib12aa1n02x5               g252(.a(new_n125), .b(new_n97), .c(new_n127), .out0(new_n348));
  aoib12aa1n02x5               g253(.a(new_n348), .b(new_n121), .c(new_n124), .out0(new_n349));
  aoi022aa1n02x5               g254(.a(new_n167), .b(new_n128), .c(new_n166), .d(new_n349), .o1(\s[9] ));
endmodule


