// Benchmark "adder" written by ABC on Wed Jul 17 23:04:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n325, new_n326, new_n328, new_n331, new_n332, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv040aa1d32x5               g002(.a(\a[9] ), .o1(new_n98));
  inv040aa1d32x5               g003(.a(\b[8] ), .o1(new_n99));
  nand02aa1n03x5               g004(.a(new_n99), .b(new_n98), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nand02aa1n06x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nand02aa1n04x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nona23aa1d18x5               g010(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\b[5] ), .o1(new_n107));
  nanb02aa1d24x5               g012(.a(\a[6] ), .b(new_n107), .out0(new_n108));
  nand02aa1n10x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  oai112aa1n06x5               g014(.a(new_n108), .b(new_n109), .c(\b[4] ), .d(\a[5] ), .o1(new_n110));
  aoi112aa1n09x5               g015(.a(new_n106), .b(new_n110), .c(\a[5] ), .d(\b[4] ), .o1(new_n111));
  and002aa1n02x7               g016(.a(\b[3] ), .b(\a[4] ), .o(new_n112));
  nand22aa1n03x5               g017(.a(\b[0] ), .b(\a[1] ), .o1(new_n113));
  nanp02aa1n12x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  nor002aa1n03x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  norb03aa1n09x5               g020(.a(new_n114), .b(new_n113), .c(new_n115), .out0(new_n116));
  nor022aa1n16x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  nand02aa1n06x5               g022(.a(\b[2] ), .b(\a[3] ), .o1(new_n118));
  nanb03aa1n12x5               g023(.a(new_n117), .b(new_n118), .c(new_n114), .out0(new_n119));
  oab012aa1n04x5               g024(.a(new_n117), .b(\a[4] ), .c(\b[3] ), .out0(new_n120));
  oaoi13aa1n06x5               g025(.a(new_n112), .b(new_n120), .c(new_n116), .d(new_n119), .o1(new_n121));
  aoi112aa1n06x5               g026(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n122));
  nano23aa1n02x4               g027(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n123));
  nanp03aa1n02x5               g028(.a(new_n123), .b(new_n109), .c(new_n110), .o1(new_n124));
  nona22aa1n02x4               g029(.a(new_n124), .b(new_n122), .c(new_n102), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n101), .b(new_n125), .c(new_n111), .d(new_n121), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n100), .out0(\s[10] ));
  and002aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  inv020aa1n02x5               g033(.a(new_n112), .o1(new_n129));
  oai012aa1n12x5               g034(.a(new_n120), .b(new_n116), .c(new_n119), .o1(new_n130));
  nand23aa1d12x5               g035(.a(new_n111), .b(new_n130), .c(new_n129), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n102), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n122), .o1(new_n133));
  nano22aa1n03x7               g038(.a(new_n106), .b(new_n110), .c(new_n109), .out0(new_n134));
  nano22aa1n09x5               g039(.a(new_n134), .b(new_n132), .c(new_n133), .out0(new_n135));
  aobi12aa1n06x5               g040(.a(new_n101), .b(new_n131), .c(new_n135), .out0(new_n136));
  nano22aa1n03x7               g041(.a(new_n136), .b(new_n97), .c(new_n100), .out0(new_n137));
  nor002aa1d32x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand42aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  oab012aa1n02x4               g045(.a(new_n140), .b(new_n137), .c(new_n128), .out0(new_n141));
  nand42aa1n20x5               g046(.a(\b[9] ), .b(\a[10] ), .o1(new_n142));
  nano22aa1n03x7               g047(.a(new_n137), .b(new_n142), .c(new_n140), .out0(new_n143));
  norp02aa1n02x5               g048(.a(new_n141), .b(new_n143), .o1(\s[11] ));
  inv000aa1n06x5               g049(.a(new_n138), .o1(new_n145));
  nor002aa1d32x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand02aa1n06x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanb02aa1n02x5               g052(.a(new_n146), .b(new_n147), .out0(new_n148));
  nano22aa1n02x4               g053(.a(new_n143), .b(new_n145), .c(new_n148), .out0(new_n149));
  oab012aa1n02x4               g054(.a(new_n148), .b(new_n143), .c(new_n138), .out0(new_n150));
  norp02aa1n02x5               g055(.a(new_n150), .b(new_n149), .o1(\s[12] ));
  nanp02aa1n24x5               g056(.a(new_n131), .b(new_n135), .o1(new_n152));
  nand22aa1n03x5               g057(.a(new_n100), .b(new_n101), .o1(new_n153));
  nona23aa1n09x5               g058(.a(new_n147), .b(new_n139), .c(new_n138), .d(new_n146), .out0(new_n154));
  norb02aa1n06x5               g059(.a(new_n97), .b(new_n154), .out0(new_n155));
  nanb03aa1n09x5               g060(.a(new_n153), .b(new_n152), .c(new_n155), .out0(new_n156));
  nor002aa1d32x5               g061(.a(\b[9] ), .b(\a[10] ), .o1(new_n157));
  aoai13aa1n12x5               g062(.a(new_n142), .b(new_n157), .c(new_n98), .d(new_n99), .o1(new_n158));
  oaoi03aa1n09x5               g063(.a(\a[12] ), .b(\b[11] ), .c(new_n145), .o1(new_n159));
  oabi12aa1n18x5               g064(.a(new_n159), .b(new_n154), .c(new_n158), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[12] ), .b(\a[13] ), .out0(new_n162));
  xobna2aa1n03x5               g067(.a(new_n162), .b(new_n156), .c(new_n161), .out0(\s[13] ));
  tech160nm_fiao0012aa1n02p5x5 g068(.a(new_n162), .b(new_n156), .c(new_n161), .o(new_n164));
  inv040aa1d32x5               g069(.a(\a[14] ), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[13] ), .o1(new_n166));
  nanp02aa1n04x5               g071(.a(new_n166), .b(new_n165), .o1(new_n167));
  nor002aa1n03x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  oaoi03aa1n12x5               g073(.a(new_n165), .b(new_n166), .c(new_n168), .o1(new_n169));
  nand42aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nano22aa1d15x5               g075(.a(new_n162), .b(new_n167), .c(new_n170), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n169), .b(new_n172), .c(new_n156), .d(new_n161), .o1(new_n173));
  aoi012aa1n02x5               g078(.a(new_n168), .b(new_n167), .c(new_n170), .o1(new_n174));
  aoi022aa1n02x5               g079(.a(new_n164), .b(new_n174), .c(new_n173), .d(new_n167), .o1(\s[14] ));
  xorb03aa1n03x5               g080(.a(new_n173), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  xnrc02aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .out0(new_n177));
  nanb02aa1n03x5               g082(.a(new_n177), .b(new_n173), .out0(new_n178));
  inv000aa1d42x5               g083(.a(\a[16] ), .o1(new_n179));
  inv000aa1d42x5               g084(.a(\b[15] ), .o1(new_n180));
  nand42aa1n02x5               g085(.a(new_n180), .b(new_n179), .o1(new_n181));
  norp02aa1n02x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n182), .b(new_n181), .c(new_n183), .o1(new_n184));
  nano22aa1n03x7               g089(.a(new_n177), .b(new_n181), .c(new_n183), .out0(new_n185));
  nano23aa1n09x5               g090(.a(new_n138), .b(new_n146), .c(new_n147), .d(new_n139), .out0(new_n186));
  nona32aa1n09x5               g091(.a(new_n186), .b(new_n153), .c(new_n128), .d(new_n157), .out0(new_n187));
  nano22aa1n12x5               g092(.a(new_n187), .b(new_n171), .c(new_n185), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n125), .c(new_n111), .d(new_n121), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n169), .o1(new_n190));
  aoai13aa1n03x5               g095(.a(new_n185), .b(new_n190), .c(new_n160), .d(new_n171), .o1(new_n191));
  oaoi03aa1n02x5               g096(.a(new_n179), .b(new_n180), .c(new_n182), .o1(new_n192));
  nand23aa1n03x5               g097(.a(new_n189), .b(new_n191), .c(new_n192), .o1(new_n193));
  aoi022aa1n02x5               g098(.a(new_n178), .b(new_n184), .c(new_n181), .d(new_n193), .o1(\s[16] ));
  xorb03aa1n02x5               g099(.a(new_n193), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor002aa1d32x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  and002aa1n03x5               g101(.a(\b[14] ), .b(\a[15] ), .o(new_n197));
  nona23aa1n06x5               g102(.a(new_n181), .b(new_n183), .c(new_n197), .d(new_n182), .out0(new_n198));
  nona23aa1n03x5               g103(.a(new_n155), .b(new_n171), .c(new_n198), .d(new_n153), .out0(new_n199));
  aoi012aa1n06x5               g104(.a(new_n199), .b(new_n131), .c(new_n135), .o1(new_n200));
  inv040aa1n02x5               g105(.a(new_n158), .o1(new_n201));
  aoai13aa1n06x5               g106(.a(new_n171), .b(new_n159), .c(new_n186), .d(new_n201), .o1(new_n202));
  aoai13aa1n12x5               g107(.a(new_n192), .b(new_n198), .c(new_n202), .d(new_n169), .o1(new_n203));
  tech160nm_fixorc02aa1n05x5   g108(.a(\a[17] ), .b(\b[16] ), .out0(new_n204));
  nand42aa1d28x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nano22aa1n12x5               g110(.a(new_n196), .b(new_n204), .c(new_n205), .out0(new_n206));
  inv040aa1d30x5               g111(.a(\a[17] ), .o1(new_n207));
  inv040aa1d32x5               g112(.a(\b[16] ), .o1(new_n208));
  aoai13aa1n12x5               g113(.a(new_n205), .b(new_n196), .c(new_n207), .d(new_n208), .o1(new_n209));
  inv000aa1n06x5               g114(.a(new_n209), .o1(new_n210));
  oaoi13aa1n06x5               g115(.a(new_n210), .b(new_n206), .c(new_n200), .d(new_n203), .o1(new_n211));
  obai22aa1n02x7               g116(.a(new_n205), .b(new_n196), .c(\a[17] ), .d(\b[16] ), .out0(new_n212));
  oaoi13aa1n02x5               g117(.a(new_n212), .b(new_n204), .c(new_n200), .d(new_n203), .o1(new_n213));
  oab012aa1n02x4               g118(.a(new_n213), .b(new_n211), .c(new_n196), .out0(\s[18] ));
  aoai13aa1n06x5               g119(.a(new_n206), .b(new_n203), .c(new_n152), .d(new_n188), .o1(new_n215));
  nor002aa1d32x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  nand42aa1n06x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nanb02aa1n12x5               g122(.a(new_n216), .b(new_n217), .out0(new_n218));
  xobna2aa1n03x5               g123(.a(new_n218), .b(new_n215), .c(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g125(.a(new_n216), .o1(new_n221));
  aoi012aa1n02x5               g126(.a(new_n218), .b(new_n215), .c(new_n209), .o1(new_n222));
  nor002aa1d24x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nand02aa1n10x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  nanb02aa1n06x5               g129(.a(new_n223), .b(new_n224), .out0(new_n225));
  nano22aa1n03x5               g130(.a(new_n222), .b(new_n221), .c(new_n225), .out0(new_n226));
  oaoi13aa1n03x5               g131(.a(new_n225), .b(new_n221), .c(new_n211), .d(new_n218), .o1(new_n227));
  norp02aa1n03x5               g132(.a(new_n227), .b(new_n226), .o1(\s[20] ));
  nano23aa1n09x5               g133(.a(new_n216), .b(new_n223), .c(new_n224), .d(new_n217), .out0(new_n229));
  nand22aa1n04x5               g134(.a(new_n206), .b(new_n229), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n203), .c(new_n152), .d(new_n188), .o1(new_n232));
  aoi012aa1n06x5               g137(.a(new_n223), .b(new_n216), .c(new_n224), .o1(new_n233));
  oai013aa1d12x5               g138(.a(new_n233), .b(new_n209), .c(new_n218), .d(new_n225), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .out0(new_n236));
  xobna2aa1n03x5               g141(.a(new_n236), .b(new_n232), .c(new_n235), .out0(\s[21] ));
  nor002aa1d32x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoi012aa1n02x7               g144(.a(new_n236), .b(new_n232), .c(new_n235), .o1(new_n240));
  tech160nm_fixnrc02aa1n04x5   g145(.a(\b[21] ), .b(\a[22] ), .out0(new_n241));
  nano22aa1n03x7               g146(.a(new_n240), .b(new_n239), .c(new_n241), .out0(new_n242));
  oaoi13aa1n03x5               g147(.a(new_n234), .b(new_n231), .c(new_n200), .d(new_n203), .o1(new_n243));
  oaoi13aa1n03x5               g148(.a(new_n241), .b(new_n239), .c(new_n243), .d(new_n236), .o1(new_n244));
  norp02aa1n03x5               g149(.a(new_n244), .b(new_n242), .o1(\s[22] ));
  nor042aa1n04x5               g150(.a(new_n241), .b(new_n236), .o1(new_n246));
  and003aa1n02x5               g151(.a(new_n206), .b(new_n246), .c(new_n229), .o(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n203), .c(new_n152), .d(new_n188), .o1(new_n248));
  oao003aa1n12x5               g153(.a(\a[22] ), .b(\b[21] ), .c(new_n239), .carry(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n250), .b(new_n234), .c(new_n246), .o1(new_n251));
  xnrc02aa1n12x5               g156(.a(\b[22] ), .b(\a[23] ), .out0(new_n252));
  xobna2aa1n03x5               g157(.a(new_n252), .b(new_n248), .c(new_n251), .out0(\s[23] ));
  nor042aa1n06x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  aoi012aa1n02x7               g160(.a(new_n252), .b(new_n248), .c(new_n251), .o1(new_n256));
  xnrc02aa1n12x5               g161(.a(\b[23] ), .b(\a[24] ), .out0(new_n257));
  nano22aa1n03x7               g162(.a(new_n256), .b(new_n255), .c(new_n257), .out0(new_n258));
  inv000aa1n03x5               g163(.a(new_n251), .o1(new_n259));
  oaoi13aa1n03x5               g164(.a(new_n259), .b(new_n247), .c(new_n200), .d(new_n203), .o1(new_n260));
  oaoi13aa1n03x5               g165(.a(new_n257), .b(new_n255), .c(new_n260), .d(new_n252), .o1(new_n261));
  norp02aa1n03x5               g166(.a(new_n261), .b(new_n258), .o1(\s[24] ));
  nor042aa1n02x5               g167(.a(new_n257), .b(new_n252), .o1(new_n263));
  nano22aa1n03x7               g168(.a(new_n230), .b(new_n246), .c(new_n263), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n203), .c(new_n152), .d(new_n188), .o1(new_n265));
  inv030aa1n02x5               g170(.a(new_n233), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n246), .b(new_n266), .c(new_n229), .d(new_n210), .o1(new_n267));
  inv000aa1n03x5               g172(.a(new_n263), .o1(new_n268));
  oao003aa1n02x5               g173(.a(\a[24] ), .b(\b[23] ), .c(new_n255), .carry(new_n269));
  aoai13aa1n12x5               g174(.a(new_n269), .b(new_n268), .c(new_n267), .d(new_n249), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  xnrc02aa1n12x5               g176(.a(\b[24] ), .b(\a[25] ), .out0(new_n272));
  xobna2aa1n03x5               g177(.a(new_n272), .b(new_n265), .c(new_n271), .out0(\s[25] ));
  nor042aa1n03x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n274), .o1(new_n275));
  tech160nm_fiaoi012aa1n02p5x5 g180(.a(new_n272), .b(new_n265), .c(new_n271), .o1(new_n276));
  xnrc02aa1n12x5               g181(.a(\b[25] ), .b(\a[26] ), .out0(new_n277));
  nano22aa1n03x7               g182(.a(new_n276), .b(new_n275), .c(new_n277), .out0(new_n278));
  oaoi13aa1n02x7               g183(.a(new_n270), .b(new_n264), .c(new_n200), .d(new_n203), .o1(new_n279));
  oaoi13aa1n03x5               g184(.a(new_n277), .b(new_n275), .c(new_n279), .d(new_n272), .o1(new_n280));
  nor002aa1n02x5               g185(.a(new_n280), .b(new_n278), .o1(\s[26] ));
  nor042aa1n06x5               g186(.a(new_n277), .b(new_n272), .o1(new_n282));
  nano32aa1d15x5               g187(.a(new_n230), .b(new_n282), .c(new_n246), .d(new_n263), .out0(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n203), .c(new_n152), .d(new_n188), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[26] ), .b(\b[25] ), .c(new_n275), .carry(new_n285));
  aobi12aa1n18x5               g190(.a(new_n285), .b(new_n270), .c(new_n282), .out0(new_n286));
  xorc02aa1n12x5               g191(.a(\a[27] ), .b(\b[26] ), .out0(new_n287));
  xnbna2aa1n03x5               g192(.a(new_n287), .b(new_n284), .c(new_n286), .out0(\s[27] ));
  norp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  inv040aa1n03x5               g194(.a(new_n289), .o1(new_n290));
  aobi12aa1n06x5               g195(.a(new_n287), .b(new_n284), .c(new_n286), .out0(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .out0(new_n292));
  nano22aa1n03x7               g197(.a(new_n291), .b(new_n290), .c(new_n292), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n263), .b(new_n250), .c(new_n234), .d(new_n246), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n282), .o1(new_n295));
  aoai13aa1n04x5               g200(.a(new_n285), .b(new_n295), .c(new_n294), .d(new_n269), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n287), .b(new_n296), .c(new_n193), .d(new_n283), .o1(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n292), .b(new_n297), .c(new_n290), .o1(new_n298));
  norp02aa1n03x5               g203(.a(new_n298), .b(new_n293), .o1(\s[28] ));
  xnrc02aa1n02x5               g204(.a(\b[28] ), .b(\a[29] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n287), .b(new_n292), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n296), .c(new_n193), .d(new_n283), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n290), .carry(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n300), .b(new_n302), .c(new_n303), .o1(new_n304));
  aobi12aa1n06x5               g209(.a(new_n301), .b(new_n284), .c(new_n286), .out0(new_n305));
  nano22aa1n03x7               g210(.a(new_n305), .b(new_n300), .c(new_n303), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n304), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n113), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g213(.a(new_n287), .b(new_n300), .c(new_n292), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n296), .c(new_n193), .d(new_n283), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .out0(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n312), .b(new_n310), .c(new_n311), .o1(new_n313));
  aobi12aa1n06x5               g218(.a(new_n309), .b(new_n284), .c(new_n286), .out0(new_n314));
  nano22aa1n03x7               g219(.a(new_n314), .b(new_n311), .c(new_n312), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n313), .b(new_n315), .o1(\s[30] ));
  xnrc02aa1n02x5               g221(.a(\b[30] ), .b(\a[31] ), .out0(new_n317));
  norb02aa1n02x7               g222(.a(new_n309), .b(new_n312), .out0(new_n318));
  aobi12aa1n06x5               g223(.a(new_n318), .b(new_n284), .c(new_n286), .out0(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n320));
  nano22aa1n03x7               g225(.a(new_n319), .b(new_n317), .c(new_n320), .out0(new_n321));
  aoai13aa1n02x5               g226(.a(new_n318), .b(new_n296), .c(new_n193), .d(new_n283), .o1(new_n322));
  tech160nm_fiaoi012aa1n02p5x5 g227(.a(new_n317), .b(new_n322), .c(new_n320), .o1(new_n323));
  norp02aa1n03x5               g228(.a(new_n323), .b(new_n321), .o1(\s[31] ));
  norb02aa1n02x5               g229(.a(new_n118), .b(new_n117), .out0(new_n325));
  oaoi13aa1n02x5               g230(.a(new_n325), .b(new_n114), .c(new_n113), .d(new_n115), .o1(new_n326));
  oab012aa1n02x4               g231(.a(new_n326), .b(new_n116), .c(new_n119), .out0(\s[3] ));
  oabi12aa1n02x5               g232(.a(new_n117), .b(new_n116), .c(new_n119), .out0(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g234(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanp02aa1n02x5               g235(.a(new_n130), .b(new_n129), .o1(new_n331));
  oao003aa1n03x5               g236(.a(\a[5] ), .b(\b[4] ), .c(new_n331), .carry(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n108), .c(new_n109), .out0(\s[6] ));
  tech160nm_fioaoi03aa1n03p5x5 g238(.a(\a[6] ), .b(\b[5] ), .c(new_n332), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  tech160nm_fiaoi012aa1n05x5   g240(.a(new_n104), .b(new_n334), .c(new_n105), .o1(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n336), .b(new_n132), .c(new_n103), .out0(\s[8] ));
  xobna2aa1n03x5               g242(.a(new_n153), .b(new_n131), .c(new_n135), .out0(\s[9] ));
endmodule


