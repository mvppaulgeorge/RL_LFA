// Benchmark "adder" written by ABC on Wed Jul 17 16:18:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n332, new_n335, new_n337, new_n338, new_n339, new_n341, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  nor042aa1n04x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n06x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand02aa1d12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  tech160nm_fiaoi012aa1n05x5   g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  inv000aa1n04x5               g007(.a(new_n102), .o1(new_n103));
  nor002aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand42aa1n20x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n06x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n08x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nano23aa1n03x5               g012(.a(new_n104), .b(new_n106), .c(new_n107), .d(new_n105), .out0(new_n108));
  inv030aa1n02x5               g013(.a(new_n106), .o1(new_n109));
  oaoi03aa1n09x5               g014(.a(\a[4] ), .b(\b[3] ), .c(new_n109), .o1(new_n110));
  aoi012aa1n06x5               g015(.a(new_n110), .b(new_n108), .c(new_n103), .o1(new_n111));
  tech160nm_fixorc02aa1n03p5x5 g016(.a(\a[5] ), .b(\b[4] ), .out0(new_n112));
  nor002aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand02aa1n08x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  norb02aa1n06x5               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  nor002aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n06x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nor002aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1n03x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nanp03aa1n04x5               g025(.a(new_n120), .b(new_n112), .c(new_n115), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\a[8] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[7] ), .o1(new_n123));
  inv000aa1n06x5               g028(.a(new_n116), .o1(new_n124));
  nor042aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  aoai13aa1n03x5               g030(.a(new_n117), .b(new_n113), .c(new_n125), .d(new_n114), .o1(new_n126));
  nanp02aa1n03x5               g031(.a(new_n126), .b(new_n124), .o1(new_n127));
  oaoi03aa1n12x5               g032(.a(new_n122), .b(new_n123), .c(new_n127), .o1(new_n128));
  oai012aa1n12x5               g033(.a(new_n128), .b(new_n111), .c(new_n121), .o1(new_n129));
  xnrc02aa1n12x5               g034(.a(\b[8] ), .b(\a[9] ), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  aoi012aa1n02x5               g036(.a(new_n98), .b(new_n129), .c(new_n131), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  xnrc02aa1n02x5               g038(.a(\b[9] ), .b(\a[10] ), .out0(new_n134));
  nor042aa1n02x5               g039(.a(new_n130), .b(new_n134), .o1(new_n135));
  inv000aa1d42x5               g040(.a(\b[9] ), .o1(new_n136));
  oao003aa1n02x5               g041(.a(new_n97), .b(new_n136), .c(new_n98), .carry(new_n137));
  xnrc02aa1n12x5               g042(.a(\b[10] ), .b(\a[11] ), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  aoai13aa1n03x5               g044(.a(new_n139), .b(new_n137), .c(new_n129), .d(new_n135), .o1(new_n140));
  aoi112aa1n02x5               g045(.a(new_n139), .b(new_n137), .c(new_n129), .d(new_n135), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(\s[11] ));
  nor042aa1n04x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n143), .o1(new_n144));
  nor022aa1n08x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand42aa1n04x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nanb02aa1n12x5               g051(.a(new_n145), .b(new_n146), .out0(new_n147));
  xobna2aa1n03x5               g052(.a(new_n147), .b(new_n140), .c(new_n144), .out0(\s[12] ));
  nanb02aa1n02x5               g053(.a(new_n104), .b(new_n105), .out0(new_n149));
  nanb02aa1n02x5               g054(.a(new_n106), .b(new_n107), .out0(new_n150));
  nor043aa1n03x5               g055(.a(new_n102), .b(new_n149), .c(new_n150), .o1(new_n151));
  nanb02aa1n02x5               g056(.a(new_n116), .b(new_n117), .out0(new_n152));
  norb02aa1n06x4               g057(.a(new_n119), .b(new_n118), .out0(new_n153));
  nano32aa1n02x4               g058(.a(new_n152), .b(new_n112), .c(new_n153), .d(new_n115), .out0(new_n154));
  oaih12aa1n06x5               g059(.a(new_n154), .b(new_n151), .c(new_n110), .o1(new_n155));
  nor042aa1n04x5               g060(.a(new_n138), .b(new_n147), .o1(new_n156));
  and002aa1n06x5               g061(.a(new_n135), .b(new_n156), .o(new_n157));
  inv000aa1n03x5               g062(.a(new_n157), .o1(new_n158));
  tech160nm_fioaoi03aa1n03p5x5 g063(.a(new_n97), .b(new_n136), .c(new_n98), .o1(new_n159));
  tech160nm_fiaoi012aa1n05x5   g064(.a(new_n145), .b(new_n143), .c(new_n146), .o1(new_n160));
  oai013aa1d12x5               g065(.a(new_n160), .b(new_n159), .c(new_n138), .d(new_n147), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n158), .c(new_n155), .d(new_n128), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand42aa1n04x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  tech160nm_fiaoi012aa1n05x5   g071(.a(new_n165), .b(new_n163), .c(new_n166), .o1(new_n167));
  xnrb03aa1n02x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1n06x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nano23aa1n06x5               g075(.a(new_n165), .b(new_n169), .c(new_n170), .d(new_n166), .out0(new_n171));
  aoai13aa1n03x5               g076(.a(new_n171), .b(new_n161), .c(new_n129), .d(new_n157), .o1(new_n172));
  aoi012aa1n09x5               g077(.a(new_n169), .b(new_n165), .c(new_n170), .o1(new_n173));
  xorc02aa1n06x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n172), .c(new_n173), .out0(\s[15] ));
  nanp02aa1n02x5               g080(.a(new_n172), .b(new_n173), .o1(new_n176));
  nor042aa1n03x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  xnrc02aa1n02x5               g082(.a(\b[15] ), .b(\a[16] ), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n177), .c(new_n176), .d(new_n174), .o1(new_n179));
  inv030aa1n02x5               g084(.a(new_n173), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n174), .b(new_n180), .c(new_n163), .d(new_n171), .o1(new_n181));
  nona22aa1n02x4               g086(.a(new_n181), .b(new_n178), .c(new_n177), .out0(new_n182));
  nanp02aa1n02x5               g087(.a(new_n179), .b(new_n182), .o1(\s[16] ));
  tech160nm_fixorc02aa1n02p5x5 g088(.a(\a[16] ), .b(\b[15] ), .out0(new_n184));
  nanp03aa1n09x5               g089(.a(new_n171), .b(new_n174), .c(new_n184), .o1(new_n185));
  nano22aa1n12x5               g090(.a(new_n185), .b(new_n135), .c(new_n156), .out0(new_n186));
  nand22aa1n03x5               g091(.a(new_n129), .b(new_n186), .o1(new_n187));
  nona23aa1n03x5               g092(.a(new_n170), .b(new_n166), .c(new_n165), .d(new_n169), .out0(new_n188));
  norb03aa1n09x5               g093(.a(new_n174), .b(new_n188), .c(new_n178), .out0(new_n189));
  nanb03aa1n02x5               g094(.a(new_n173), .b(new_n184), .c(new_n174), .out0(new_n190));
  inv000aa1d42x5               g095(.a(\a[16] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[15] ), .o1(new_n192));
  tech160nm_fioaoi03aa1n03p5x5 g097(.a(new_n191), .b(new_n192), .c(new_n177), .o1(new_n193));
  nand22aa1n02x5               g098(.a(new_n190), .b(new_n193), .o1(new_n194));
  aoi012aa1d18x5               g099(.a(new_n194), .b(new_n161), .c(new_n189), .o1(new_n195));
  xorc02aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n187), .c(new_n195), .out0(\s[17] ));
  inv040aa1d32x5               g102(.a(\a[18] ), .o1(new_n198));
  inv000aa1n06x5               g103(.a(new_n186), .o1(new_n199));
  aoai13aa1n12x5               g104(.a(new_n195), .b(new_n199), .c(new_n155), .d(new_n128), .o1(new_n200));
  norp02aa1n02x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  tech160nm_fiaoi012aa1n05x5   g106(.a(new_n201), .b(new_n200), .c(new_n196), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[17] ), .c(new_n198), .out0(\s[18] ));
  nona22aa1n09x5               g108(.a(new_n137), .b(new_n138), .c(new_n147), .out0(new_n204));
  inv030aa1n02x5               g109(.a(new_n193), .o1(new_n205));
  aoi013aa1n02x4               g110(.a(new_n205), .b(new_n180), .c(new_n174), .d(new_n184), .o1(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n185), .c(new_n204), .d(new_n160), .o1(new_n207));
  inv000aa1d42x5               g112(.a(\a[17] ), .o1(new_n208));
  xroi22aa1d06x4               g113(.a(new_n208), .b(\b[16] ), .c(new_n198), .d(\b[17] ), .out0(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n207), .c(new_n129), .d(new_n186), .o1(new_n210));
  nor002aa1n02x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  aoi112aa1n09x5               g116(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n212));
  nor002aa1n02x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  norp02aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand42aa1n06x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norb02aa1n06x4               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n210), .c(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand22aa1n03x5               g123(.a(new_n210), .b(new_n213), .o1(new_n219));
  nor002aa1n06x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nanp02aa1n24x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  norb02aa1n12x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n214), .c(new_n219), .d(new_n215), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n213), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n216), .b(new_n225), .c(new_n200), .d(new_n209), .o1(new_n226));
  nona22aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n214), .out0(new_n227));
  nanp02aa1n03x5               g132(.a(new_n224), .b(new_n227), .o1(\s[20] ));
  nano23aa1n06x5               g133(.a(new_n214), .b(new_n220), .c(new_n221), .d(new_n215), .out0(new_n229));
  nand02aa1d04x5               g134(.a(new_n209), .b(new_n229), .o1(new_n230));
  oai112aa1n06x5               g135(.a(new_n216), .b(new_n222), .c(new_n212), .d(new_n211), .o1(new_n231));
  aoi012aa1n02x7               g136(.a(new_n220), .b(new_n214), .c(new_n221), .o1(new_n232));
  nand02aa1d08x5               g137(.a(new_n231), .b(new_n232), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n230), .c(new_n187), .d(new_n195), .o1(new_n235));
  xorb03aa1n02x5               g140(.a(new_n235), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n04x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[21] ), .b(\b[20] ), .out0(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  aoai13aa1n02x7               g144(.a(new_n239), .b(new_n237), .c(new_n235), .d(new_n238), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n230), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n238), .b(new_n233), .c(new_n200), .d(new_n241), .o1(new_n242));
  nona22aa1n03x5               g147(.a(new_n242), .b(new_n239), .c(new_n237), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n240), .b(new_n243), .o1(\s[22] ));
  nanb02aa1n02x5               g149(.a(new_n239), .b(new_n238), .out0(new_n245));
  nano22aa1n02x4               g150(.a(new_n245), .b(new_n209), .c(new_n229), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n207), .c(new_n129), .d(new_n186), .o1(new_n247));
  norb02aa1n03x5               g152(.a(new_n238), .b(new_n239), .out0(new_n248));
  inv000aa1d42x5               g153(.a(\a[22] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\b[21] ), .o1(new_n250));
  oao003aa1n03x5               g155(.a(new_n249), .b(new_n250), .c(new_n237), .carry(new_n251));
  aoi012aa1n02x7               g156(.a(new_n251), .b(new_n233), .c(new_n248), .o1(new_n252));
  tech160nm_fixorc02aa1n03p5x5 g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  xnbna2aa1n03x5               g158(.a(new_n253), .b(new_n247), .c(new_n252), .out0(\s[23] ));
  nanp02aa1n02x5               g159(.a(new_n247), .b(new_n252), .o1(new_n255));
  norp02aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  xnrc02aa1n12x5               g161(.a(\b[23] ), .b(\a[24] ), .out0(new_n257));
  aoai13aa1n02x5               g162(.a(new_n257), .b(new_n256), .c(new_n255), .d(new_n253), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n252), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n253), .b(new_n259), .c(new_n200), .d(new_n246), .o1(new_n260));
  nona22aa1n03x5               g165(.a(new_n260), .b(new_n257), .c(new_n256), .out0(new_n261));
  nanp02aa1n03x5               g166(.a(new_n258), .b(new_n261), .o1(\s[24] ));
  tech160nm_fixnrc02aa1n02p5x5 g167(.a(\b[22] ), .b(\a[23] ), .out0(new_n263));
  nor042aa1n02x5               g168(.a(new_n257), .b(new_n263), .o1(new_n264));
  nano32aa1n03x7               g169(.a(new_n245), .b(new_n209), .c(new_n264), .d(new_n229), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n207), .c(new_n129), .d(new_n186), .o1(new_n266));
  norp02aa1n02x5               g171(.a(\b[23] ), .b(\a[24] ), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n268));
  nona22aa1n02x4               g173(.a(new_n251), .b(new_n263), .c(new_n257), .out0(new_n269));
  nona22aa1n02x4               g174(.a(new_n269), .b(new_n268), .c(new_n267), .out0(new_n270));
  aoi013aa1n09x5               g175(.a(new_n270), .b(new_n233), .c(new_n248), .d(new_n264), .o1(new_n271));
  tech160nm_fixorc02aa1n03p5x5 g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n266), .c(new_n271), .out0(\s[25] ));
  nand42aa1n03x5               g178(.a(new_n266), .b(new_n271), .o1(new_n274));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  aoai13aa1n02x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .d(new_n272), .o1(new_n277));
  inv020aa1n02x5               g182(.a(new_n271), .o1(new_n278));
  aoai13aa1n02x7               g183(.a(new_n272), .b(new_n278), .c(new_n200), .d(new_n265), .o1(new_n279));
  nona22aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n275), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n277), .b(new_n280), .o1(\s[26] ));
  norb02aa1n02x5               g186(.a(new_n272), .b(new_n276), .out0(new_n282));
  nano32aa1n03x7               g187(.a(new_n230), .b(new_n282), .c(new_n248), .d(new_n264), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n207), .c(new_n129), .d(new_n186), .o1(new_n284));
  nanb02aa1n02x5               g189(.a(new_n257), .b(new_n253), .out0(new_n285));
  aoi112aa1n03x5               g190(.a(new_n245), .b(new_n285), .c(new_n231), .d(new_n232), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\a[26] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[25] ), .o1(new_n288));
  tech160nm_fioaoi03aa1n03p5x5 g193(.a(new_n287), .b(new_n288), .c(new_n275), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  oaoi13aa1n04x5               g195(.a(new_n290), .b(new_n282), .c(new_n286), .d(new_n270), .o1(new_n291));
  xorc02aa1n12x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  xnbna2aa1n03x5               g197(.a(new_n292), .b(new_n284), .c(new_n291), .out0(\s[27] ));
  nand02aa1n03x5               g198(.a(new_n284), .b(new_n291), .o1(new_n294));
  norp02aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  xnrc02aa1n06x5               g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n295), .c(new_n294), .d(new_n292), .o1(new_n297));
  oai012aa1n03x5               g202(.a(new_n282), .b(new_n286), .c(new_n270), .o1(new_n298));
  nand42aa1n03x5               g203(.a(new_n298), .b(new_n289), .o1(new_n299));
  aoai13aa1n02x7               g204(.a(new_n292), .b(new_n299), .c(new_n200), .d(new_n283), .o1(new_n300));
  nona22aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n297), .b(new_n301), .o1(\s[28] ));
  norb02aa1n12x5               g207(.a(new_n292), .b(new_n296), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n299), .c(new_n200), .d(new_n283), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n303), .o1(new_n305));
  orn002aa1n03x5               g210(.a(\a[27] ), .b(\b[26] ), .o(new_n306));
  oao003aa1n02x5               g211(.a(\a[28] ), .b(\b[27] ), .c(new_n306), .carry(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n305), .c(new_n284), .d(new_n291), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n307), .b(new_n309), .out0(new_n310));
  aoi022aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n304), .d(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g216(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g217(.a(new_n296), .b(new_n292), .c(new_n309), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n299), .c(new_n200), .d(new_n283), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  oaoi03aa1n09x5               g220(.a(\a[29] ), .b(\b[28] ), .c(new_n307), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n316), .o1(new_n317));
  aoai13aa1n02x5               g222(.a(new_n317), .b(new_n315), .c(new_n284), .d(new_n291), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  and002aa1n02x5               g224(.a(\b[28] ), .b(\a[29] ), .o(new_n320));
  oabi12aa1n02x5               g225(.a(new_n319), .b(\a[29] ), .c(\b[28] ), .out0(new_n321));
  oab012aa1n02x4               g226(.a(new_n321), .b(new_n307), .c(new_n320), .out0(new_n322));
  aoi022aa1n03x5               g227(.a(new_n318), .b(new_n319), .c(new_n314), .d(new_n322), .o1(\s[30] ));
  nanp03aa1n02x5               g228(.a(new_n303), .b(new_n309), .c(new_n319), .o1(new_n324));
  nanb02aa1n03x5               g229(.a(new_n324), .b(new_n294), .out0(new_n325));
  xorc02aa1n02x5               g230(.a(\a[31] ), .b(\b[30] ), .out0(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n327));
  norb02aa1n02x5               g232(.a(new_n327), .b(new_n326), .out0(new_n328));
  aoai13aa1n03x5               g233(.a(new_n327), .b(new_n324), .c(new_n284), .d(new_n291), .o1(new_n329));
  aoi022aa1n03x5               g234(.a(new_n325), .b(new_n328), .c(new_n329), .d(new_n326), .o1(\s[31] ));
  xnbna2aa1n03x5               g235(.a(new_n102), .b(new_n107), .c(new_n109), .out0(\s[3] ));
  oai112aa1n02x5               g236(.a(new_n109), .b(new_n149), .c(new_n102), .d(new_n150), .o1(new_n332));
  oa0012aa1n02x5               g237(.a(new_n332), .b(new_n111), .c(new_n104), .o(\s[4] ));
  xnrc02aa1n02x5               g238(.a(new_n111), .b(new_n112), .out0(\s[5] ));
  oaoi13aa1n04x5               g239(.a(new_n125), .b(new_n112), .c(new_n151), .d(new_n110), .o1(new_n335));
  xnrc02aa1n02x5               g240(.a(new_n335), .b(new_n115), .out0(\s[6] ));
  aob012aa1n02x5               g241(.a(new_n114), .b(new_n335), .c(new_n115), .out0(new_n337));
  and002aa1n03x5               g242(.a(new_n335), .b(new_n115), .o(new_n338));
  nano32aa1n02x5               g243(.a(new_n338), .b(new_n117), .c(new_n124), .d(new_n114), .out0(new_n339));
  aoi012aa1n02x5               g244(.a(new_n339), .b(new_n152), .c(new_n337), .o1(\s[7] ));
  oabi12aa1n02x5               g245(.a(new_n153), .b(new_n339), .c(new_n116), .out0(new_n341));
  nano22aa1n03x7               g246(.a(new_n339), .b(new_n124), .c(new_n153), .out0(new_n342));
  nanb02aa1n02x5               g247(.a(new_n342), .b(new_n341), .out0(\s[8] ));
  xorb03aa1n02x5               g248(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


