// Benchmark "adder" written by ABC on Wed Jul 17 19:13:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n176,
    new_n177, new_n178, new_n179, new_n180, new_n181, new_n182, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n361, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n387,
    new_n388, new_n390, new_n391, new_n392, new_n394, new_n395, new_n397,
    new_n398, new_n400, new_n401, new_n403;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n03x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  oai112aa1n06x5               g002(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n98));
  nand42aa1n03x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nor022aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1n03x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  norb02aa1n03x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  tech160nm_finand02aa1n03p5x5 g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nona22aa1n02x4               g009(.a(new_n103), .b(new_n104), .c(new_n100), .out0(new_n105));
  aoi013aa1n06x4               g010(.a(new_n105), .b(new_n102), .c(new_n99), .d(new_n98), .o1(new_n106));
  nor042aa1d18x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  norp02aa1n04x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand42aa1n08x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  norb03aa1n09x5               g014(.a(new_n109), .b(new_n107), .c(new_n108), .out0(new_n110));
  aob012aa1n02x5               g015(.a(new_n103), .b(\b[4] ), .c(\a[5] ), .out0(new_n111));
  oai022aa1n02x5               g016(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n112));
  aoi022aa1d24x5               g017(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n113));
  nona23aa1n09x5               g018(.a(new_n110), .b(new_n113), .c(new_n111), .d(new_n112), .out0(new_n114));
  inv000aa1n02x5               g019(.a(new_n107), .o1(new_n115));
  oaoi03aa1n03x5               g020(.a(\a[8] ), .b(\b[7] ), .c(new_n115), .o1(new_n116));
  norp02aa1n06x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  inv000aa1n02x5               g022(.a(new_n117), .o1(new_n118));
  nand22aa1n02x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  oai112aa1n06x5               g024(.a(new_n118), .b(new_n119), .c(\b[4] ), .d(\a[5] ), .o1(new_n120));
  aoi013aa1n06x4               g025(.a(new_n116), .b(new_n120), .c(new_n110), .d(new_n113), .o1(new_n121));
  oai012aa1d24x5               g026(.a(new_n121), .b(new_n106), .c(new_n114), .o1(new_n122));
  nor042aa1n06x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  tech160nm_fixorc02aa1n02p5x5 g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoi112aa1n02x5               g029(.a(new_n123), .b(new_n97), .c(new_n122), .d(new_n124), .o1(new_n125));
  inv020aa1n02x5               g030(.a(new_n98), .o1(new_n126));
  nanb03aa1n06x5               g031(.a(new_n100), .b(new_n101), .c(new_n99), .out0(new_n127));
  norb03aa1n03x4               g032(.a(new_n103), .b(new_n100), .c(new_n104), .out0(new_n128));
  tech160nm_fioai012aa1n05x5   g033(.a(new_n128), .b(new_n127), .c(new_n126), .o1(new_n129));
  aoi022aa1n06x5               g034(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n130));
  nor042aa1n02x5               g035(.a(\b[4] ), .b(\a[5] ), .o1(new_n131));
  nona23aa1n02x4               g036(.a(new_n130), .b(new_n113), .c(new_n117), .d(new_n131), .out0(new_n132));
  norb02aa1n03x5               g037(.a(new_n110), .b(new_n132), .out0(new_n133));
  nanp02aa1n02x5               g038(.a(new_n133), .b(new_n129), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n123), .o1(new_n135));
  xnrc02aa1n02x5               g040(.a(\b[8] ), .b(\a[9] ), .out0(new_n136));
  aoai13aa1n02x5               g041(.a(new_n135), .b(new_n136), .c(new_n134), .d(new_n121), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n125), .b(new_n97), .c(new_n137), .o1(\s[10] ));
  aoai13aa1n06x5               g043(.a(new_n97), .b(new_n123), .c(new_n122), .d(new_n124), .o1(new_n139));
  tech160nm_fioaoi03aa1n02p5x5 g044(.a(\a[10] ), .b(\b[9] ), .c(new_n135), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  nor002aa1n16x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand42aa1n06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n139), .c(new_n141), .out0(\s[11] ));
  aoai13aa1n06x5               g050(.a(new_n144), .b(new_n140), .c(new_n137), .d(new_n97), .o1(new_n146));
  nor042aa1n09x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanp02aa1n12x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(\a[11] ), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\b[10] ), .o1(new_n151));
  aboi22aa1n03x5               g056(.a(new_n147), .b(new_n148), .c(new_n150), .d(new_n151), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n142), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n144), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n153), .b(new_n154), .c(new_n139), .d(new_n141), .o1(new_n155));
  aoi022aa1n02x5               g060(.a(new_n155), .b(new_n149), .c(new_n146), .d(new_n152), .o1(\s[12] ));
  norb03aa1n02x5               g061(.a(new_n119), .b(new_n131), .c(new_n117), .out0(new_n157));
  nona23aa1n02x4               g062(.a(new_n113), .b(new_n109), .c(new_n107), .d(new_n108), .out0(new_n158));
  oabi12aa1n03x5               g063(.a(new_n116), .b(new_n158), .c(new_n157), .out0(new_n159));
  xnrc02aa1n02x5               g064(.a(\b[9] ), .b(\a[10] ), .out0(new_n160));
  nona23aa1n06x5               g065(.a(new_n148), .b(new_n143), .c(new_n142), .d(new_n147), .out0(new_n161));
  nor043aa1n02x5               g066(.a(new_n161), .b(new_n160), .c(new_n136), .o1(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n159), .c(new_n133), .d(new_n129), .o1(new_n163));
  nano23aa1n02x4               g068(.a(new_n142), .b(new_n147), .c(new_n148), .d(new_n143), .out0(new_n164));
  nand23aa1n02x5               g069(.a(new_n164), .b(new_n124), .c(new_n97), .o1(new_n165));
  nand42aa1n16x5               g070(.a(\b[9] ), .b(\a[10] ), .o1(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  oai022aa1d18x5               g072(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n168));
  nor022aa1n04x5               g073(.a(new_n168), .b(new_n167), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n148), .b(new_n147), .c(new_n150), .d(new_n151), .o1(new_n170));
  oai012aa1d24x5               g075(.a(new_n166), .b(\b[10] ), .c(\a[11] ), .o1(new_n171));
  nanb03aa1d24x5               g076(.a(new_n147), .b(new_n148), .c(new_n143), .out0(new_n172));
  oai013aa1d12x5               g077(.a(new_n170), .b(new_n169), .c(new_n172), .d(new_n171), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n165), .c(new_n134), .d(new_n121), .o1(new_n175));
  nor042aa1n06x5               g080(.a(\b[12] ), .b(\a[13] ), .o1(new_n176));
  nand42aa1n03x5               g081(.a(\b[12] ), .b(\a[13] ), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  inv000aa1d42x5               g083(.a(new_n171), .o1(new_n179));
  nano22aa1n02x4               g084(.a(new_n147), .b(new_n143), .c(new_n148), .out0(new_n180));
  oai112aa1n03x5               g085(.a(new_n180), .b(new_n179), .c(new_n168), .d(new_n167), .o1(new_n181));
  nano22aa1n02x4               g086(.a(new_n178), .b(new_n181), .c(new_n170), .out0(new_n182));
  aoi022aa1n02x5               g087(.a(new_n175), .b(new_n178), .c(new_n163), .d(new_n182), .o1(\s[13] ));
  inv000aa1n02x5               g088(.a(new_n176), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n178), .b(new_n173), .c(new_n122), .d(new_n162), .o1(new_n185));
  nor002aa1n03x5               g090(.a(\b[13] ), .b(\a[14] ), .o1(new_n186));
  nanp02aa1n04x5               g091(.a(\b[13] ), .b(\a[14] ), .o1(new_n187));
  norb02aa1n02x5               g092(.a(new_n187), .b(new_n186), .out0(new_n188));
  xnbna2aa1n03x5               g093(.a(new_n188), .b(new_n185), .c(new_n184), .out0(\s[14] ));
  tech160nm_fioaoi03aa1n02p5x5 g094(.a(\a[14] ), .b(\b[13] ), .c(new_n184), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n190), .o1(new_n191));
  nano23aa1n06x5               g096(.a(new_n176), .b(new_n186), .c(new_n187), .d(new_n177), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n173), .c(new_n122), .d(new_n162), .o1(new_n193));
  nor002aa1d32x5               g098(.a(\b[14] ), .b(\a[15] ), .o1(new_n194));
  nand42aa1n08x5               g099(.a(\b[14] ), .b(\a[15] ), .o1(new_n195));
  norb02aa1n12x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n193), .c(new_n191), .out0(\s[15] ));
  aoai13aa1n02x5               g102(.a(new_n196), .b(new_n190), .c(new_n175), .d(new_n192), .o1(new_n198));
  xorc02aa1n02x5               g103(.a(\a[16] ), .b(\b[15] ), .out0(new_n199));
  inv000aa1d42x5               g104(.a(\a[16] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[15] ), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(new_n201), .b(new_n200), .o1(new_n202));
  and002aa1n18x5               g107(.a(\b[15] ), .b(\a[16] ), .o(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoi012aa1n02x5               g109(.a(new_n194), .b(new_n202), .c(new_n204), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n194), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n196), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n206), .b(new_n207), .c(new_n193), .d(new_n191), .o1(new_n208));
  aoi022aa1n02x5               g113(.a(new_n208), .b(new_n199), .c(new_n198), .d(new_n205), .o1(\s[16] ));
  aoi012aa1n06x5               g114(.a(new_n159), .b(new_n133), .c(new_n129), .o1(new_n210));
  nona23aa1n02x4               g115(.a(new_n187), .b(new_n177), .c(new_n176), .d(new_n186), .out0(new_n211));
  nano32aa1n03x7               g116(.a(new_n211), .b(new_n204), .c(new_n196), .d(new_n202), .out0(new_n212));
  nand22aa1n03x5               g117(.a(new_n212), .b(new_n162), .o1(new_n213));
  oai022aa1n02x5               g118(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n214));
  oaib12aa1n02x5               g119(.a(new_n214), .b(new_n201), .c(\a[16] ), .out0(new_n215));
  nona22aa1n02x4               g120(.a(new_n187), .b(new_n186), .c(new_n176), .out0(new_n216));
  oai012aa1n02x5               g121(.a(new_n187), .b(\b[14] ), .c(\a[15] ), .o1(new_n217));
  oai012aa1n02x5               g122(.a(new_n195), .b(\b[15] ), .c(\a[16] ), .o1(new_n218));
  nor003aa1n02x5               g123(.a(new_n218), .b(new_n217), .c(new_n203), .o1(new_n219));
  nanp02aa1n02x5               g124(.a(new_n219), .b(new_n216), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(new_n220), .b(new_n215), .o1(new_n221));
  tech160nm_fiaoi012aa1n05x5   g126(.a(new_n221), .b(new_n173), .c(new_n212), .o1(new_n222));
  oai012aa1n12x5               g127(.a(new_n222), .b(new_n210), .c(new_n213), .o1(new_n223));
  xorc02aa1n02x5               g128(.a(\a[17] ), .b(\b[16] ), .out0(new_n224));
  nanp03aa1n03x5               g129(.a(new_n192), .b(new_n196), .c(new_n199), .o1(new_n225));
  nor042aa1n04x5               g130(.a(new_n225), .b(new_n165), .o1(new_n226));
  nanb03aa1n02x5               g131(.a(new_n224), .b(new_n220), .c(new_n215), .out0(new_n227));
  aoi122aa1n02x5               g132(.a(new_n227), .b(new_n173), .c(new_n212), .d(new_n122), .e(new_n226), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n223), .c(new_n224), .o1(\s[17] ));
  inv000aa1d42x5               g134(.a(\a[17] ), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(\b[16] ), .b(new_n230), .out0(new_n231));
  aoi022aa1n02x5               g136(.a(new_n219), .b(new_n216), .c(new_n204), .d(new_n214), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n225), .c(new_n181), .d(new_n170), .o1(new_n233));
  aoai13aa1n06x5               g138(.a(new_n224), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n234));
  xorc02aa1n02x5               g139(.a(\a[18] ), .b(\b[17] ), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n234), .c(new_n231), .out0(\s[18] ));
  inv000aa1d42x5               g141(.a(\a[18] ), .o1(new_n237));
  xroi22aa1d04x5               g142(.a(new_n230), .b(\b[16] ), .c(new_n237), .d(\b[17] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n239));
  oaoi03aa1n02x5               g144(.a(\a[18] ), .b(\b[17] ), .c(new_n231), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  nor022aa1n16x5               g146(.a(\b[18] ), .b(\a[19] ), .o1(new_n242));
  nanp02aa1n04x5               g147(.a(\b[18] ), .b(\a[19] ), .o1(new_n243));
  norb02aa1n02x7               g148(.a(new_n243), .b(new_n242), .out0(new_n244));
  xnbna2aa1n03x5               g149(.a(new_n244), .b(new_n239), .c(new_n241), .out0(\s[19] ));
  xnrc02aa1n02x5               g150(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g151(.a(new_n244), .b(new_n240), .c(new_n223), .d(new_n238), .o1(new_n247));
  nor042aa1n04x5               g152(.a(\b[19] ), .b(\a[20] ), .o1(new_n248));
  nanp02aa1n06x5               g153(.a(\b[19] ), .b(\a[20] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  inv000aa1d42x5               g155(.a(\a[19] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\b[18] ), .o1(new_n252));
  aboi22aa1n03x5               g157(.a(new_n248), .b(new_n249), .c(new_n251), .d(new_n252), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n242), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n244), .o1(new_n255));
  aoai13aa1n02x5               g160(.a(new_n254), .b(new_n255), .c(new_n239), .d(new_n241), .o1(new_n256));
  aoi022aa1n02x5               g161(.a(new_n256), .b(new_n250), .c(new_n247), .d(new_n253), .o1(\s[20] ));
  nano23aa1n02x5               g162(.a(new_n242), .b(new_n248), .c(new_n249), .d(new_n243), .out0(new_n258));
  and003aa1n02x5               g163(.a(new_n258), .b(new_n235), .c(new_n224), .o(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n260));
  nanp02aa1n04x5               g165(.a(\b[17] ), .b(\a[18] ), .o1(new_n261));
  inv040aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  oai022aa1d18x5               g167(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n263));
  tech160nm_fiaoi012aa1n04x5   g168(.a(new_n242), .b(\a[18] ), .c(\b[17] ), .o1(new_n264));
  nano22aa1n03x7               g169(.a(new_n248), .b(new_n243), .c(new_n249), .out0(new_n265));
  oai112aa1n06x5               g170(.a(new_n265), .b(new_n264), .c(new_n263), .d(new_n262), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n249), .b(new_n248), .c(new_n251), .d(new_n252), .o1(new_n267));
  nand02aa1d10x5               g172(.a(new_n266), .b(new_n267), .o1(new_n268));
  nor022aa1n16x5               g173(.a(\b[20] ), .b(\a[21] ), .o1(new_n269));
  tech160nm_finand02aa1n03p5x5 g174(.a(\b[20] ), .b(\a[21] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n270), .b(new_n269), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n268), .c(new_n223), .d(new_n259), .o1(new_n272));
  nanb03aa1n02x5               g177(.a(new_n248), .b(new_n249), .c(new_n243), .out0(new_n273));
  nano32aa1n02x4               g178(.a(new_n273), .b(new_n263), .c(new_n254), .d(new_n261), .out0(new_n274));
  inv000aa1d42x5               g179(.a(new_n271), .o1(new_n275));
  nano22aa1n02x4               g180(.a(new_n274), .b(new_n267), .c(new_n275), .out0(new_n276));
  aobi12aa1n02x7               g181(.a(new_n272), .b(new_n276), .c(new_n260), .out0(\s[21] ));
  nor002aa1d32x5               g182(.a(\b[21] ), .b(\a[22] ), .o1(new_n278));
  nand42aa1d28x5               g183(.a(\b[21] ), .b(\a[22] ), .o1(new_n279));
  norb02aa1n02x5               g184(.a(new_n279), .b(new_n278), .out0(new_n280));
  inv040aa1n09x5               g185(.a(new_n278), .o1(new_n281));
  aoi012aa1n02x5               g186(.a(new_n269), .b(new_n281), .c(new_n279), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n268), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n269), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n275), .c(new_n260), .d(new_n283), .o1(new_n285));
  aoi022aa1n02x5               g190(.a(new_n285), .b(new_n280), .c(new_n272), .d(new_n282), .o1(\s[22] ));
  nona23aa1n02x4               g191(.a(new_n279), .b(new_n270), .c(new_n269), .d(new_n278), .out0(new_n287));
  nano32aa1n03x7               g192(.a(new_n287), .b(new_n258), .c(new_n235), .d(new_n224), .out0(new_n288));
  aoai13aa1n04x5               g193(.a(new_n288), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n289));
  nano23aa1n09x5               g194(.a(new_n269), .b(new_n278), .c(new_n279), .d(new_n270), .out0(new_n290));
  oai112aa1n06x5               g195(.a(new_n281), .b(new_n279), .c(\b[20] ), .d(\a[21] ), .o1(new_n291));
  aoi022aa1n12x5               g196(.a(new_n268), .b(new_n290), .c(new_n279), .d(new_n291), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[23] ), .b(\b[22] ), .out0(new_n294));
  aoai13aa1n06x5               g199(.a(new_n294), .b(new_n293), .c(new_n223), .d(new_n288), .o1(new_n295));
  aoi122aa1n02x5               g200(.a(new_n294), .b(new_n279), .c(new_n291), .d(new_n268), .e(new_n290), .o1(new_n296));
  aobi12aa1n02x5               g201(.a(new_n295), .b(new_n296), .c(new_n289), .out0(\s[23] ));
  tech160nm_fixorc02aa1n02p5x5 g202(.a(\a[24] ), .b(\b[23] ), .out0(new_n298));
  inv040aa1d32x5               g203(.a(\a[23] ), .o1(new_n299));
  inv000aa1d42x5               g204(.a(\b[22] ), .o1(new_n300));
  aoi012aa1n02x5               g205(.a(new_n298), .b(new_n299), .c(new_n300), .o1(new_n301));
  nanp02aa1n02x5               g206(.a(new_n300), .b(new_n299), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n294), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n302), .b(new_n303), .c(new_n289), .d(new_n292), .o1(new_n304));
  aoi022aa1n02x5               g209(.a(new_n304), .b(new_n298), .c(new_n295), .d(new_n301), .o1(\s[24] ));
  nand23aa1n04x5               g210(.a(new_n290), .b(new_n294), .c(new_n298), .o1(new_n306));
  nano32aa1n02x4               g211(.a(new_n306), .b(new_n258), .c(new_n235), .d(new_n224), .out0(new_n307));
  and002aa1n02x5               g212(.a(\b[23] ), .b(\a[24] ), .o(new_n308));
  tech160nm_fioai012aa1n04x5   g213(.a(new_n279), .b(\b[22] ), .c(\a[23] ), .o1(new_n309));
  nanp02aa1n02x5               g214(.a(\b[22] ), .b(\a[23] ), .o1(new_n310));
  oai012aa1n02x5               g215(.a(new_n310), .b(\b[23] ), .c(\a[24] ), .o1(new_n311));
  nor043aa1n02x5               g216(.a(new_n311), .b(new_n309), .c(new_n308), .o1(new_n312));
  tech160nm_fioaoi03aa1n04x5   g217(.a(\a[24] ), .b(\b[23] ), .c(new_n302), .o1(new_n313));
  aoi012aa1n12x5               g218(.a(new_n313), .b(new_n312), .c(new_n291), .o1(new_n314));
  aoai13aa1n12x5               g219(.a(new_n314), .b(new_n306), .c(new_n266), .d(new_n267), .o1(new_n315));
  xorc02aa1n12x5               g220(.a(\a[25] ), .b(\b[24] ), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n223), .d(new_n307), .o1(new_n317));
  aoai13aa1n06x5               g222(.a(new_n307), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n318));
  nano22aa1n03x5               g223(.a(new_n287), .b(new_n294), .c(new_n298), .out0(new_n319));
  oaib12aa1n09x5               g224(.a(new_n319), .b(new_n274), .c(new_n267), .out0(new_n320));
  aoi112aa1n02x5               g225(.a(new_n313), .b(new_n316), .c(new_n312), .d(new_n291), .o1(new_n321));
  and003aa1n03x5               g226(.a(new_n318), .b(new_n321), .c(new_n320), .o(new_n322));
  norb02aa1n03x4               g227(.a(new_n317), .b(new_n322), .out0(\s[25] ));
  xorc02aa1n02x5               g228(.a(\a[26] ), .b(\b[25] ), .out0(new_n324));
  nor042aa1n06x5               g229(.a(\b[24] ), .b(\a[25] ), .o1(new_n325));
  norp02aa1n02x5               g230(.a(new_n324), .b(new_n325), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n315), .o1(new_n327));
  inv000aa1n06x5               g232(.a(new_n325), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n316), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n328), .b(new_n329), .c(new_n318), .d(new_n327), .o1(new_n330));
  aoi022aa1n03x5               g235(.a(new_n330), .b(new_n324), .c(new_n317), .d(new_n326), .o1(\s[26] ));
  nanp02aa1n02x5               g236(.a(\b[24] ), .b(\a[25] ), .o1(new_n332));
  xnrc02aa1n02x5               g237(.a(\b[25] ), .b(\a[26] ), .out0(new_n333));
  nano22aa1n06x5               g238(.a(new_n333), .b(new_n328), .c(new_n332), .out0(new_n334));
  nano32aa1n03x7               g239(.a(new_n306), .b(new_n238), .c(new_n334), .d(new_n258), .out0(new_n335));
  aoai13aa1n06x5               g240(.a(new_n335), .b(new_n233), .c(new_n122), .d(new_n226), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n334), .o1(new_n337));
  oaoi03aa1n02x5               g242(.a(\a[26] ), .b(\b[25] ), .c(new_n328), .o1(new_n338));
  inv000aa1n02x5               g243(.a(new_n338), .o1(new_n339));
  aoai13aa1n04x5               g244(.a(new_n339), .b(new_n337), .c(new_n320), .d(new_n314), .o1(new_n340));
  xorc02aa1n12x5               g245(.a(\a[27] ), .b(\b[26] ), .out0(new_n341));
  aoai13aa1n06x5               g246(.a(new_n341), .b(new_n340), .c(new_n223), .d(new_n335), .o1(new_n342));
  aoi112aa1n02x5               g247(.a(new_n341), .b(new_n338), .c(new_n315), .d(new_n334), .o1(new_n343));
  aobi12aa1n02x5               g248(.a(new_n342), .b(new_n343), .c(new_n336), .out0(\s[27] ));
  xorc02aa1n02x5               g249(.a(\a[28] ), .b(\b[27] ), .out0(new_n345));
  norp02aa1n02x5               g250(.a(\b[26] ), .b(\a[27] ), .o1(new_n346));
  norp02aa1n02x5               g251(.a(new_n345), .b(new_n346), .o1(new_n347));
  aoi012aa1n09x5               g252(.a(new_n338), .b(new_n315), .c(new_n334), .o1(new_n348));
  inv000aa1n03x5               g253(.a(new_n346), .o1(new_n349));
  inv000aa1n02x5               g254(.a(new_n341), .o1(new_n350));
  aoai13aa1n03x5               g255(.a(new_n349), .b(new_n350), .c(new_n336), .d(new_n348), .o1(new_n351));
  aoi022aa1n03x5               g256(.a(new_n351), .b(new_n345), .c(new_n342), .d(new_n347), .o1(\s[28] ));
  and002aa1n02x5               g257(.a(new_n345), .b(new_n341), .o(new_n353));
  aoai13aa1n02x5               g258(.a(new_n353), .b(new_n340), .c(new_n223), .d(new_n335), .o1(new_n354));
  inv000aa1d42x5               g259(.a(new_n353), .o1(new_n355));
  oao003aa1n02x5               g260(.a(\a[28] ), .b(\b[27] ), .c(new_n349), .carry(new_n356));
  aoai13aa1n03x5               g261(.a(new_n356), .b(new_n355), .c(new_n336), .d(new_n348), .o1(new_n357));
  xorc02aa1n02x5               g262(.a(\a[29] ), .b(\b[28] ), .out0(new_n358));
  norb02aa1n02x5               g263(.a(new_n356), .b(new_n358), .out0(new_n359));
  aoi022aa1n03x5               g264(.a(new_n357), .b(new_n358), .c(new_n354), .d(new_n359), .o1(\s[29] ));
  nanp02aa1n02x5               g265(.a(\b[0] ), .b(\a[1] ), .o1(new_n361));
  xorb03aa1n02x5               g266(.a(new_n361), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g267(.a(new_n350), .b(new_n345), .c(new_n358), .out0(new_n363));
  aoai13aa1n04x5               g268(.a(new_n363), .b(new_n340), .c(new_n223), .d(new_n335), .o1(new_n364));
  inv000aa1n02x5               g269(.a(new_n363), .o1(new_n365));
  inv000aa1d42x5               g270(.a(\b[28] ), .o1(new_n366));
  inv000aa1d42x5               g271(.a(\a[29] ), .o1(new_n367));
  oaib12aa1n02x5               g272(.a(new_n356), .b(\b[28] ), .c(new_n367), .out0(new_n368));
  oaib12aa1n02x5               g273(.a(new_n368), .b(new_n366), .c(\a[29] ), .out0(new_n369));
  aoai13aa1n03x5               g274(.a(new_n369), .b(new_n365), .c(new_n336), .d(new_n348), .o1(new_n370));
  xorc02aa1n02x5               g275(.a(\a[30] ), .b(\b[29] ), .out0(new_n371));
  oaoi13aa1n02x5               g276(.a(new_n371), .b(new_n368), .c(new_n367), .d(new_n366), .o1(new_n372));
  aoi022aa1n03x5               g277(.a(new_n370), .b(new_n371), .c(new_n364), .d(new_n372), .o1(\s[30] ));
  nano32aa1n03x7               g278(.a(new_n350), .b(new_n371), .c(new_n345), .d(new_n358), .out0(new_n374));
  aoai13aa1n02x5               g279(.a(new_n374), .b(new_n340), .c(new_n223), .d(new_n335), .o1(new_n375));
  aoi022aa1n02x5               g280(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n376));
  norb02aa1n02x5               g281(.a(\b[30] ), .b(\a[31] ), .out0(new_n377));
  obai22aa1n02x7               g282(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n378));
  aoi112aa1n02x5               g283(.a(new_n378), .b(new_n377), .c(new_n368), .d(new_n376), .o1(new_n379));
  inv000aa1d42x5               g284(.a(new_n374), .o1(new_n380));
  norp02aa1n02x5               g285(.a(\b[29] ), .b(\a[30] ), .o1(new_n381));
  aoi012aa1n02x5               g286(.a(new_n381), .b(new_n368), .c(new_n376), .o1(new_n382));
  aoai13aa1n03x5               g287(.a(new_n382), .b(new_n380), .c(new_n336), .d(new_n348), .o1(new_n383));
  xorc02aa1n02x5               g288(.a(\a[31] ), .b(\b[30] ), .out0(new_n384));
  aoi022aa1n03x5               g289(.a(new_n383), .b(new_n384), .c(new_n379), .d(new_n375), .o1(\s[31] ));
  xobna2aa1n03x5               g290(.a(new_n102), .b(new_n99), .c(new_n98), .out0(\s[3] ));
  norb02aa1n02x5               g291(.a(new_n103), .b(new_n104), .out0(new_n387));
  aoi013aa1n02x4               g292(.a(new_n100), .b(new_n98), .c(new_n99), .d(new_n101), .o1(new_n388));
  oai012aa1n02x5               g293(.a(new_n129), .b(new_n388), .c(new_n387), .o1(\s[4] ));
  nona22aa1n02x4               g294(.a(new_n129), .b(new_n111), .c(new_n131), .out0(new_n390));
  xorc02aa1n02x5               g295(.a(\a[5] ), .b(\b[4] ), .out0(new_n391));
  aoi012aa1n02x5               g296(.a(new_n391), .b(new_n129), .c(new_n103), .o1(new_n392));
  norb02aa1n02x5               g297(.a(new_n390), .b(new_n392), .out0(\s[5] ));
  aoi012aa1n02x5               g298(.a(new_n131), .b(new_n129), .c(new_n130), .o1(new_n394));
  nanp02aa1n02x5               g299(.a(new_n390), .b(new_n157), .o1(new_n395));
  aoai13aa1n02x5               g300(.a(new_n395), .b(new_n394), .c(new_n118), .d(new_n119), .o1(\s[6] ));
  nanp02aa1n02x5               g301(.a(\b[6] ), .b(\a[7] ), .o1(new_n397));
  aoi022aa1n02x5               g302(.a(new_n395), .b(new_n119), .c(new_n115), .d(new_n397), .o1(new_n398));
  aoi013aa1n02x4               g303(.a(new_n398), .b(new_n395), .c(new_n113), .d(new_n115), .o1(\s[7] ));
  norb02aa1n02x5               g304(.a(new_n109), .b(new_n108), .out0(new_n400));
  nanp03aa1n02x5               g305(.a(new_n395), .b(new_n115), .c(new_n113), .o1(new_n401));
  xnbna2aa1n03x5               g306(.a(new_n400), .b(new_n401), .c(new_n115), .out0(\s[8] ));
  aoi113aa1n02x5               g307(.a(new_n116), .b(new_n124), .c(new_n120), .d(new_n110), .e(new_n113), .o1(new_n403));
  aoi022aa1n02x5               g308(.a(new_n122), .b(new_n124), .c(new_n134), .d(new_n403), .o1(\s[9] ));
endmodule


