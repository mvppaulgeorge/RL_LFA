// Benchmark "adder" written by ABC on Wed Jul 17 17:31:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n331,
    new_n334, new_n336, new_n337, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  tech160nm_finand02aa1n05x5   g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  norp02aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  tech160nm_fiao0012aa1n02p5x5 g005(.a(new_n98), .b(new_n100), .c(new_n99), .o(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand02aa1n02x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oao003aa1n02x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .carry(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano23aa1n02x4               g011(.a(new_n98), .b(new_n100), .c(new_n106), .d(new_n99), .out0(new_n107));
  aoi012aa1n03x5               g012(.a(new_n101), .b(new_n107), .c(new_n105), .o1(new_n108));
  tech160nm_finand02aa1n03p5x5 g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  norp02aa1n03x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  norp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nand42aa1n16x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nano23aa1n02x4               g017(.a(new_n111), .b(new_n110), .c(new_n112), .d(new_n109), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  tech160nm_fixnrc02aa1n04x5   g019(.a(\b[7] ), .b(\a[8] ), .out0(new_n115));
  nona22aa1n02x4               g020(.a(new_n113), .b(new_n114), .c(new_n115), .out0(new_n116));
  oai022aa1n02x5               g021(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  nanp03aa1n03x5               g022(.a(new_n117), .b(new_n109), .c(new_n112), .o1(new_n118));
  oab012aa1n03x5               g023(.a(new_n110), .b(\a[8] ), .c(\b[7] ), .out0(new_n119));
  aoi022aa1n12x5               g024(.a(new_n118), .b(new_n119), .c(\b[7] ), .d(\a[8] ), .o1(new_n120));
  inv000aa1n02x5               g025(.a(new_n120), .o1(new_n121));
  oai012aa1n02x5               g026(.a(new_n121), .b(new_n108), .c(new_n116), .o1(new_n122));
  nand42aa1n06x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  norb02aa1n02x5               g028(.a(new_n123), .b(new_n97), .out0(new_n124));
  nor042aa1n02x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nand02aa1n04x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  norb02aa1n06x4               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  aoai13aa1n03x5               g032(.a(new_n127), .b(new_n97), .c(new_n122), .d(new_n124), .o1(new_n128));
  aoi112aa1n02x5               g033(.a(new_n127), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n128), .b(new_n129), .out0(\s[10] ));
  tech160nm_fiaoi012aa1n04x5   g035(.a(new_n125), .b(new_n97), .c(new_n126), .o1(new_n131));
  nand42aa1n06x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nor042aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n06x4               g038(.a(new_n132), .b(new_n133), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n128), .c(new_n131), .out0(\s[11] ));
  and002aa1n02x5               g040(.a(new_n131), .b(new_n134), .o(new_n136));
  nanp02aa1n02x5               g041(.a(new_n128), .b(new_n136), .o1(new_n137));
  nor042aa1n03x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoi012aa1n02x5               g045(.a(new_n140), .b(new_n137), .c(new_n132), .o1(new_n141));
  nanp03aa1n02x5               g046(.a(new_n137), .b(new_n132), .c(new_n140), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(\s[12] ));
  oaoi03aa1n02x5               g048(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n144));
  nona23aa1n02x4               g049(.a(new_n106), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n145));
  oabi12aa1n09x5               g050(.a(new_n101), .b(new_n145), .c(new_n144), .out0(new_n146));
  norb02aa1n02x5               g051(.a(new_n109), .b(new_n110), .out0(new_n147));
  norb02aa1n06x4               g052(.a(new_n112), .b(new_n111), .out0(new_n148));
  nano23aa1n06x5               g053(.a(new_n115), .b(new_n114), .c(new_n148), .d(new_n147), .out0(new_n149));
  nona23aa1n03x5               g054(.a(new_n132), .b(new_n139), .c(new_n138), .d(new_n133), .out0(new_n150));
  nano22aa1n03x7               g055(.a(new_n150), .b(new_n124), .c(new_n127), .out0(new_n151));
  aoai13aa1n03x5               g056(.a(new_n151), .b(new_n120), .c(new_n149), .d(new_n146), .o1(new_n152));
  inv030aa1n06x5               g057(.a(new_n131), .o1(new_n153));
  nano23aa1n03x7               g058(.a(new_n138), .b(new_n133), .c(new_n139), .d(new_n132), .out0(new_n154));
  aoi012aa1n02x5               g059(.a(new_n138), .b(new_n133), .c(new_n139), .o1(new_n155));
  inv000aa1n02x5               g060(.a(new_n155), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n156), .b(new_n154), .c(new_n153), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(new_n152), .b(new_n157), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nand42aa1n02x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nor002aa1n02x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n161), .b(new_n158), .c(new_n160), .o1(new_n162));
  xnrb03aa1n02x5               g067(.a(new_n162), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nand02aa1n03x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n160), .b(new_n165), .c(new_n164), .d(new_n161), .out0(new_n166));
  aoi012aa1n02x5               g071(.a(new_n164), .b(new_n161), .c(new_n165), .o1(new_n167));
  aoai13aa1n03x5               g072(.a(new_n167), .b(new_n166), .c(new_n152), .d(new_n157), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand42aa1n03x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nor022aa1n03x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norp02aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand42aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  aoai13aa1n02x5               g080(.a(new_n175), .b(new_n171), .c(new_n168), .d(new_n170), .o1(new_n176));
  aoi112aa1n02x5               g081(.a(new_n175), .b(new_n171), .c(new_n168), .d(new_n170), .o1(new_n177));
  nanb02aa1n03x5               g082(.a(new_n177), .b(new_n176), .out0(\s[16] ));
  nano23aa1n06x5               g083(.a(new_n164), .b(new_n161), .c(new_n165), .d(new_n160), .out0(new_n179));
  nano23aa1n03x5               g084(.a(new_n172), .b(new_n171), .c(new_n173), .d(new_n170), .out0(new_n180));
  nanp02aa1n02x5               g085(.a(new_n180), .b(new_n179), .o1(new_n181));
  nano32aa1n03x7               g086(.a(new_n181), .b(new_n154), .c(new_n127), .d(new_n124), .out0(new_n182));
  aoai13aa1n06x5               g087(.a(new_n182), .b(new_n120), .c(new_n149), .d(new_n146), .o1(new_n183));
  aoi112aa1n02x5               g088(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n184));
  oai112aa1n03x5               g089(.a(new_n134), .b(new_n140), .c(new_n184), .d(new_n125), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n167), .b(new_n166), .c(new_n185), .d(new_n155), .o1(new_n186));
  nand42aa1n02x5               g091(.a(new_n186), .b(new_n180), .o1(new_n187));
  oai012aa1n02x5               g092(.a(new_n173), .b(new_n172), .c(new_n171), .o1(new_n188));
  nand23aa1n06x5               g093(.a(new_n183), .b(new_n187), .c(new_n188), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g095(.a(\a[18] ), .o1(new_n191));
  inv040aa1d32x5               g096(.a(\a[17] ), .o1(new_n192));
  inv030aa1d32x5               g097(.a(\b[16] ), .o1(new_n193));
  oaoi03aa1n03x5               g098(.a(new_n192), .b(new_n193), .c(new_n189), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[17] ), .c(new_n191), .out0(\s[18] ));
  aobi12aa1n06x5               g100(.a(new_n188), .b(new_n186), .c(new_n180), .out0(new_n196));
  xroi22aa1d06x4               g101(.a(new_n192), .b(\b[16] ), .c(new_n191), .d(\b[17] ), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  oai022aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n199));
  oaib12aa1n03x5               g104(.a(new_n199), .b(new_n191), .c(\b[17] ), .out0(new_n200));
  aoai13aa1n03x5               g105(.a(new_n200), .b(new_n198), .c(new_n196), .d(new_n183), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nand42aa1n06x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  nor002aa1n20x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand42aa1n08x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n204), .c(new_n201), .d(new_n207), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(new_n193), .b(new_n192), .o1(new_n212));
  oaoi03aa1n09x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n212), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n207), .b(new_n213), .c(new_n189), .d(new_n197), .o1(new_n214));
  nona22aa1n03x5               g119(.a(new_n214), .b(new_n210), .c(new_n204), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n211), .b(new_n215), .o1(\s[20] ));
  nano23aa1d12x5               g121(.a(new_n208), .b(new_n204), .c(new_n209), .d(new_n205), .out0(new_n217));
  nand22aa1n09x5               g122(.a(new_n197), .b(new_n217), .o1(new_n218));
  nona23aa1n03x5               g123(.a(new_n205), .b(new_n209), .c(new_n208), .d(new_n204), .out0(new_n219));
  oa0012aa1n12x5               g124(.a(new_n209), .b(new_n208), .c(new_n204), .o(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  oai012aa1n09x5               g126(.a(new_n221), .b(new_n219), .c(new_n200), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n218), .c(new_n196), .d(new_n183), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  tech160nm_fixnrc02aa1n04x5   g133(.a(\b[21] ), .b(\a[22] ), .out0(new_n229));
  aoai13aa1n02x5               g134(.a(new_n229), .b(new_n226), .c(new_n224), .d(new_n228), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n218), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n228), .b(new_n222), .c(new_n189), .d(new_n231), .o1(new_n232));
  nona22aa1n02x4               g137(.a(new_n232), .b(new_n229), .c(new_n226), .out0(new_n233));
  nanp02aa1n02x5               g138(.a(new_n230), .b(new_n233), .o1(\s[22] ));
  nona23aa1n03x5               g139(.a(new_n170), .b(new_n173), .c(new_n172), .d(new_n171), .out0(new_n235));
  nona22aa1n03x5               g140(.a(new_n151), .b(new_n166), .c(new_n235), .out0(new_n236));
  oaoi13aa1n06x5               g141(.a(new_n236), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n179), .b(new_n156), .c(new_n154), .d(new_n153), .o1(new_n238));
  aoai13aa1n06x5               g143(.a(new_n188), .b(new_n235), .c(new_n238), .d(new_n167), .o1(new_n239));
  nor042aa1n09x5               g144(.a(new_n229), .b(new_n227), .o1(new_n240));
  nano22aa1n02x4               g145(.a(new_n198), .b(new_n240), .c(new_n217), .out0(new_n241));
  tech160nm_fioai012aa1n05x5   g146(.a(new_n241), .b(new_n239), .c(new_n237), .o1(new_n242));
  aoai13aa1n12x5               g147(.a(new_n240), .b(new_n220), .c(new_n217), .d(new_n213), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  inv000aa1d42x5               g149(.a(\a[22] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\b[21] ), .o1(new_n246));
  oao003aa1n02x5               g151(.a(new_n245), .b(new_n246), .c(new_n226), .carry(new_n247));
  nona22aa1n02x4               g152(.a(new_n242), .b(new_n244), .c(new_n247), .out0(new_n248));
  nor042aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  and002aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .o(new_n250));
  norp02aa1n03x5               g155(.a(new_n250), .b(new_n249), .o1(new_n251));
  nona32aa1n02x4               g156(.a(new_n242), .b(new_n251), .c(new_n247), .d(new_n244), .out0(new_n252));
  aobi12aa1n02x5               g157(.a(new_n252), .b(new_n251), .c(new_n248), .out0(\s[23] ));
  norp02aa1n02x5               g158(.a(new_n247), .b(new_n249), .o1(new_n254));
  aoi013aa1n02x4               g159(.a(new_n250), .b(new_n242), .c(new_n243), .d(new_n254), .o1(new_n255));
  xnrc02aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .out0(new_n256));
  nona32aa1n03x5               g161(.a(new_n242), .b(new_n249), .c(new_n247), .d(new_n244), .out0(new_n257));
  nanb03aa1n03x5               g162(.a(new_n250), .b(new_n257), .c(new_n256), .out0(new_n258));
  oaih12aa1n02x5               g163(.a(new_n258), .b(new_n255), .c(new_n256), .o1(\s[24] ));
  norb02aa1n03x5               g164(.a(new_n251), .b(new_n256), .out0(new_n260));
  nano22aa1n06x5               g165(.a(new_n218), .b(new_n240), .c(new_n260), .out0(new_n261));
  inv020aa1n03x5               g166(.a(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n247), .o1(new_n263));
  inv000aa1n02x5               g168(.a(new_n260), .o1(new_n264));
  inv000aa1d42x5               g169(.a(\a[24] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(\b[23] ), .o1(new_n266));
  oao003aa1n02x5               g171(.a(new_n265), .b(new_n266), .c(new_n249), .carry(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n12x5               g173(.a(new_n268), .b(new_n264), .c(new_n243), .d(new_n263), .o1(new_n269));
  inv040aa1n03x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n262), .c(new_n196), .d(new_n183), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n276));
  aoai13aa1n02x5               g181(.a(new_n274), .b(new_n269), .c(new_n189), .d(new_n261), .o1(new_n277));
  nona22aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .out0(new_n278));
  nanp02aa1n03x5               g183(.a(new_n276), .b(new_n278), .o1(\s[26] ));
  nor002aa1d32x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  and002aa1n24x5               g185(.a(\b[26] ), .b(\a[27] ), .o(new_n281));
  nor042aa1n06x5               g186(.a(new_n281), .b(new_n280), .o1(new_n282));
  norb02aa1n06x5               g187(.a(new_n274), .b(new_n275), .out0(new_n283));
  nano32aa1d12x5               g188(.a(new_n218), .b(new_n283), .c(new_n240), .d(new_n260), .out0(new_n284));
  oai012aa1n12x5               g189(.a(new_n284), .b(new_n239), .c(new_n237), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(\b[25] ), .b(\a[26] ), .o1(new_n286));
  oai022aa1n02x5               g191(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n287));
  aoi022aa1n12x5               g192(.a(new_n269), .b(new_n283), .c(new_n286), .d(new_n287), .o1(new_n288));
  xnbna2aa1n06x5               g193(.a(new_n282), .b(new_n285), .c(new_n288), .out0(\s[27] ));
  inv000aa1d42x5               g194(.a(new_n281), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n260), .b(new_n247), .c(new_n222), .d(new_n240), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n283), .o1(new_n292));
  nanp02aa1n02x5               g197(.a(new_n287), .b(new_n286), .o1(new_n293));
  aoai13aa1n04x5               g198(.a(new_n293), .b(new_n292), .c(new_n291), .d(new_n268), .o1(new_n294));
  aoai13aa1n02x5               g199(.a(new_n290), .b(new_n294), .c(new_n284), .d(new_n189), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .out0(new_n296));
  norp02aa1n02x5               g201(.a(new_n296), .b(new_n280), .o1(new_n297));
  inv040aa1n08x5               g202(.a(new_n280), .o1(new_n298));
  aoai13aa1n06x5               g203(.a(new_n298), .b(new_n281), .c(new_n285), .d(new_n288), .o1(new_n299));
  aoi022aa1n03x5               g204(.a(new_n299), .b(new_n296), .c(new_n295), .d(new_n297), .o1(\s[28] ));
  and002aa1n06x5               g205(.a(new_n296), .b(new_n282), .o(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n294), .c(new_n189), .d(new_n284), .o1(new_n302));
  inv000aa1n02x5               g207(.a(new_n301), .o1(new_n303));
  oao003aa1n03x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n298), .carry(new_n304));
  aoai13aa1n04x5               g209(.a(new_n304), .b(new_n303), .c(new_n285), .d(new_n288), .o1(new_n305));
  xorc02aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n304), .b(new_n306), .out0(new_n307));
  aoi022aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n302), .d(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g214(.a(new_n296), .b(new_n306), .c(new_n282), .o(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n294), .c(new_n189), .d(new_n284), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n310), .o1(new_n312));
  tech160nm_fioaoi03aa1n02p5x5 g217(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n313), .o1(new_n314));
  aoai13aa1n04x5               g219(.a(new_n314), .b(new_n312), .c(new_n285), .d(new_n288), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .out0(new_n316));
  norp02aa1n02x5               g221(.a(new_n313), .b(new_n316), .o1(new_n317));
  aoi022aa1n02x7               g222(.a(new_n315), .b(new_n316), .c(new_n311), .d(new_n317), .o1(\s[30] ));
  nano22aa1d15x5               g223(.a(new_n303), .b(new_n306), .c(new_n316), .out0(new_n319));
  aoai13aa1n02x5               g224(.a(new_n319), .b(new_n294), .c(new_n189), .d(new_n284), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n319), .o1(new_n321));
  inv000aa1d42x5               g226(.a(\a[30] ), .o1(new_n322));
  inv000aa1d42x5               g227(.a(\b[29] ), .o1(new_n323));
  oaoi03aa1n03x5               g228(.a(new_n322), .b(new_n323), .c(new_n313), .o1(new_n324));
  aoai13aa1n06x5               g229(.a(new_n324), .b(new_n321), .c(new_n285), .d(new_n288), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[31] ), .b(\b[30] ), .out0(new_n326));
  oabi12aa1n02x5               g231(.a(new_n326), .b(\a[30] ), .c(\b[29] ), .out0(new_n327));
  oaoi13aa1n04x5               g232(.a(new_n327), .b(new_n313), .c(new_n322), .d(new_n323), .o1(new_n328));
  aoi022aa1n03x5               g233(.a(new_n325), .b(new_n326), .c(new_n320), .d(new_n328), .o1(\s[31] ));
  xnrb03aa1n02x5               g234(.a(new_n144), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g235(.a(\a[3] ), .b(\b[2] ), .c(new_n144), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g237(.a(new_n146), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oao003aa1n02x5               g238(.a(\a[5] ), .b(\b[4] ), .c(new_n108), .carry(new_n334));
  xnrc02aa1n02x5               g239(.a(new_n334), .b(new_n148), .out0(\s[6] ));
  inv000aa1d42x5               g240(.a(new_n112), .o1(new_n336));
  aoai13aa1n02x5               g241(.a(new_n147), .b(new_n336), .c(new_n334), .d(new_n148), .o1(new_n337));
  aoi112aa1n02x5               g242(.a(new_n147), .b(new_n336), .c(new_n334), .d(new_n148), .o1(new_n338));
  nanb02aa1n02x5               g243(.a(new_n338), .b(new_n337), .out0(\s[7] ));
  xnbna2aa1n03x5               g244(.a(new_n115), .b(new_n337), .c(new_n109), .out0(\s[8] ));
  xorb03aa1n02x5               g245(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


