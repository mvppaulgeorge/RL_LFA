// Benchmark "adder" written by ABC on Wed Jul 17 14:56:02 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n316, new_n317,
    new_n320, new_n321, new_n322, new_n323, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand02aa1n03x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nanp02aa1n03x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  aoi012aa1n06x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor002aa1n12x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  tech160nm_finand02aa1n03p5x5 g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n09x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  tech160nm_fiaoi012aa1n03p5x5 g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  nand02aa1d16x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  inv000aa1n03x5               g019(.a(new_n114), .o1(new_n115));
  oai112aa1n03x5               g020(.a(new_n115), .b(new_n113), .c(\b[6] ), .d(\a[7] ), .o1(new_n116));
  tech160nm_finand02aa1n03p5x5 g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nor002aa1n04x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanp02aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor042aa1n04x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n119), .b(new_n117), .c(new_n120), .d(new_n118), .out0(new_n121));
  aoi112aa1n06x5               g026(.a(new_n121), .b(new_n116), .c(\a[7] ), .d(\b[6] ), .o1(new_n122));
  inv040aa1d32x5               g027(.a(\a[7] ), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\b[6] ), .o1(new_n124));
  nand42aa1n02x5               g029(.a(new_n124), .b(new_n123), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[8] ), .b(\b[7] ), .c(new_n125), .o1(new_n126));
  tech160nm_fixnrc02aa1n05x5   g031(.a(\b[6] ), .b(\a[7] ), .out0(new_n127));
  norb02aa1n12x5               g032(.a(new_n113), .b(new_n114), .out0(new_n128));
  oai112aa1n02x7               g033(.a(new_n128), .b(new_n119), .c(new_n120), .d(new_n118), .o1(new_n129));
  oabi12aa1n06x5               g034(.a(new_n126), .b(new_n129), .c(new_n127), .out0(new_n130));
  nanp02aa1n04x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nanb02aa1n18x5               g036(.a(new_n100), .b(new_n131), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n130), .c(new_n112), .d(new_n122), .o1(new_n134));
  xobna2aa1n03x5               g039(.a(new_n99), .b(new_n134), .c(new_n101), .out0(\s[10] ));
  norp02aa1n02x5               g040(.a(new_n100), .b(new_n97), .o1(new_n136));
  aoi022aa1n02x5               g041(.a(new_n134), .b(new_n136), .c(\b[9] ), .d(\a[10] ), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand02aa1n06x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n139), .b(new_n137), .c(new_n140), .o1(new_n141));
  xnrb03aa1n02x5               g046(.a(new_n141), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor022aa1n16x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand22aa1n12x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nona23aa1n09x5               g049(.a(new_n144), .b(new_n140), .c(new_n139), .d(new_n143), .out0(new_n145));
  nor043aa1n03x5               g050(.a(new_n145), .b(new_n132), .c(new_n99), .o1(new_n146));
  aoai13aa1n06x5               g051(.a(new_n146), .b(new_n130), .c(new_n112), .d(new_n122), .o1(new_n147));
  oai012aa1d24x5               g052(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n148));
  ao0012aa1n03x7               g053(.a(new_n143), .b(new_n139), .c(new_n144), .o(new_n149));
  oabi12aa1n18x5               g054(.a(new_n149), .b(new_n145), .c(new_n148), .out0(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[12] ), .b(\a[13] ), .out0(new_n152));
  xobna2aa1n03x5               g057(.a(new_n152), .b(new_n147), .c(new_n151), .out0(\s[13] ));
  orn002aa1n24x5               g058(.a(\a[13] ), .b(\b[12] ), .o(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n152), .c(new_n147), .d(new_n151), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nanp02aa1n03x5               g061(.a(new_n147), .b(new_n151), .o1(new_n157));
  tech160nm_fixnrc02aa1n02p5x5 g062(.a(\b[13] ), .b(\a[14] ), .out0(new_n158));
  nor042aa1n04x5               g063(.a(new_n158), .b(new_n152), .o1(new_n159));
  oaoi03aa1n12x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n154), .o1(new_n160));
  nor042aa1n03x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(new_n161), .b(new_n162), .out0(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n160), .c(new_n157), .d(new_n159), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n164), .b(new_n160), .c(new_n157), .d(new_n159), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(\s[15] ));
  nor042aa1n03x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  nanp02aa1n04x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nanb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(new_n170));
  oai112aa1n02x7               g075(.a(new_n165), .b(new_n170), .c(\b[14] ), .d(\a[15] ), .o1(new_n171));
  oaoi13aa1n06x5               g076(.a(new_n170), .b(new_n165), .c(\a[15] ), .d(\b[14] ), .o1(new_n172));
  norb02aa1n03x4               g077(.a(new_n171), .b(new_n172), .out0(\s[16] ));
  aoi012aa1n12x5               g078(.a(new_n130), .b(new_n112), .c(new_n122), .o1(new_n174));
  nano23aa1d15x5               g079(.a(new_n161), .b(new_n168), .c(new_n169), .d(new_n162), .out0(new_n175));
  nand23aa1n03x5               g080(.a(new_n146), .b(new_n159), .c(new_n175), .o1(new_n176));
  aoai13aa1n12x5               g081(.a(new_n175), .b(new_n160), .c(new_n150), .d(new_n159), .o1(new_n177));
  tech160nm_fiaoi012aa1n03p5x5 g082(.a(new_n168), .b(new_n161), .c(new_n169), .o1(new_n178));
  oai112aa1n06x5               g083(.a(new_n177), .b(new_n178), .c(new_n174), .d(new_n176), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  inv040aa1d32x5               g086(.a(\a[17] ), .o1(new_n182));
  inv030aa1d32x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n03x5               g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  nor042aa1n04x5               g090(.a(new_n174), .b(new_n176), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n160), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n175), .o1(new_n188));
  nano23aa1n06x5               g093(.a(new_n139), .b(new_n143), .c(new_n144), .d(new_n140), .out0(new_n189));
  inv040aa1n02x5               g094(.a(new_n148), .o1(new_n190));
  aoai13aa1n06x5               g095(.a(new_n159), .b(new_n149), .c(new_n189), .d(new_n190), .o1(new_n191));
  aoai13aa1n04x5               g096(.a(new_n178), .b(new_n188), .c(new_n191), .d(new_n187), .o1(new_n192));
  xroi22aa1d06x4               g097(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n193));
  tech160nm_fioai012aa1n03p5x5 g098(.a(new_n193), .b(new_n186), .c(new_n192), .o1(new_n194));
  oai022aa1n09x5               g099(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n195));
  oaib12aa1n06x5               g100(.a(new_n195), .b(new_n181), .c(\b[17] ), .out0(new_n196));
  nor002aa1d32x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nand42aa1d28x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nanb02aa1n02x5               g103(.a(new_n197), .b(new_n198), .out0(new_n199));
  inv000aa1d42x5               g104(.a(new_n199), .o1(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n200), .b(new_n194), .c(new_n196), .out0(\s[19] ));
  xnrc02aa1n02x5               g106(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g107(.a(new_n197), .o1(new_n203));
  tech160nm_fiaoi012aa1n03p5x5 g108(.a(new_n199), .b(new_n194), .c(new_n196), .o1(new_n204));
  nor042aa1n09x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand42aa1d28x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  nano22aa1n03x5               g112(.a(new_n204), .b(new_n203), .c(new_n207), .out0(new_n208));
  nand02aa1n03x5               g113(.a(new_n183), .b(new_n182), .o1(new_n209));
  oaoi03aa1n12x5               g114(.a(\a[18] ), .b(\b[17] ), .c(new_n209), .o1(new_n210));
  aoai13aa1n03x5               g115(.a(new_n200), .b(new_n210), .c(new_n179), .d(new_n193), .o1(new_n211));
  aoi012aa1n03x5               g116(.a(new_n207), .b(new_n211), .c(new_n203), .o1(new_n212));
  nor002aa1n02x5               g117(.a(new_n212), .b(new_n208), .o1(\s[20] ));
  nano23aa1n09x5               g118(.a(new_n197), .b(new_n205), .c(new_n206), .d(new_n198), .out0(new_n214));
  nand22aa1n03x5               g119(.a(new_n193), .b(new_n214), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  oai012aa1n03x5               g121(.a(new_n216), .b(new_n186), .c(new_n192), .o1(new_n217));
  nona23aa1d18x5               g122(.a(new_n206), .b(new_n198), .c(new_n197), .d(new_n205), .out0(new_n218));
  aoi012aa1n12x5               g123(.a(new_n205), .b(new_n197), .c(new_n206), .o1(new_n219));
  oai012aa1n18x5               g124(.a(new_n219), .b(new_n218), .c(new_n196), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  nor042aa1d18x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  nand42aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  xnbna2aa1n03x5               g129(.a(new_n224), .b(new_n217), .c(new_n221), .out0(\s[21] ));
  inv000aa1d42x5               g130(.a(new_n222), .o1(new_n226));
  aobi12aa1n02x5               g131(.a(new_n224), .b(new_n217), .c(new_n221), .out0(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  nano22aa1n02x4               g133(.a(new_n227), .b(new_n226), .c(new_n228), .out0(new_n229));
  aoai13aa1n03x5               g134(.a(new_n224), .b(new_n220), .c(new_n179), .d(new_n216), .o1(new_n230));
  aoi012aa1n03x5               g135(.a(new_n228), .b(new_n230), .c(new_n226), .o1(new_n231));
  nor002aa1n02x5               g136(.a(new_n231), .b(new_n229), .o1(\s[22] ));
  nano22aa1n12x5               g137(.a(new_n228), .b(new_n226), .c(new_n223), .out0(new_n233));
  and003aa1n02x5               g138(.a(new_n193), .b(new_n233), .c(new_n214), .o(new_n234));
  oai012aa1n03x5               g139(.a(new_n234), .b(new_n186), .c(new_n192), .o1(new_n235));
  oao003aa1n09x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n226), .carry(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi012aa1n02x5               g142(.a(new_n237), .b(new_n220), .c(new_n233), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[22] ), .b(\a[23] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  xnbna2aa1n03x5               g145(.a(new_n240), .b(new_n235), .c(new_n238), .out0(\s[23] ));
  nor042aa1n06x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n239), .b(new_n235), .c(new_n238), .o1(new_n244));
  xnrc02aa1n12x5               g149(.a(\b[23] ), .b(\a[24] ), .out0(new_n245));
  nano22aa1n02x4               g150(.a(new_n244), .b(new_n243), .c(new_n245), .out0(new_n246));
  inv000aa1n02x5               g151(.a(new_n238), .o1(new_n247));
  aoai13aa1n03x5               g152(.a(new_n240), .b(new_n247), .c(new_n179), .d(new_n234), .o1(new_n248));
  aoi012aa1n03x5               g153(.a(new_n245), .b(new_n248), .c(new_n243), .o1(new_n249));
  nor002aa1n02x5               g154(.a(new_n249), .b(new_n246), .o1(\s[24] ));
  norp02aa1n09x5               g155(.a(new_n245), .b(new_n239), .o1(new_n251));
  nano22aa1n03x7               g156(.a(new_n215), .b(new_n233), .c(new_n251), .out0(new_n252));
  oai012aa1n02x5               g157(.a(new_n252), .b(new_n186), .c(new_n192), .o1(new_n253));
  inv020aa1n04x5               g158(.a(new_n219), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n233), .b(new_n254), .c(new_n214), .d(new_n210), .o1(new_n255));
  inv000aa1n03x5               g160(.a(new_n251), .o1(new_n256));
  oao003aa1n02x5               g161(.a(\a[24] ), .b(\b[23] ), .c(new_n243), .carry(new_n257));
  aoai13aa1n12x5               g162(.a(new_n257), .b(new_n256), .c(new_n255), .d(new_n236), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[24] ), .b(\a[25] ), .out0(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n253), .c(new_n259), .out0(\s[25] ));
  nor042aa1n03x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aoi012aa1n02x7               g169(.a(new_n260), .b(new_n253), .c(new_n259), .o1(new_n265));
  xnrc02aa1n02x5               g170(.a(\b[25] ), .b(\a[26] ), .out0(new_n266));
  nano22aa1n02x5               g171(.a(new_n265), .b(new_n264), .c(new_n266), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n261), .b(new_n258), .c(new_n179), .d(new_n252), .o1(new_n268));
  aoi012aa1n03x5               g173(.a(new_n266), .b(new_n268), .c(new_n264), .o1(new_n269));
  nor002aa1n02x5               g174(.a(new_n269), .b(new_n267), .o1(\s[26] ));
  nor042aa1n06x5               g175(.a(new_n266), .b(new_n260), .o1(new_n271));
  nano32aa1n03x7               g176(.a(new_n215), .b(new_n271), .c(new_n233), .d(new_n251), .out0(new_n272));
  oai012aa1n06x5               g177(.a(new_n272), .b(new_n186), .c(new_n192), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .c(new_n264), .carry(new_n274));
  aobi12aa1n12x5               g179(.a(new_n274), .b(new_n258), .c(new_n271), .out0(new_n275));
  xorc02aa1n12x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n273), .c(new_n275), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  inv040aa1n03x5               g183(.a(new_n278), .o1(new_n279));
  aobi12aa1n06x5               g184(.a(new_n276), .b(new_n273), .c(new_n275), .out0(new_n280));
  xnrc02aa1n02x5               g185(.a(\b[27] ), .b(\a[28] ), .out0(new_n281));
  nano22aa1n03x7               g186(.a(new_n280), .b(new_n279), .c(new_n281), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n251), .b(new_n237), .c(new_n220), .d(new_n233), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n271), .o1(new_n284));
  aoai13aa1n04x5               g189(.a(new_n274), .b(new_n284), .c(new_n283), .d(new_n257), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n276), .b(new_n285), .c(new_n179), .d(new_n272), .o1(new_n286));
  aoi012aa1n02x5               g191(.a(new_n281), .b(new_n286), .c(new_n279), .o1(new_n287));
  norp02aa1n03x5               g192(.a(new_n287), .b(new_n282), .o1(\s[28] ));
  norb02aa1n02x5               g193(.a(new_n276), .b(new_n281), .out0(new_n289));
  aoai13aa1n02x7               g194(.a(new_n289), .b(new_n285), .c(new_n179), .d(new_n272), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n279), .carry(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[28] ), .b(\a[29] ), .out0(new_n292));
  aoi012aa1n02x7               g197(.a(new_n292), .b(new_n290), .c(new_n291), .o1(new_n293));
  aobi12aa1n06x5               g198(.a(new_n289), .b(new_n273), .c(new_n275), .out0(new_n294));
  nano22aa1n03x7               g199(.a(new_n294), .b(new_n291), .c(new_n292), .out0(new_n295));
  norp02aa1n03x5               g200(.a(new_n293), .b(new_n295), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g202(.a(new_n276), .b(new_n292), .c(new_n281), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n285), .c(new_n179), .d(new_n272), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[29] ), .b(\a[30] ), .out0(new_n301));
  aoi012aa1n02x5               g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  aobi12aa1n06x5               g207(.a(new_n298), .b(new_n273), .c(new_n275), .out0(new_n303));
  nano22aa1n03x7               g208(.a(new_n303), .b(new_n300), .c(new_n301), .out0(new_n304));
  norp02aa1n03x5               g209(.a(new_n302), .b(new_n304), .o1(\s[30] ));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n298), .b(new_n301), .out0(new_n307));
  aoai13aa1n02x7               g212(.a(new_n307), .b(new_n285), .c(new_n179), .d(new_n272), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  aobi12aa1n06x5               g215(.a(new_n307), .b(new_n273), .c(new_n275), .out0(new_n311));
  nano22aa1n03x7               g216(.a(new_n311), .b(new_n306), .c(new_n309), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n310), .b(new_n312), .o1(\s[31] ));
  xnrb03aa1n02x5               g218(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g219(.a(new_n106), .o1(new_n315));
  nona22aa1n02x4               g220(.a(new_n109), .b(new_n105), .c(new_n108), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n108), .b(new_n315), .c(new_n107), .o1(new_n317));
  aoi022aa1n02x5               g222(.a(new_n112), .b(new_n315), .c(new_n316), .d(new_n317), .o1(\s[4] ));
  xorb03aa1n02x5               g223(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g224(.a(new_n119), .b(new_n118), .out0(new_n320));
  aoi012aa1n02x5               g225(.a(new_n120), .b(new_n112), .c(new_n117), .o1(new_n321));
  nanb03aa1n02x5               g226(.a(new_n120), .b(new_n112), .c(new_n117), .out0(new_n322));
  oai112aa1n02x5               g227(.a(new_n322), .b(new_n320), .c(\b[4] ), .d(\a[5] ), .o1(new_n323));
  oai012aa1n02x5               g228(.a(new_n323), .b(new_n321), .c(new_n320), .o1(\s[6] ));
  xnbna2aa1n03x5               g229(.a(new_n127), .b(new_n323), .c(new_n119), .out0(\s[7] ));
  nanb03aa1n02x5               g230(.a(new_n127), .b(new_n323), .c(new_n119), .out0(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n128), .b(new_n326), .c(new_n125), .out0(\s[8] ));
  xnbna2aa1n03x5               g232(.a(new_n174), .b(new_n131), .c(new_n101), .out0(\s[9] ));
endmodule


