// Benchmark "adder" written by ABC on Thu Jul 18 10:38:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n179, new_n180, new_n181,
    new_n182, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n307, new_n310, new_n312, new_n313,
    new_n314;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n15x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  orn002aa1n02x5               g004(.a(\a[9] ), .b(\b[8] ), .o(new_n100));
  inv040aa1d32x5               g005(.a(\a[5] ), .o1(new_n101));
  inv040aa1n16x5               g006(.a(\b[4] ), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  aoi012aa1n06x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .o1(new_n104));
  xnrc02aa1n12x5               g009(.a(\b[7] ), .b(\a[8] ), .out0(new_n105));
  inv000aa1d42x5               g010(.a(\a[6] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[5] ), .o1(new_n107));
  orn002aa1n24x5               g012(.a(\a[7] ), .b(\b[6] ), .o(new_n108));
  nand42aa1n04x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  oai112aa1n06x5               g014(.a(new_n108), .b(new_n109), .c(new_n107), .d(new_n106), .o1(new_n110));
  oao003aa1n03x5               g015(.a(\a[8] ), .b(\b[7] ), .c(new_n108), .carry(new_n111));
  oai013aa1n09x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .d(new_n104), .o1(new_n112));
  nor002aa1n02x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand02aa1d04x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nand22aa1n09x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  tech160nm_fiaoi012aa1n04x5   g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nor022aa1n08x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  tech160nm_finand02aa1n03p5x5 g022(.a(\b[3] ), .b(\a[4] ), .o1(new_n118));
  nor022aa1n16x5               g023(.a(\b[2] ), .b(\a[3] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n120), .b(new_n118), .c(new_n117), .d(new_n119), .out0(new_n121));
  tech160nm_fioai012aa1n03p5x5 g026(.a(new_n118), .b(new_n119), .c(new_n117), .o1(new_n122));
  oai012aa1n12x5               g027(.a(new_n122), .b(new_n121), .c(new_n116), .o1(new_n123));
  nand42aa1n03x5               g028(.a(new_n102), .b(new_n101), .o1(new_n124));
  nand42aa1n03x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  oai112aa1n02x5               g030(.a(new_n124), .b(new_n125), .c(\b[5] ), .d(\a[6] ), .o1(new_n126));
  nor043aa1n06x5               g031(.a(new_n110), .b(new_n126), .c(new_n105), .o1(new_n127));
  nor002aa1d24x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nand02aa1d16x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  norb02aa1d27x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n112), .c(new_n123), .d(new_n127), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n99), .b(new_n131), .c(new_n100), .out0(\s[10] ));
  inv040aa1n02x5               g037(.a(new_n99), .o1(new_n133));
  oai012aa1d24x5               g038(.a(new_n98), .b(new_n128), .c(new_n97), .o1(new_n134));
  inv040aa1n02x5               g039(.a(new_n134), .o1(new_n135));
  oab012aa1n06x5               g040(.a(new_n135), .b(new_n131), .c(new_n133), .out0(new_n136));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  inv040aa1n03x5               g042(.a(new_n137), .o1(new_n138));
  nand42aa1d28x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n136), .b(new_n139), .c(new_n138), .out0(\s[11] ));
  oaoi03aa1n03x5               g045(.a(\a[11] ), .b(\b[10] ), .c(new_n136), .o1(new_n141));
  xorb03aa1n02x5               g046(.a(new_n141), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  aoi012aa1d18x5               g047(.a(new_n112), .b(new_n123), .c(new_n127), .o1(new_n143));
  norb02aa1n15x5               g048(.a(new_n139), .b(new_n137), .out0(new_n144));
  nor042aa1n06x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nanp02aa1n12x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  norb02aa1d21x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  nano32aa1d15x5               g052(.a(new_n133), .b(new_n147), .c(new_n130), .d(new_n144), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  oaoi03aa1n02x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n138), .o1(new_n150));
  nona23aa1n03x5               g055(.a(new_n146), .b(new_n139), .c(new_n137), .d(new_n145), .out0(new_n151));
  oabi12aa1n02x7               g056(.a(new_n150), .b(new_n151), .c(new_n134), .out0(new_n152));
  oabi12aa1n06x5               g057(.a(new_n152), .b(new_n143), .c(new_n149), .out0(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  orn002aa1n24x5               g059(.a(\a[13] ), .b(\b[12] ), .o(new_n155));
  nand42aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  aobi12aa1n02x5               g061(.a(new_n155), .b(new_n153), .c(new_n156), .out0(new_n157));
  xnrb03aa1n03x5               g062(.a(new_n157), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nano23aa1n02x5               g063(.a(new_n137), .b(new_n145), .c(new_n146), .d(new_n139), .out0(new_n159));
  tech160nm_fixnrc02aa1n05x5   g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  nano22aa1d15x5               g065(.a(new_n160), .b(new_n155), .c(new_n156), .out0(new_n161));
  aoai13aa1n03x5               g066(.a(new_n161), .b(new_n150), .c(new_n159), .d(new_n135), .o1(new_n162));
  tech160nm_fioaoi03aa1n02p5x5 g067(.a(\a[14] ), .b(\b[13] ), .c(new_n155), .o1(new_n163));
  inv000aa1n02x5               g068(.a(new_n163), .o1(new_n164));
  nano22aa1n03x7               g069(.a(new_n143), .b(new_n148), .c(new_n161), .out0(new_n165));
  nano22aa1n03x7               g070(.a(new_n165), .b(new_n162), .c(new_n164), .out0(new_n166));
  xnrb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  oaoi03aa1n03x5               g072(.a(\a[15] ), .b(\b[14] ), .c(new_n166), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  tech160nm_fixnrc02aa1n02p5x5 g074(.a(\b[14] ), .b(\a[15] ), .out0(new_n170));
  tech160nm_fixnrc02aa1n02p5x5 g075(.a(\b[15] ), .b(\a[16] ), .out0(new_n171));
  nor042aa1n06x5               g076(.a(new_n171), .b(new_n170), .o1(new_n172));
  aoai13aa1n02x7               g077(.a(new_n172), .b(new_n163), .c(new_n152), .d(new_n161), .o1(new_n173));
  oai022aa1n02x5               g078(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n174));
  aob012aa1n02x5               g079(.a(new_n174), .b(\b[15] ), .c(\a[16] ), .out0(new_n175));
  nand23aa1d12x5               g080(.a(new_n148), .b(new_n161), .c(new_n172), .o1(new_n176));
  oai112aa1n06x5               g081(.a(new_n175), .b(new_n173), .c(new_n143), .d(new_n176), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g083(.a(\a[18] ), .o1(new_n179));
  inv040aa1d32x5               g084(.a(\a[17] ), .o1(new_n180));
  inv030aa1d32x5               g085(.a(\b[16] ), .o1(new_n181));
  oaoi03aa1n03x5               g086(.a(new_n180), .b(new_n181), .c(new_n177), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[17] ), .c(new_n179), .out0(\s[18] ));
  inv040aa1n03x5               g088(.a(new_n143), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n172), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n175), .b(new_n185), .c(new_n162), .d(new_n164), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n176), .o1(new_n187));
  xroi22aa1d06x4               g092(.a(new_n180), .b(\b[16] ), .c(new_n179), .d(\b[17] ), .out0(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n186), .c(new_n184), .d(new_n187), .o1(new_n189));
  oaih22aa1n04x5               g094(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n190));
  oaib12aa1n06x5               g095(.a(new_n190), .b(new_n179), .c(\b[17] ), .out0(new_n191));
  nor002aa1d32x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nand42aa1d28x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  norb02aa1n02x5               g098(.a(new_n193), .b(new_n192), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n189), .c(new_n191), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g101(.a(new_n192), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n181), .b(new_n180), .o1(new_n198));
  oaoi03aa1n12x5               g103(.a(\a[18] ), .b(\b[17] ), .c(new_n198), .o1(new_n199));
  aoai13aa1n03x5               g104(.a(new_n194), .b(new_n199), .c(new_n177), .d(new_n188), .o1(new_n200));
  nor042aa1n12x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand02aa1d28x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n03x4               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  inv000aa1n02x5               g108(.a(new_n203), .o1(new_n204));
  aoi012aa1n03x5               g109(.a(new_n204), .b(new_n200), .c(new_n197), .o1(new_n205));
  nona22aa1n03x5               g110(.a(new_n200), .b(new_n203), .c(new_n192), .out0(new_n206));
  norb02aa1n02x7               g111(.a(new_n206), .b(new_n205), .out0(\s[20] ));
  nona23aa1d18x5               g112(.a(new_n188), .b(new_n193), .c(new_n204), .d(new_n192), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n186), .c(new_n184), .d(new_n187), .o1(new_n210));
  tech160nm_fioaoi03aa1n03p5x5 g115(.a(\a[20] ), .b(\b[19] ), .c(new_n197), .o1(new_n211));
  inv040aa1n03x5               g116(.a(new_n211), .o1(new_n212));
  nona23aa1n12x5               g117(.a(new_n202), .b(new_n193), .c(new_n192), .d(new_n201), .out0(new_n213));
  oai012aa1n18x5               g118(.a(new_n212), .b(new_n213), .c(new_n191), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n210), .c(new_n215), .out0(\s[21] ));
  orn002aa1n24x5               g122(.a(\a[21] ), .b(\b[20] ), .o(new_n218));
  aoai13aa1n03x5               g123(.a(new_n216), .b(new_n214), .c(new_n177), .d(new_n209), .o1(new_n219));
  xnrc02aa1n12x5               g124(.a(\b[21] ), .b(\a[22] ), .out0(new_n220));
  aoi012aa1n03x5               g125(.a(new_n220), .b(new_n219), .c(new_n218), .o1(new_n221));
  aobi12aa1n02x5               g126(.a(new_n216), .b(new_n210), .c(new_n215), .out0(new_n222));
  nano22aa1n02x4               g127(.a(new_n222), .b(new_n218), .c(new_n220), .out0(new_n223));
  nor002aa1n02x5               g128(.a(new_n221), .b(new_n223), .o1(\s[22] ));
  nanp02aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  nano22aa1n12x5               g130(.a(new_n220), .b(new_n218), .c(new_n225), .out0(new_n226));
  norb02aa1n03x5               g131(.a(new_n226), .b(new_n208), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n186), .c(new_n184), .d(new_n187), .o1(new_n228));
  oaoi03aa1n12x5               g133(.a(\a[22] ), .b(\b[21] ), .c(new_n218), .o1(new_n229));
  aoi012aa1n02x5               g134(.a(new_n229), .b(new_n214), .c(new_n226), .o1(new_n230));
  xnrc02aa1n12x5               g135(.a(\b[22] ), .b(\a[23] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  xnbna2aa1n03x5               g137(.a(new_n232), .b(new_n228), .c(new_n230), .out0(\s[23] ));
  orn002aa1n02x5               g138(.a(\a[23] ), .b(\b[22] ), .o(new_n234));
  inv030aa1n02x5               g139(.a(new_n230), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n232), .b(new_n235), .c(new_n177), .d(new_n227), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[23] ), .b(\a[24] ), .out0(new_n237));
  aoi012aa1n03x5               g142(.a(new_n237), .b(new_n236), .c(new_n234), .o1(new_n238));
  tech160nm_fiaoi012aa1n02p5x5 g143(.a(new_n231), .b(new_n228), .c(new_n230), .o1(new_n239));
  nano22aa1n02x4               g144(.a(new_n239), .b(new_n234), .c(new_n237), .out0(new_n240));
  nor002aa1n02x5               g145(.a(new_n238), .b(new_n240), .o1(\s[24] ));
  nano23aa1n03x7               g146(.a(new_n192), .b(new_n201), .c(new_n202), .d(new_n193), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n226), .b(new_n211), .c(new_n242), .d(new_n199), .o1(new_n243));
  inv000aa1n02x5               g148(.a(new_n229), .o1(new_n244));
  nor042aa1n06x5               g149(.a(new_n237), .b(new_n231), .o1(new_n245));
  inv030aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  oao003aa1n02x5               g151(.a(\a[24] ), .b(\b[23] ), .c(new_n234), .carry(new_n247));
  aoai13aa1n12x5               g152(.a(new_n247), .b(new_n246), .c(new_n243), .d(new_n244), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  nano22aa1n03x7               g154(.a(new_n208), .b(new_n226), .c(new_n245), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n186), .c(new_n184), .d(new_n187), .o1(new_n251));
  xnrc02aa1n12x5               g156(.a(\b[24] ), .b(\a[25] ), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  xnbna2aa1n03x5               g158(.a(new_n253), .b(new_n251), .c(new_n249), .out0(\s[25] ));
  nor042aa1n03x5               g159(.a(\b[24] ), .b(\a[25] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n03x5               g161(.a(new_n253), .b(new_n248), .c(new_n177), .d(new_n250), .o1(new_n257));
  tech160nm_fixnrc02aa1n05x5   g162(.a(\b[25] ), .b(\a[26] ), .out0(new_n258));
  aoi012aa1n03x5               g163(.a(new_n258), .b(new_n257), .c(new_n256), .o1(new_n259));
  aoi012aa1n02x5               g164(.a(new_n252), .b(new_n251), .c(new_n249), .o1(new_n260));
  nano22aa1n03x5               g165(.a(new_n260), .b(new_n256), .c(new_n258), .out0(new_n261));
  nor002aa1n02x5               g166(.a(new_n259), .b(new_n261), .o1(\s[26] ));
  nor042aa1n06x5               g167(.a(new_n258), .b(new_n252), .o1(new_n263));
  nano32aa1d12x5               g168(.a(new_n208), .b(new_n263), .c(new_n226), .d(new_n245), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n186), .c(new_n184), .d(new_n187), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[26] ), .b(\b[25] ), .c(new_n256), .carry(new_n266));
  aobi12aa1n12x5               g171(.a(new_n266), .b(new_n248), .c(new_n263), .out0(new_n267));
  xorc02aa1n12x5               g172(.a(\a[27] ), .b(\b[26] ), .out0(new_n268));
  xnbna2aa1n03x5               g173(.a(new_n268), .b(new_n265), .c(new_n267), .out0(\s[27] ));
  norp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  inv040aa1n03x5               g175(.a(new_n270), .o1(new_n271));
  aoai13aa1n03x5               g176(.a(new_n245), .b(new_n229), .c(new_n214), .d(new_n226), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n263), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n266), .b(new_n273), .c(new_n272), .d(new_n247), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n268), .b(new_n274), .c(new_n177), .d(new_n264), .o1(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[27] ), .b(\a[28] ), .out0(new_n276));
  aoi012aa1n02x5               g181(.a(new_n276), .b(new_n275), .c(new_n271), .o1(new_n277));
  aobi12aa1n03x5               g182(.a(new_n268), .b(new_n265), .c(new_n267), .out0(new_n278));
  nano22aa1n03x5               g183(.a(new_n278), .b(new_n271), .c(new_n276), .out0(new_n279));
  norp02aa1n03x5               g184(.a(new_n277), .b(new_n279), .o1(\s[28] ));
  xnrc02aa1n02x5               g185(.a(\b[28] ), .b(\a[29] ), .out0(new_n281));
  norb02aa1n02x5               g186(.a(new_n268), .b(new_n276), .out0(new_n282));
  aoai13aa1n02x7               g187(.a(new_n282), .b(new_n274), .c(new_n177), .d(new_n264), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .c(new_n271), .carry(new_n284));
  aoi012aa1n03x5               g189(.a(new_n281), .b(new_n283), .c(new_n284), .o1(new_n285));
  aobi12aa1n03x5               g190(.a(new_n282), .b(new_n265), .c(new_n267), .out0(new_n286));
  nano22aa1n03x5               g191(.a(new_n286), .b(new_n281), .c(new_n284), .out0(new_n287));
  norp02aa1n03x5               g192(.a(new_n285), .b(new_n287), .o1(\s[29] ));
  xorb03aa1n02x5               g193(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  norb03aa1n02x5               g195(.a(new_n268), .b(new_n281), .c(new_n276), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n274), .c(new_n177), .d(new_n264), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .carry(new_n293));
  aoi012aa1n03x5               g198(.a(new_n290), .b(new_n292), .c(new_n293), .o1(new_n294));
  aobi12aa1n06x5               g199(.a(new_n291), .b(new_n265), .c(new_n267), .out0(new_n295));
  nano22aa1n03x7               g200(.a(new_n295), .b(new_n290), .c(new_n293), .out0(new_n296));
  norp02aa1n03x5               g201(.a(new_n294), .b(new_n296), .o1(\s[30] ));
  xnrc02aa1n02x5               g202(.a(\b[30] ), .b(\a[31] ), .out0(new_n298));
  norb02aa1n03x4               g203(.a(new_n291), .b(new_n290), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n274), .c(new_n177), .d(new_n264), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n301));
  aoi012aa1n03x5               g206(.a(new_n298), .b(new_n300), .c(new_n301), .o1(new_n302));
  aobi12aa1n06x5               g207(.a(new_n299), .b(new_n265), .c(new_n267), .out0(new_n303));
  nano22aa1n03x7               g208(.a(new_n303), .b(new_n298), .c(new_n301), .out0(new_n304));
  norp02aa1n03x5               g209(.a(new_n302), .b(new_n304), .o1(\s[31] ));
  xnrb03aa1n02x5               g210(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g211(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g213(.a(new_n123), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aob012aa1n02x5               g214(.a(new_n124), .b(new_n123), .c(new_n125), .out0(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oabi12aa1n02x5               g216(.a(new_n110), .b(new_n310), .c(new_n103), .out0(new_n312));
  xorc02aa1n02x5               g217(.a(\a[6] ), .b(\b[5] ), .out0(new_n313));
  aoi122aa1n02x5               g218(.a(new_n103), .b(new_n109), .c(new_n108), .d(new_n310), .e(new_n313), .o1(new_n314));
  norb02aa1n02x5               g219(.a(new_n312), .b(new_n314), .out0(\s[7] ));
  xobna2aa1n03x5               g220(.a(new_n105), .b(new_n312), .c(new_n108), .out0(\s[8] ));
  xnbna2aa1n03x5               g221(.a(new_n143), .b(new_n129), .c(new_n100), .out0(\s[9] ));
endmodule


