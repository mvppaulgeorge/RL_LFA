// Benchmark "adder" written by ABC on Wed Jul 17 22:59:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n319, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n341, new_n342, new_n344, new_n346,
    new_n348, new_n350, new_n351, new_n352, new_n354, new_n356, new_n357,
    new_n358;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1n03x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norp02aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  aoi012aa1n02x7               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  nand42aa1n16x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand42aa1d28x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano22aa1n03x7               g010(.a(new_n102), .b(new_n104), .c(new_n105), .out0(new_n106));
  nor042aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nand03aa1n02x5               g012(.a(new_n104), .b(\a[1] ), .c(\b[0] ), .o1(new_n108));
  norb02aa1n06x5               g013(.a(new_n101), .b(new_n100), .out0(new_n109));
  oai112aa1n06x5               g014(.a(new_n106), .b(new_n109), .c(new_n108), .d(new_n107), .o1(new_n110));
  nor022aa1n08x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nano23aa1n06x5               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  xorc02aa1n02x5               g020(.a(\a[6] ), .b(\b[5] ), .out0(new_n116));
  xorc02aa1n02x5               g021(.a(\a[5] ), .b(\b[4] ), .out0(new_n117));
  nanp03aa1n02x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  nor042aa1n06x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  inv040aa1n02x5               g024(.a(new_n119), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[6] ), .b(\b[5] ), .c(new_n120), .o1(new_n121));
  oai012aa1n02x5               g026(.a(new_n112), .b(new_n113), .c(new_n111), .o1(new_n122));
  aobi12aa1n06x5               g027(.a(new_n122), .b(new_n115), .c(new_n121), .out0(new_n123));
  aoai13aa1n06x5               g028(.a(new_n123), .b(new_n118), .c(new_n110), .d(new_n103), .o1(new_n124));
  aob012aa1n06x5               g029(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n97), .b(new_n125), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g031(.a(new_n97), .o1(new_n127));
  nona22aa1n06x5               g032(.a(new_n125), .b(new_n98), .c(new_n127), .out0(new_n128));
  and002aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o(new_n129));
  nanp02aa1n04x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor022aa1n08x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb03aa1n02x5               g036(.a(new_n130), .b(new_n129), .c(new_n131), .out0(new_n132));
  nanb02aa1n02x5               g037(.a(new_n131), .b(new_n130), .out0(new_n133));
  nanb02aa1n02x5               g038(.a(new_n129), .b(new_n128), .out0(new_n134));
  aoi022aa1n02x5               g039(.a(new_n134), .b(new_n133), .c(new_n128), .d(new_n132), .o1(\s[11] ));
  nor002aa1n20x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n136), .o1(new_n137));
  nanp02aa1n06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  aoi122aa1n02x5               g043(.a(new_n131), .b(new_n137), .c(new_n138), .d(new_n128), .e(new_n132), .o1(new_n139));
  tech160nm_fiao0012aa1n02p5x5 g044(.a(new_n131), .b(new_n128), .c(new_n132), .o(new_n140));
  aoi013aa1n02x4               g045(.a(new_n139), .b(new_n140), .c(new_n137), .d(new_n138), .o1(\s[12] ));
  nand02aa1d06x5               g046(.a(new_n110), .b(new_n103), .o1(new_n142));
  nona23aa1n03x5               g047(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n143));
  xnrc02aa1n02x5               g048(.a(\b[5] ), .b(\a[6] ), .out0(new_n144));
  norb03aa1n03x5               g049(.a(new_n117), .b(new_n143), .c(new_n144), .out0(new_n145));
  oaib12aa1n03x5               g050(.a(new_n122), .b(new_n143), .c(new_n121), .out0(new_n146));
  nano23aa1n06x5               g051(.a(new_n136), .b(new_n131), .c(new_n138), .d(new_n130), .out0(new_n147));
  xorc02aa1n12x5               g052(.a(\a[9] ), .b(\b[8] ), .out0(new_n148));
  nand23aa1d12x5               g053(.a(new_n147), .b(new_n97), .c(new_n148), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n146), .c(new_n142), .d(new_n145), .o1(new_n151));
  nona23aa1n02x4               g056(.a(new_n130), .b(new_n138), .c(new_n136), .d(new_n131), .out0(new_n152));
  oai022aa1n02x5               g057(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n153));
  aob012aa1n02x5               g058(.a(new_n153), .b(\b[9] ), .c(\a[10] ), .out0(new_n154));
  aob012aa1d15x5               g059(.a(new_n137), .b(new_n131), .c(new_n138), .out0(new_n155));
  oabi12aa1n06x5               g060(.a(new_n155), .b(new_n152), .c(new_n154), .out0(new_n156));
  xnrc02aa1n12x5               g061(.a(\b[12] ), .b(\a[13] ), .out0(new_n157));
  aoib12aa1n06x5               g062(.a(new_n157), .b(new_n151), .c(new_n156), .out0(new_n158));
  oaoi03aa1n02x5               g063(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n157), .o1(new_n160));
  aoi112aa1n02x5               g065(.a(new_n160), .b(new_n155), .c(new_n147), .d(new_n159), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n158), .b(new_n151), .c(new_n161), .o1(\s[13] ));
  nor042aa1n03x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  inv000aa1d42x5               g068(.a(\a[14] ), .o1(new_n164));
  inv000aa1d42x5               g069(.a(\b[13] ), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(new_n165), .b(new_n164), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  aoi112aa1n02x5               g072(.a(new_n158), .b(new_n163), .c(new_n166), .d(new_n167), .o1(new_n168));
  oai112aa1n02x5               g073(.a(new_n166), .b(new_n167), .c(new_n158), .d(new_n163), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(\s[14] ));
  nano22aa1n09x5               g075(.a(new_n157), .b(new_n166), .c(new_n167), .out0(new_n171));
  nanp03aa1n03x5               g076(.a(new_n124), .b(new_n150), .c(new_n171), .o1(new_n172));
  oaoi03aa1n06x5               g077(.a(new_n164), .b(new_n165), .c(new_n163), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  aoi012aa1n02x5               g079(.a(new_n174), .b(new_n156), .c(new_n171), .o1(new_n175));
  nor042aa1n04x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nand42aa1n03x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  aobi12aa1n06x5               g083(.a(new_n178), .b(new_n172), .c(new_n175), .out0(new_n179));
  aoi112aa1n02x5               g084(.a(new_n178), .b(new_n174), .c(new_n156), .d(new_n171), .o1(new_n180));
  aoi012aa1n02x5               g085(.a(new_n179), .b(new_n172), .c(new_n180), .o1(\s[15] ));
  nand42aa1n06x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nor042aa1n04x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  norp03aa1n02x5               g089(.a(new_n179), .b(new_n184), .c(new_n176), .o1(new_n185));
  oab012aa1n02x4               g090(.a(new_n183), .b(new_n179), .c(new_n176), .out0(new_n186));
  aoi012aa1n02x5               g091(.a(new_n185), .b(new_n186), .c(new_n182), .o1(\s[16] ));
  nano23aa1d15x5               g092(.a(new_n176), .b(new_n183), .c(new_n182), .d(new_n177), .out0(new_n188));
  nano22aa1d15x5               g093(.a(new_n149), .b(new_n171), .c(new_n188), .out0(new_n189));
  aoai13aa1n09x5               g094(.a(new_n189), .b(new_n146), .c(new_n142), .d(new_n145), .o1(new_n190));
  aoai13aa1n06x5               g095(.a(new_n188), .b(new_n174), .c(new_n156), .d(new_n171), .o1(new_n191));
  aoi012aa1n12x5               g096(.a(new_n183), .b(new_n176), .c(new_n182), .o1(new_n192));
  nanp03aa1d12x5               g097(.a(new_n190), .b(new_n191), .c(new_n192), .o1(new_n193));
  tech160nm_fixnrc02aa1n04x5   g098(.a(\b[16] ), .b(\a[17] ), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n171), .b(new_n155), .c(new_n147), .d(new_n159), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n188), .o1(new_n196));
  tech160nm_fiaoi012aa1n04x5   g101(.a(new_n196), .b(new_n195), .c(new_n173), .o1(new_n197));
  nano22aa1n02x4               g102(.a(new_n197), .b(new_n192), .c(new_n194), .out0(new_n198));
  aboi22aa1n03x5               g103(.a(new_n194), .b(new_n193), .c(new_n198), .d(new_n190), .out0(\s[17] ));
  inv000aa1d42x5               g104(.a(\a[18] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[17] ), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(new_n201), .b(new_n200), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norp02aa1n02x5               g108(.a(\b[16] ), .b(\a[17] ), .o1(new_n204));
  aoi013aa1n02x4               g109(.a(new_n194), .b(new_n190), .c(new_n191), .d(new_n192), .o1(new_n205));
  aoi112aa1n02x5               g110(.a(new_n205), .b(new_n204), .c(new_n202), .d(new_n203), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n192), .o1(new_n207));
  aoi112aa1n03x5               g112(.a(new_n197), .b(new_n207), .c(new_n124), .d(new_n189), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(\a[17] ), .b(\b[16] ), .c(new_n208), .o1(new_n209));
  aoi013aa1n02x4               g114(.a(new_n206), .b(new_n209), .c(new_n202), .d(new_n203), .o1(\s[18] ));
  nano22aa1n02x4               g115(.a(new_n194), .b(new_n202), .c(new_n203), .out0(new_n211));
  aob012aa1n02x5               g116(.a(new_n202), .b(new_n204), .c(new_n203), .out0(new_n212));
  nor042aa1n06x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n212), .c(new_n193), .d(new_n211), .o1(new_n216));
  aoi112aa1n02x5               g121(.a(new_n215), .b(new_n212), .c(new_n193), .d(new_n211), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n216), .b(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g124(.a(new_n213), .o1(new_n220));
  nor002aa1n04x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand22aa1n09x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n222), .o1(new_n224));
  oai022aa1n02x5               g129(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n225));
  nona22aa1n03x5               g130(.a(new_n216), .b(new_n224), .c(new_n225), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n220), .d(new_n216), .o1(\s[20] ));
  nona23aa1n09x5               g132(.a(new_n222), .b(new_n214), .c(new_n213), .d(new_n221), .out0(new_n228));
  nano23aa1n03x7               g133(.a(new_n228), .b(new_n194), .c(new_n202), .d(new_n203), .out0(new_n229));
  oaoi03aa1n02x5               g134(.a(new_n200), .b(new_n201), .c(new_n204), .o1(new_n230));
  aoi012aa1d18x5               g135(.a(new_n221), .b(new_n213), .c(new_n222), .o1(new_n231));
  tech160nm_fioai012aa1n05x5   g136(.a(new_n231), .b(new_n228), .c(new_n230), .o1(new_n232));
  nor042aa1n03x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  nanp02aa1n02x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n232), .c(new_n193), .d(new_n229), .o1(new_n236));
  nano23aa1n06x5               g141(.a(new_n213), .b(new_n221), .c(new_n222), .d(new_n214), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n231), .o1(new_n238));
  aoi112aa1n02x5               g143(.a(new_n238), .b(new_n235), .c(new_n237), .d(new_n212), .o1(new_n239));
  aobi12aa1n02x5               g144(.a(new_n239), .b(new_n193), .c(new_n229), .out0(new_n240));
  norb02aa1n02x5               g145(.a(new_n236), .b(new_n240), .out0(\s[21] ));
  inv000aa1n06x5               g146(.a(new_n233), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  and002aa1n02x5               g149(.a(\b[21] ), .b(\a[22] ), .o(new_n245));
  oai022aa1n02x5               g150(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n246));
  nona22aa1n03x5               g151(.a(new_n236), .b(new_n245), .c(new_n246), .out0(new_n247));
  aoai13aa1n03x5               g152(.a(new_n247), .b(new_n244), .c(new_n242), .d(new_n236), .o1(\s[22] ));
  nano22aa1d18x5               g153(.a(new_n243), .b(new_n242), .c(new_n234), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  nano22aa1n02x4               g155(.a(new_n250), .b(new_n211), .c(new_n237), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n249), .b(new_n238), .c(new_n237), .d(new_n212), .o1(new_n252));
  oao003aa1n02x5               g157(.a(\a[22] ), .b(\b[21] ), .c(new_n242), .carry(new_n253));
  nanp02aa1n02x5               g158(.a(new_n252), .b(new_n253), .o1(new_n254));
  tech160nm_fixorc02aa1n03p5x5 g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n193), .d(new_n251), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n253), .o1(new_n257));
  nona22aa1n02x4               g162(.a(new_n252), .b(new_n257), .c(new_n255), .out0(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(new_n193), .c(new_n251), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n256), .b(new_n259), .out0(\s[23] ));
  nor042aa1n03x5               g165(.a(\b[22] ), .b(\a[23] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .out0(new_n263));
  and002aa1n02x5               g168(.a(\b[23] ), .b(\a[24] ), .o(new_n264));
  oai022aa1n02x5               g169(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n265));
  nona22aa1n03x5               g170(.a(new_n256), .b(new_n264), .c(new_n265), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n266), .b(new_n263), .c(new_n262), .d(new_n256), .o1(\s[24] ));
  and002aa1n18x5               g172(.a(new_n263), .b(new_n255), .o(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  nano32aa1n02x4               g174(.a(new_n269), .b(new_n249), .c(new_n211), .d(new_n237), .out0(new_n270));
  oao003aa1n03x5               g175(.a(\a[24] ), .b(\b[23] ), .c(new_n262), .carry(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n269), .c(new_n252), .d(new_n253), .o1(new_n272));
  xorc02aa1n12x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n272), .c(new_n193), .d(new_n270), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n268), .b(new_n257), .c(new_n232), .d(new_n249), .o1(new_n275));
  nanb03aa1n02x5               g180(.a(new_n273), .b(new_n275), .c(new_n271), .out0(new_n276));
  aoi012aa1n02x5               g181(.a(new_n276), .b(new_n193), .c(new_n270), .o1(new_n277));
  norb02aa1n02x5               g182(.a(new_n274), .b(new_n277), .out0(\s[25] ));
  nor042aa1n03x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  xorc02aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .out0(new_n281));
  and002aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .o(new_n282));
  oai022aa1n02x5               g187(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n283));
  nona22aa1n03x5               g188(.a(new_n274), .b(new_n282), .c(new_n283), .out0(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n281), .c(new_n280), .d(new_n274), .o1(\s[26] ));
  and002aa1n02x5               g190(.a(new_n281), .b(new_n273), .o(new_n286));
  inv000aa1n02x5               g191(.a(new_n286), .o1(new_n287));
  nano32aa1n03x7               g192(.a(new_n287), .b(new_n229), .c(new_n249), .d(new_n268), .out0(new_n288));
  nanp02aa1n02x5               g193(.a(new_n193), .b(new_n288), .o1(new_n289));
  inv000aa1n02x5               g194(.a(new_n288), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n280), .carry(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoi012aa1n02x5               g197(.a(new_n292), .b(new_n272), .c(new_n286), .o1(new_n293));
  oai012aa1n04x7               g198(.a(new_n293), .b(new_n208), .c(new_n290), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoi112aa1n02x5               g200(.a(new_n295), .b(new_n292), .c(new_n272), .d(new_n286), .o1(new_n296));
  aoi022aa1n02x5               g201(.a(new_n294), .b(new_n295), .c(new_n289), .d(new_n296), .o1(\s[27] ));
  nor042aa1n03x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[27] ), .b(\a[28] ), .out0(new_n299));
  aoai13aa1n02x5               g204(.a(new_n299), .b(new_n298), .c(new_n294), .d(new_n295), .o1(new_n300));
  aoai13aa1n04x5               g205(.a(new_n291), .b(new_n287), .c(new_n275), .d(new_n271), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n295), .b(new_n301), .c(new_n193), .d(new_n288), .o1(new_n302));
  and002aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .o(new_n303));
  oai022aa1n02x5               g208(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n304));
  nona22aa1n02x4               g209(.a(new_n302), .b(new_n303), .c(new_n304), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n300), .b(new_n305), .o1(\s[28] ));
  norb02aa1n02x5               g211(.a(new_n295), .b(new_n299), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n301), .c(new_n193), .d(new_n288), .o1(new_n308));
  inv000aa1d42x5               g213(.a(\a[28] ), .o1(new_n309));
  inv000aa1d42x5               g214(.a(\b[27] ), .o1(new_n310));
  norp02aa1n02x5               g215(.a(\b[28] ), .b(\a[29] ), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n311), .o1(new_n312));
  oaib12aa1n02x5               g217(.a(new_n312), .b(new_n303), .c(new_n298), .out0(new_n313));
  aoi122aa1n02x5               g218(.a(new_n313), .b(\b[28] ), .c(\a[29] ), .d(new_n310), .e(new_n309), .o1(new_n314));
  nanp02aa1n03x5               g219(.a(new_n308), .b(new_n314), .o1(new_n315));
  tech160nm_fioaoi03aa1n03p5x5 g220(.a(new_n309), .b(new_n310), .c(new_n298), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n315), .b(new_n317), .c(new_n308), .d(new_n316), .o1(\s[29] ));
  nanp02aa1n02x5               g223(.a(\b[0] ), .b(\a[1] ), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g225(.a(new_n299), .b(new_n295), .c(new_n317), .out0(new_n321));
  aoai13aa1n06x5               g226(.a(new_n321), .b(new_n301), .c(new_n193), .d(new_n288), .o1(new_n322));
  oaoi03aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .o1(new_n323));
  inv000aa1d42x5               g228(.a(new_n323), .o1(new_n324));
  norp02aa1n02x5               g229(.a(\b[29] ), .b(\a[30] ), .o1(new_n325));
  nanp02aa1n02x5               g230(.a(\b[29] ), .b(\a[30] ), .o1(new_n326));
  norb02aa1n02x5               g231(.a(new_n326), .b(new_n325), .out0(new_n327));
  aoi012aa1n02x5               g232(.a(new_n316), .b(\a[29] ), .c(\b[28] ), .o1(new_n328));
  nano23aa1n02x4               g233(.a(new_n328), .b(new_n325), .c(new_n326), .d(new_n312), .out0(new_n329));
  nanp02aa1n06x5               g234(.a(new_n322), .b(new_n329), .o1(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n327), .c(new_n322), .d(new_n324), .o1(\s[30] ));
  and003aa1n02x5               g236(.a(new_n307), .b(new_n327), .c(new_n317), .o(new_n332));
  aoai13aa1n06x5               g237(.a(new_n332), .b(new_n301), .c(new_n193), .d(new_n288), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  oai012aa1n02x5               g239(.a(new_n334), .b(\b[29] ), .c(\a[30] ), .o1(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n323), .c(new_n327), .o1(new_n336));
  nanp02aa1n03x5               g241(.a(new_n333), .b(new_n336), .o1(new_n337));
  aoi012aa1n02x5               g242(.a(new_n325), .b(new_n323), .c(new_n327), .o1(new_n338));
  aoai13aa1n03x5               g243(.a(new_n337), .b(new_n334), .c(new_n333), .d(new_n338), .o1(\s[31] ));
  norb03aa1n02x5               g244(.a(new_n104), .b(new_n319), .c(new_n107), .out0(new_n340));
  norb02aa1n02x5               g245(.a(new_n105), .b(new_n102), .out0(new_n341));
  oaoi13aa1n02x5               g246(.a(new_n341), .b(new_n104), .c(new_n319), .d(new_n107), .o1(new_n342));
  aoib12aa1n02x5               g247(.a(new_n342), .b(new_n106), .c(new_n340), .out0(\s[3] ));
  aoai13aa1n02x5               g248(.a(new_n341), .b(new_n340), .c(\b[1] ), .d(\a[2] ), .o1(new_n344));
  xobna2aa1n03x5               g249(.a(new_n109), .b(new_n344), .c(new_n105), .out0(\s[4] ));
  aoi112aa1n02x5               g250(.a(new_n117), .b(new_n100), .c(new_n101), .d(new_n102), .o1(new_n346));
  aoi022aa1n02x5               g251(.a(new_n142), .b(new_n117), .c(new_n110), .d(new_n346), .o1(\s[5] ));
  nanp02aa1n02x5               g252(.a(new_n142), .b(new_n117), .o1(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n116), .b(new_n348), .c(new_n120), .out0(\s[6] ));
  nanb02aa1n02x5               g254(.a(new_n113), .b(new_n114), .out0(new_n350));
  nanp02aa1n02x5               g255(.a(\b[5] ), .b(\a[6] ), .o1(new_n351));
  nona22aa1n02x4               g256(.a(new_n348), .b(new_n119), .c(new_n144), .out0(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n350), .b(new_n352), .c(new_n351), .out0(\s[7] ));
  aoi013aa1n02x4               g258(.a(new_n113), .b(new_n352), .c(new_n351), .d(new_n114), .o1(new_n354));
  xnrb03aa1n02x5               g259(.a(new_n354), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  nanp02aa1n02x5               g260(.a(new_n148), .b(new_n122), .o1(new_n356));
  aoi012aa1n02x5               g261(.a(new_n356), .b(new_n115), .c(new_n121), .o1(new_n357));
  aoai13aa1n02x5               g262(.a(new_n357), .b(new_n118), .c(new_n110), .d(new_n103), .o1(new_n358));
  oaib12aa1n02x5               g263(.a(new_n358), .b(new_n148), .c(new_n124), .out0(\s[9] ));
endmodule


