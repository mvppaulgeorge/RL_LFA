// Benchmark "adder" written by ABC on Thu Jul 18 01:53:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n342, new_n345, new_n346, new_n348,
    new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d48x5               g002(.a(\b[8] ), .o1(new_n98));
  nand42aa1n16x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1d16x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai012aa1d24x5               g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  tech160nm_fixorc02aa1n03p5x5 g007(.a(\a[4] ), .b(\b[3] ), .out0(new_n103));
  nor042aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  norb02aa1n09x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nanb03aa1n06x5               g011(.a(new_n102), .b(new_n103), .c(new_n106), .out0(new_n107));
  inv040aa1d32x5               g012(.a(\a[3] ), .o1(new_n108));
  inv040aa1d28x5               g013(.a(\b[2] ), .o1(new_n109));
  nand42aa1n20x5               g014(.a(new_n109), .b(new_n108), .o1(new_n110));
  oaoi03aa1n09x5               g015(.a(\a[4] ), .b(\b[3] ), .c(new_n110), .o1(new_n111));
  inv040aa1n02x5               g016(.a(new_n111), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1d28x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n24x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n09x5               g021(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n117));
  xorc02aa1n02x5               g022(.a(\a[6] ), .b(\b[5] ), .out0(new_n118));
  xorc02aa1n02x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nand03aa1n02x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  inv040aa1d32x5               g025(.a(\a[6] ), .o1(new_n121));
  inv040aa1d32x5               g026(.a(\b[5] ), .o1(new_n122));
  norp02aa1n12x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  oao003aa1n03x5               g028(.a(new_n121), .b(new_n122), .c(new_n123), .carry(new_n124));
  ao0012aa1n03x7               g029(.a(new_n113), .b(new_n115), .c(new_n114), .o(new_n125));
  aoi012aa1n06x5               g030(.a(new_n125), .b(new_n117), .c(new_n124), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n120), .c(new_n107), .d(new_n112), .o1(new_n127));
  oaoi03aa1n02x5               g032(.a(new_n97), .b(new_n98), .c(new_n127), .o1(new_n128));
  xnrb03aa1n03x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1d32x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand22aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nor042aa1n04x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  nand02aa1d04x5               g037(.a(\b[8] ), .b(\a[9] ), .o1(new_n133));
  nano23aa1n09x5               g038(.a(new_n130), .b(new_n132), .c(new_n133), .d(new_n131), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n135));
  inv000aa1n02x5               g040(.a(new_n135), .o1(new_n136));
  nor002aa1n16x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand02aa1d28x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  aoai13aa1n03x5               g044(.a(new_n139), .b(new_n136), .c(new_n127), .d(new_n134), .o1(new_n140));
  aoi112aa1n02x5               g045(.a(new_n139), .b(new_n136), .c(new_n127), .d(new_n134), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(\s[11] ));
  tech160nm_fioai012aa1n03p5x5 g047(.a(new_n140), .b(\b[10] ), .c(\a[11] ), .o1(new_n143));
  xorb03aa1n02x5               g048(.a(new_n143), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv040aa1d32x5               g049(.a(\a[4] ), .o1(new_n145));
  inv040aa1n20x5               g050(.a(\b[3] ), .o1(new_n146));
  nanp02aa1n04x5               g051(.a(new_n146), .b(new_n145), .o1(new_n147));
  nanp02aa1n04x5               g052(.a(\b[3] ), .b(\a[4] ), .o1(new_n148));
  nand42aa1n08x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  nanp02aa1n04x5               g054(.a(new_n110), .b(new_n105), .o1(new_n150));
  nor043aa1n02x5               g055(.a(new_n102), .b(new_n149), .c(new_n150), .o1(new_n151));
  nona23aa1n09x5               g056(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n152));
  xnrc02aa1n03x5               g057(.a(\b[5] ), .b(\a[6] ), .out0(new_n153));
  xnrc02aa1n12x5               g058(.a(\b[4] ), .b(\a[5] ), .out0(new_n154));
  nor043aa1n03x5               g059(.a(new_n152), .b(new_n153), .c(new_n154), .o1(new_n155));
  tech160nm_fioai012aa1n03p5x5 g060(.a(new_n155), .b(new_n151), .c(new_n111), .o1(new_n156));
  nor022aa1n16x5               g061(.a(\b[11] ), .b(\a[12] ), .o1(new_n157));
  nand22aa1n12x5               g062(.a(\b[11] ), .b(\a[12] ), .o1(new_n158));
  nano23aa1n03x7               g063(.a(new_n137), .b(new_n157), .c(new_n158), .d(new_n138), .out0(new_n159));
  nanp02aa1n03x5               g064(.a(new_n159), .b(new_n134), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n157), .b(new_n137), .c(new_n158), .o1(new_n161));
  aobi12aa1n06x5               g066(.a(new_n161), .b(new_n159), .c(new_n136), .out0(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n160), .c(new_n156), .d(new_n126), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d28x5               g069(.a(\a[13] ), .o1(new_n165));
  inv040aa1d32x5               g070(.a(\b[12] ), .o1(new_n166));
  oaoi03aa1n03x5               g071(.a(new_n165), .b(new_n166), .c(new_n163), .o1(new_n167));
  xnrb03aa1n03x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  oai013aa1n03x5               g073(.a(new_n112), .b(new_n149), .c(new_n102), .d(new_n150), .o1(new_n169));
  oaoi03aa1n02x5               g074(.a(new_n121), .b(new_n122), .c(new_n123), .o1(new_n170));
  oabi12aa1n02x7               g075(.a(new_n125), .b(new_n152), .c(new_n170), .out0(new_n171));
  inv000aa1n02x5               g076(.a(new_n160), .o1(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n171), .c(new_n169), .d(new_n155), .o1(new_n173));
  nor022aa1n16x5               g078(.a(\b[12] ), .b(\a[13] ), .o1(new_n174));
  nand02aa1n03x5               g079(.a(\b[12] ), .b(\a[13] ), .o1(new_n175));
  nor002aa1d32x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  nand42aa1d28x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nona23aa1n02x4               g082(.a(new_n177), .b(new_n175), .c(new_n174), .d(new_n176), .out0(new_n178));
  aoai13aa1n12x5               g083(.a(new_n177), .b(new_n176), .c(new_n165), .d(new_n166), .o1(new_n179));
  aoai13aa1n03x5               g084(.a(new_n179), .b(new_n178), .c(new_n173), .d(new_n162), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nand22aa1n12x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  nanb02aa1d24x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  inv000aa1d42x5               g089(.a(new_n184), .o1(new_n185));
  nor002aa1d32x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nand02aa1d08x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nanb02aa1n12x5               g092(.a(new_n186), .b(new_n187), .out0(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  aoi112aa1n03x4               g094(.a(new_n189), .b(new_n182), .c(new_n180), .d(new_n185), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n182), .o1(new_n191));
  nano23aa1n03x7               g096(.a(new_n174), .b(new_n176), .c(new_n177), .d(new_n175), .out0(new_n192));
  inv000aa1d42x5               g097(.a(new_n179), .o1(new_n193));
  aoai13aa1n03x5               g098(.a(new_n185), .b(new_n193), .c(new_n163), .d(new_n192), .o1(new_n194));
  tech160nm_fiaoi012aa1n02p5x5 g099(.a(new_n188), .b(new_n194), .c(new_n191), .o1(new_n195));
  norp02aa1n03x5               g100(.a(new_n195), .b(new_n190), .o1(\s[16] ));
  nona23aa1n03x5               g101(.a(new_n158), .b(new_n138), .c(new_n137), .d(new_n157), .out0(new_n197));
  nona23aa1n09x5               g102(.a(new_n187), .b(new_n183), .c(new_n182), .d(new_n186), .out0(new_n198));
  nona23aa1n03x5               g103(.a(new_n192), .b(new_n134), .c(new_n198), .d(new_n197), .out0(new_n199));
  tech160nm_fioai012aa1n03p5x5 g104(.a(new_n161), .b(new_n197), .c(new_n135), .o1(new_n200));
  nor042aa1n02x5               g105(.a(new_n198), .b(new_n178), .o1(new_n201));
  tech160nm_fiaoi012aa1n03p5x5 g106(.a(new_n186), .b(new_n182), .c(new_n187), .o1(new_n202));
  oai012aa1n06x5               g107(.a(new_n202), .b(new_n198), .c(new_n179), .o1(new_n203));
  aoi012aa1n12x5               g108(.a(new_n203), .b(new_n200), .c(new_n201), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n199), .c(new_n156), .d(new_n126), .o1(new_n205));
  xorb03aa1n03x5               g110(.a(new_n205), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g111(.a(\a[18] ), .o1(new_n207));
  inv040aa1n09x5               g112(.a(\a[17] ), .o1(new_n208));
  inv000aa1d42x5               g113(.a(\b[16] ), .o1(new_n209));
  oaoi03aa1n03x5               g114(.a(new_n208), .b(new_n209), .c(new_n205), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[17] ), .c(new_n207), .out0(\s[18] ));
  nona22aa1n03x5               g116(.a(new_n192), .b(new_n188), .c(new_n184), .out0(new_n212));
  nor042aa1n03x5               g117(.a(new_n212), .b(new_n160), .o1(new_n213));
  aoai13aa1n06x5               g118(.a(new_n213), .b(new_n171), .c(new_n169), .d(new_n155), .o1(new_n214));
  xroi22aa1d06x4               g119(.a(new_n208), .b(\b[16] ), .c(new_n207), .d(\b[17] ), .out0(new_n215));
  inv000aa1n02x5               g120(.a(new_n215), .o1(new_n216));
  inv040aa1d28x5               g121(.a(\b[17] ), .o1(new_n217));
  oai022aa1d24x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  oaib12aa1n18x5               g123(.a(new_n218), .b(new_n217), .c(\a[18] ), .out0(new_n219));
  aoai13aa1n02x7               g124(.a(new_n219), .b(new_n216), .c(new_n214), .d(new_n204), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1d18x5               g127(.a(\b[18] ), .b(\a[19] ), .o1(new_n223));
  xorc02aa1n12x5               g128(.a(\a[19] ), .b(\b[18] ), .out0(new_n224));
  xorc02aa1n06x5               g129(.a(\a[20] ), .b(\b[19] ), .out0(new_n225));
  aoi112aa1n02x5               g130(.a(new_n223), .b(new_n225), .c(new_n220), .d(new_n224), .o1(new_n226));
  inv030aa1n02x5               g131(.a(new_n223), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n219), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n224), .b(new_n228), .c(new_n205), .d(new_n215), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[19] ), .b(\a[20] ), .out0(new_n230));
  aoi012aa1n03x5               g135(.a(new_n230), .b(new_n229), .c(new_n227), .o1(new_n231));
  nor002aa1n02x5               g136(.a(new_n231), .b(new_n226), .o1(\s[20] ));
  nanp02aa1n02x5               g137(.a(new_n225), .b(new_n224), .o1(new_n233));
  norb02aa1n06x5               g138(.a(new_n215), .b(new_n233), .out0(new_n234));
  inv000aa1n02x5               g139(.a(new_n234), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[18] ), .b(\a[19] ), .out0(new_n236));
  oao003aa1n02x5               g141(.a(\a[20] ), .b(\b[19] ), .c(new_n227), .carry(new_n237));
  oai013aa1d12x5               g142(.a(new_n237), .b(new_n236), .c(new_n230), .d(new_n219), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  aoai13aa1n02x5               g144(.a(new_n239), .b(new_n235), .c(new_n214), .d(new_n204), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  nand02aa1d06x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  nor002aa1d32x5               g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  nand02aa1n06x5               g151(.a(\b[21] ), .b(\a[22] ), .o1(new_n247));
  nanb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(new_n242), .b(new_n249), .c(new_n240), .d(new_n245), .o1(new_n250));
  inv020aa1n04x5               g155(.a(new_n242), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n245), .b(new_n238), .c(new_n205), .d(new_n234), .o1(new_n252));
  aoi012aa1n03x5               g157(.a(new_n248), .b(new_n252), .c(new_n251), .o1(new_n253));
  norp02aa1n03x5               g158(.a(new_n253), .b(new_n250), .o1(\s[22] ));
  nona23aa1n12x5               g159(.a(new_n247), .b(new_n243), .c(new_n242), .d(new_n246), .out0(new_n255));
  nona32aa1n03x5               g160(.a(new_n215), .b(new_n255), .c(new_n230), .d(new_n236), .out0(new_n256));
  nano23aa1n06x5               g161(.a(new_n242), .b(new_n246), .c(new_n247), .d(new_n243), .out0(new_n257));
  oaoi03aa1n02x5               g162(.a(\a[22] ), .b(\b[21] ), .c(new_n251), .o1(new_n258));
  tech160nm_fiaoi012aa1n05x5   g163(.a(new_n258), .b(new_n238), .c(new_n257), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n256), .c(new_n214), .d(new_n204), .o1(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1d32x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  nand42aa1n20x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  norb02aa1n12x5               g168(.a(new_n263), .b(new_n262), .out0(new_n264));
  xorc02aa1n12x5               g169(.a(\a[24] ), .b(\b[23] ), .out0(new_n265));
  aoi112aa1n02x5               g170(.a(new_n262), .b(new_n265), .c(new_n260), .d(new_n264), .o1(new_n266));
  inv000aa1n02x5               g171(.a(new_n262), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n256), .o1(new_n268));
  inv000aa1n02x5               g173(.a(new_n259), .o1(new_n269));
  aoai13aa1n03x5               g174(.a(new_n264), .b(new_n269), .c(new_n205), .d(new_n268), .o1(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[23] ), .b(\a[24] ), .out0(new_n271));
  aoi012aa1n03x5               g176(.a(new_n271), .b(new_n270), .c(new_n267), .o1(new_n272));
  nor002aa1n02x5               g177(.a(new_n272), .b(new_n266), .o1(\s[24] ));
  nano22aa1n03x7               g178(.a(new_n256), .b(new_n264), .c(new_n265), .out0(new_n274));
  inv020aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nanb03aa1n03x5               g180(.a(new_n219), .b(new_n225), .c(new_n224), .out0(new_n276));
  nand03aa1n02x5               g181(.a(new_n257), .b(new_n264), .c(new_n265), .o1(new_n277));
  oaoi03aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .o1(new_n278));
  aoi013aa1n03x5               g183(.a(new_n278), .b(new_n258), .c(new_n265), .d(new_n264), .o1(new_n279));
  aoai13aa1n06x5               g184(.a(new_n279), .b(new_n277), .c(new_n276), .d(new_n237), .o1(new_n280));
  inv040aa1n03x5               g185(.a(new_n280), .o1(new_n281));
  aoai13aa1n02x7               g186(.a(new_n281), .b(new_n275), .c(new_n214), .d(new_n204), .o1(new_n282));
  xorb03aa1n02x5               g187(.a(new_n282), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  tech160nm_fixorc02aa1n03p5x5 g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  xorc02aa1n12x5               g190(.a(\a[26] ), .b(\b[25] ), .out0(new_n286));
  aoi112aa1n02x5               g191(.a(new_n284), .b(new_n286), .c(new_n282), .d(new_n285), .o1(new_n287));
  inv000aa1n02x5               g192(.a(new_n284), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n285), .b(new_n280), .c(new_n205), .d(new_n274), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n286), .o1(new_n290));
  aoi012aa1n03x5               g195(.a(new_n290), .b(new_n289), .c(new_n288), .o1(new_n291));
  nor002aa1n02x5               g196(.a(new_n291), .b(new_n287), .o1(\s[26] ));
  oabi12aa1n02x5               g197(.a(new_n203), .b(new_n162), .c(new_n212), .out0(new_n293));
  and002aa1n02x7               g198(.a(new_n286), .b(new_n285), .o(new_n294));
  nano32aa1n03x7               g199(.a(new_n256), .b(new_n294), .c(new_n264), .d(new_n265), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n293), .c(new_n127), .d(new_n213), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[26] ), .b(\b[25] ), .c(new_n288), .carry(new_n297));
  aobi12aa1n06x5               g202(.a(new_n297), .b(new_n280), .c(new_n294), .out0(new_n298));
  xnrc02aa1n12x5               g203(.a(\b[26] ), .b(\a[27] ), .out0(new_n299));
  xobna2aa1n03x5               g204(.a(new_n299), .b(new_n296), .c(new_n298), .out0(\s[27] ));
  and002aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  xorc02aa1n06x5               g207(.a(\a[28] ), .b(\b[27] ), .out0(new_n303));
  nano22aa1n02x4               g208(.a(new_n255), .b(new_n265), .c(new_n264), .out0(new_n304));
  nand02aa1n02x5               g209(.a(new_n238), .b(new_n304), .o1(new_n305));
  inv000aa1n02x5               g210(.a(new_n294), .o1(new_n306));
  aoai13aa1n09x5               g211(.a(new_n297), .b(new_n306), .c(new_n305), .d(new_n279), .o1(new_n307));
  nor042aa1n03x5               g212(.a(\b[26] ), .b(\a[27] ), .o1(new_n308));
  aoi112aa1n03x4               g213(.a(new_n307), .b(new_n308), .c(new_n205), .d(new_n295), .o1(new_n309));
  nano22aa1n03x5               g214(.a(new_n309), .b(new_n302), .c(new_n303), .out0(new_n310));
  inv000aa1n03x5               g215(.a(new_n308), .o1(new_n311));
  nanp03aa1n02x5               g216(.a(new_n296), .b(new_n298), .c(new_n311), .o1(new_n312));
  aoi012aa1n02x5               g217(.a(new_n303), .b(new_n312), .c(new_n302), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n313), .b(new_n310), .o1(\s[28] ));
  norb02aa1n02x5               g219(.a(new_n303), .b(new_n299), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n307), .c(new_n205), .d(new_n295), .o1(new_n316));
  oao003aa1n03x5               g221(.a(\a[28] ), .b(\b[27] ), .c(new_n311), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[28] ), .b(\a[29] ), .out0(new_n318));
  aoi012aa1n03x5               g223(.a(new_n318), .b(new_n316), .c(new_n317), .o1(new_n319));
  aobi12aa1n02x5               g224(.a(new_n315), .b(new_n296), .c(new_n298), .out0(new_n320));
  nano22aa1n02x4               g225(.a(new_n320), .b(new_n317), .c(new_n318), .out0(new_n321));
  nor002aa1n02x5               g226(.a(new_n319), .b(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g228(.a(new_n303), .b(new_n299), .c(new_n318), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n307), .c(new_n205), .d(new_n295), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .c(new_n317), .carry(new_n326));
  xnrc02aa1n02x5               g231(.a(\b[29] ), .b(\a[30] ), .out0(new_n327));
  aoi012aa1n03x5               g232(.a(new_n327), .b(new_n325), .c(new_n326), .o1(new_n328));
  aobi12aa1n02x5               g233(.a(new_n324), .b(new_n296), .c(new_n298), .out0(new_n329));
  nano22aa1n02x4               g234(.a(new_n329), .b(new_n326), .c(new_n327), .out0(new_n330));
  nor002aa1n02x5               g235(.a(new_n328), .b(new_n330), .o1(\s[30] ));
  nona22aa1n02x4               g236(.a(new_n315), .b(new_n318), .c(new_n327), .out0(new_n332));
  aoi012aa1n02x5               g237(.a(new_n332), .b(new_n296), .c(new_n298), .o1(new_n333));
  oao003aa1n02x5               g238(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n334));
  xnrc02aa1n02x5               g239(.a(\b[30] ), .b(\a[31] ), .out0(new_n335));
  nano22aa1n02x4               g240(.a(new_n333), .b(new_n334), .c(new_n335), .out0(new_n336));
  inv000aa1n02x5               g241(.a(new_n332), .o1(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n307), .c(new_n205), .d(new_n295), .o1(new_n338));
  aoi012aa1n03x5               g243(.a(new_n335), .b(new_n338), .c(new_n334), .o1(new_n339));
  nor002aa1n02x5               g244(.a(new_n339), .b(new_n336), .o1(\s[31] ));
  xnbna2aa1n03x5               g245(.a(new_n102), .b(new_n105), .c(new_n110), .out0(\s[3] ));
  oaoi03aa1n02x5               g246(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n342));
  xorb03aa1n02x5               g247(.a(new_n342), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g248(.a(new_n169), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanp02aa1n02x5               g249(.a(\b[4] ), .b(\a[5] ), .o1(new_n345));
  oai013aa1n02x5               g250(.a(new_n345), .b(new_n151), .c(new_n111), .d(new_n123), .o1(new_n346));
  xorb03aa1n02x5               g251(.a(new_n346), .b(\b[5] ), .c(new_n121), .out0(\s[6] ));
  oaoi03aa1n03x5               g252(.a(\a[6] ), .b(\b[5] ), .c(new_n346), .o1(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n03x5               g254(.a(new_n115), .b(new_n348), .c(new_n116), .o1(new_n350));
  xnrb03aa1n03x5               g255(.a(new_n350), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g256(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


