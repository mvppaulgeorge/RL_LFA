// Benchmark "adder" written by ABC on Thu Jul 18 11:50:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n345, new_n346, new_n348, new_n349, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n357, new_n358, new_n359, new_n361, new_n362,
    new_n364, new_n365, new_n366, new_n368;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nand02aa1d28x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nor042aa1d18x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand02aa1d28x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor042aa1d18x5               g006(.a(new_n100), .b(new_n101), .o1(new_n102));
  nand42aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano23aa1n09x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .d(new_n99), .out0(new_n105));
  oai022aa1n04x7               g010(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n106));
  nand42aa1n16x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nor042aa1d18x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  tech160nm_fiaoi012aa1n03p5x5 g013(.a(new_n108), .b(\a[5] ), .c(\b[4] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  aoi012aa1n06x5               g015(.a(new_n110), .b(\a[4] ), .c(\b[3] ), .o1(new_n111));
  nand02aa1d16x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nanp02aa1n24x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor022aa1n16x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nona23aa1n09x5               g020(.a(new_n114), .b(new_n112), .c(new_n115), .d(new_n113), .out0(new_n116));
  nano32aa1n03x7               g021(.a(new_n116), .b(new_n111), .c(new_n109), .d(new_n107), .out0(new_n117));
  oai012aa1n12x5               g022(.a(new_n117), .b(new_n105), .c(new_n106), .o1(new_n118));
  nano22aa1n03x7               g023(.a(new_n108), .b(new_n107), .c(new_n114), .out0(new_n119));
  oai022aa1d18x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  norb02aa1n06x5               g025(.a(new_n112), .b(new_n110), .out0(new_n121));
  aoi012aa1n06x5               g026(.a(new_n108), .b(new_n110), .c(new_n107), .o1(new_n122));
  inv020aa1n02x5               g027(.a(new_n122), .o1(new_n123));
  aoi013aa1n06x4               g028(.a(new_n123), .b(new_n119), .c(new_n121), .d(new_n120), .o1(new_n124));
  xnrc02aa1n12x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n98), .b(new_n125), .c(new_n118), .d(new_n124), .o1(new_n126));
  nor002aa1d32x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand02aa1d24x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n15x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nand22aa1n03x5               g034(.a(new_n118), .b(new_n124), .o1(new_n130));
  inv000aa1d42x5               g035(.a(new_n125), .o1(new_n131));
  aoi112aa1n02x5               g036(.a(new_n129), .b(new_n97), .c(new_n130), .d(new_n131), .o1(new_n132));
  aoi012aa1n02x5               g037(.a(new_n132), .b(new_n126), .c(new_n129), .o1(\s[10] ));
  oaoi03aa1n02x5               g038(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanp02aa1n09x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  aoai13aa1n06x5               g042(.a(new_n137), .b(new_n134), .c(new_n126), .d(new_n129), .o1(new_n138));
  aoi112aa1n02x5               g043(.a(new_n137), .b(new_n134), .c(new_n126), .d(new_n129), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n138), .b(new_n139), .out0(\s[11] ));
  nor002aa1d32x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand02aa1d28x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  aoib12aa1n02x5               g048(.a(new_n135), .b(new_n142), .c(new_n141), .out0(new_n144));
  tech160nm_fioai012aa1n03p5x5 g049(.a(new_n138), .b(\b[10] ), .c(\a[11] ), .o1(new_n145));
  aboi22aa1n03x5               g050(.a(new_n143), .b(new_n145), .c(new_n138), .d(new_n144), .out0(\s[12] ));
  nanb03aa1n12x5               g051(.a(new_n104), .b(new_n99), .c(new_n103), .out0(new_n147));
  oab012aa1n09x5               g052(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .out0(new_n148));
  aoai13aa1n12x5               g053(.a(new_n148), .b(new_n147), .c(new_n99), .d(new_n102), .o1(new_n149));
  nand23aa1n03x5               g054(.a(new_n119), .b(new_n121), .c(new_n120), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n150), .b(new_n122), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(\b[8] ), .b(\a[9] ), .o1(new_n152));
  nona23aa1n09x5               g057(.a(new_n142), .b(new_n136), .c(new_n135), .d(new_n141), .out0(new_n153));
  nano32aa1n03x7               g058(.a(new_n153), .b(new_n129), .c(new_n152), .d(new_n98), .out0(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n151), .c(new_n149), .d(new_n117), .o1(new_n155));
  nano22aa1n03x7               g060(.a(new_n141), .b(new_n136), .c(new_n142), .out0(new_n156));
  oai012aa1n04x7               g061(.a(new_n128), .b(\b[10] ), .c(\a[11] ), .o1(new_n157));
  oab012aa1n06x5               g062(.a(new_n157), .b(new_n97), .c(new_n127), .out0(new_n158));
  tech160nm_fiaoi012aa1n05x5   g063(.a(new_n141), .b(new_n135), .c(new_n142), .o1(new_n159));
  aob012aa1n02x5               g064(.a(new_n159), .b(new_n158), .c(new_n156), .out0(new_n160));
  nanb02aa1n03x5               g065(.a(new_n160), .b(new_n155), .out0(new_n161));
  nor002aa1d32x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanp02aa1n24x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  inv020aa1n03x5               g069(.a(new_n159), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n164), .c(new_n158), .d(new_n156), .o1(new_n166));
  aoi022aa1n02x5               g071(.a(new_n161), .b(new_n164), .c(new_n155), .d(new_n166), .o1(\s[13] ));
  nor022aa1n12x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand42aa1n16x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  aoi112aa1n02x7               g075(.a(new_n162), .b(new_n170), .c(new_n161), .d(new_n164), .o1(new_n171));
  aoai13aa1n02x5               g076(.a(new_n170), .b(new_n162), .c(new_n161), .d(new_n163), .o1(new_n172));
  norb02aa1n03x4               g077(.a(new_n172), .b(new_n171), .out0(\s[14] ));
  nano23aa1d15x5               g078(.a(new_n162), .b(new_n168), .c(new_n169), .d(new_n163), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n160), .c(new_n130), .d(new_n154), .o1(new_n175));
  oai012aa1n12x5               g080(.a(new_n169), .b(new_n168), .c(new_n162), .o1(new_n176));
  nor002aa1d32x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand02aa1d06x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n175), .c(new_n176), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(new_n176), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n180), .b(new_n182), .c(new_n161), .d(new_n174), .o1(new_n183));
  nor022aa1n16x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand22aa1n09x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nanb02aa1n02x5               g090(.a(new_n184), .b(new_n185), .out0(new_n186));
  aoib12aa1n02x5               g091(.a(new_n177), .b(new_n185), .c(new_n184), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n177), .o1(new_n188));
  aoai13aa1n02x7               g093(.a(new_n188), .b(new_n179), .c(new_n175), .d(new_n176), .o1(new_n189));
  aboi22aa1n03x5               g094(.a(new_n186), .b(new_n189), .c(new_n183), .d(new_n187), .out0(\s[16] ));
  nona23aa1d18x5               g095(.a(new_n185), .b(new_n178), .c(new_n177), .d(new_n184), .out0(new_n191));
  inv020aa1n02x5               g096(.a(new_n191), .o1(new_n192));
  nand23aa1n03x5               g097(.a(new_n154), .b(new_n174), .c(new_n192), .o1(new_n193));
  aoi012aa1n12x5               g098(.a(new_n193), .b(new_n118), .c(new_n124), .o1(new_n194));
  aoai13aa1n04x5               g099(.a(new_n174), .b(new_n165), .c(new_n158), .d(new_n156), .o1(new_n195));
  tech160nm_fiaoi012aa1n03p5x5 g100(.a(new_n184), .b(new_n177), .c(new_n185), .o1(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n191), .c(new_n195), .d(new_n176), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  tech160nm_fioai012aa1n03p5x5 g103(.a(new_n198), .b(new_n197), .c(new_n194), .o1(new_n199));
  aob012aa1n02x5               g104(.a(new_n192), .b(new_n195), .c(new_n176), .out0(new_n200));
  nano23aa1n02x4               g105(.a(new_n198), .b(new_n194), .c(new_n200), .d(new_n196), .out0(new_n201));
  norb02aa1n02x5               g106(.a(new_n199), .b(new_n201), .out0(\s[17] ));
  nor002aa1d32x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  nor002aa1n16x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nand22aa1n09x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  norb02aa1n06x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n199), .c(new_n204), .out0(\s[18] ));
  and002aa1n02x5               g113(.a(new_n198), .b(new_n207), .o(new_n209));
  oaih12aa1n02x5               g114(.a(new_n209), .b(new_n197), .c(new_n194), .o1(new_n210));
  oaoi03aa1n09x5               g115(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor042aa1d18x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand02aa1d16x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n12x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n210), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fiaoi012aa1n05x5   g122(.a(new_n151), .b(new_n149), .c(new_n117), .o1(new_n218));
  oai112aa1n06x5               g123(.a(new_n200), .b(new_n196), .c(new_n218), .d(new_n193), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n215), .b(new_n211), .c(new_n219), .d(new_n209), .o1(new_n220));
  nor002aa1n20x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1d28x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1n03x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  inv000aa1d42x5               g128(.a(\a[19] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\b[18] ), .o1(new_n225));
  aboi22aa1n03x5               g130(.a(new_n221), .b(new_n222), .c(new_n224), .d(new_n225), .out0(new_n226));
  inv030aa1n03x5               g131(.a(new_n213), .o1(new_n227));
  inv030aa1n02x5               g132(.a(new_n215), .o1(new_n228));
  aoai13aa1n02x7               g133(.a(new_n227), .b(new_n228), .c(new_n210), .d(new_n212), .o1(new_n229));
  aoi022aa1n03x5               g134(.a(new_n229), .b(new_n223), .c(new_n220), .d(new_n226), .o1(\s[20] ));
  nano32aa1n03x7               g135(.a(new_n228), .b(new_n198), .c(new_n223), .d(new_n207), .out0(new_n231));
  oaih12aa1n02x5               g136(.a(new_n231), .b(new_n197), .c(new_n194), .o1(new_n232));
  nanb03aa1n12x5               g137(.a(new_n221), .b(new_n222), .c(new_n214), .out0(new_n233));
  oai112aa1n06x5               g138(.a(new_n227), .b(new_n206), .c(new_n205), .d(new_n203), .o1(new_n234));
  aoi012aa1n06x5               g139(.a(new_n221), .b(new_n213), .c(new_n222), .o1(new_n235));
  oai012aa1d24x5               g140(.a(new_n235), .b(new_n234), .c(new_n233), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[20] ), .b(\a[21] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n236), .c(new_n219), .d(new_n231), .o1(new_n239));
  nano22aa1n02x5               g144(.a(new_n221), .b(new_n214), .c(new_n222), .out0(new_n240));
  oai012aa1n02x5               g145(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .o1(new_n241));
  oab012aa1n02x4               g146(.a(new_n241), .b(new_n203), .c(new_n205), .out0(new_n242));
  inv000aa1n02x5               g147(.a(new_n235), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(new_n238), .b(new_n243), .c(new_n242), .d(new_n240), .o1(new_n244));
  aobi12aa1n02x7               g149(.a(new_n239), .b(new_n244), .c(new_n232), .out0(\s[21] ));
  xnrc02aa1n12x5               g150(.a(\b[21] ), .b(\a[22] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  nor042aa1n03x5               g152(.a(\b[20] ), .b(\a[21] ), .o1(new_n248));
  norb02aa1n02x5               g153(.a(new_n246), .b(new_n248), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n236), .o1(new_n250));
  inv000aa1n03x5               g155(.a(new_n248), .o1(new_n251));
  aoai13aa1n02x7               g156(.a(new_n251), .b(new_n237), .c(new_n232), .d(new_n250), .o1(new_n252));
  aoi022aa1n03x5               g157(.a(new_n252), .b(new_n247), .c(new_n239), .d(new_n249), .o1(\s[22] ));
  nor042aa1n06x5               g158(.a(new_n246), .b(new_n237), .o1(new_n254));
  and002aa1n02x5               g159(.a(new_n231), .b(new_n254), .o(new_n255));
  oaih12aa1n02x5               g160(.a(new_n255), .b(new_n197), .c(new_n194), .o1(new_n256));
  oao003aa1n02x5               g161(.a(\a[22] ), .b(\b[21] ), .c(new_n251), .carry(new_n257));
  inv030aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(new_n236), .c(new_n254), .o1(new_n259));
  inv040aa1n03x5               g164(.a(new_n259), .o1(new_n260));
  xorc02aa1n12x5               g165(.a(\a[23] ), .b(\b[22] ), .out0(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n260), .c(new_n219), .d(new_n255), .o1(new_n262));
  aoi112aa1n02x5               g167(.a(new_n261), .b(new_n258), .c(new_n236), .d(new_n254), .o1(new_n263));
  aobi12aa1n02x7               g168(.a(new_n262), .b(new_n263), .c(new_n256), .out0(\s[23] ));
  xorc02aa1n03x5               g169(.a(\a[24] ), .b(\b[23] ), .out0(new_n265));
  nor042aa1n09x5               g170(.a(\b[22] ), .b(\a[23] ), .o1(new_n266));
  norp02aa1n02x5               g171(.a(new_n265), .b(new_n266), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n266), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n261), .o1(new_n269));
  aoai13aa1n02x7               g174(.a(new_n268), .b(new_n269), .c(new_n256), .d(new_n259), .o1(new_n270));
  aoi022aa1n03x5               g175(.a(new_n270), .b(new_n265), .c(new_n262), .d(new_n267), .o1(\s[24] ));
  inv030aa1n02x5               g176(.a(new_n231), .o1(new_n272));
  and002aa1n06x5               g177(.a(new_n265), .b(new_n261), .o(new_n273));
  nano22aa1n06x5               g178(.a(new_n272), .b(new_n273), .c(new_n254), .out0(new_n274));
  oaih12aa1n02x5               g179(.a(new_n274), .b(new_n197), .c(new_n194), .o1(new_n275));
  aoai13aa1n06x5               g180(.a(new_n254), .b(new_n243), .c(new_n242), .d(new_n240), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n273), .o1(new_n277));
  oao003aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .c(new_n268), .carry(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n276), .d(new_n257), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[25] ), .b(\b[24] ), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n279), .c(new_n219), .d(new_n274), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n273), .b(new_n258), .c(new_n236), .d(new_n254), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n280), .o1(new_n283));
  and003aa1n02x5               g188(.a(new_n282), .b(new_n283), .c(new_n278), .o(new_n284));
  aobi12aa1n02x7               g189(.a(new_n281), .b(new_n284), .c(new_n275), .out0(\s[25] ));
  tech160nm_fixorc02aa1n03p5x5 g190(.a(\a[26] ), .b(\b[25] ), .out0(new_n286));
  nor042aa1n06x5               g191(.a(\b[24] ), .b(\a[25] ), .o1(new_n287));
  norp02aa1n02x5               g192(.a(new_n286), .b(new_n287), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n279), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n287), .o1(new_n290));
  aoai13aa1n02x7               g195(.a(new_n290), .b(new_n283), .c(new_n275), .d(new_n289), .o1(new_n291));
  aoi022aa1n03x5               g196(.a(new_n291), .b(new_n286), .c(new_n281), .d(new_n288), .o1(\s[26] ));
  and002aa1n12x5               g197(.a(new_n286), .b(new_n280), .o(new_n293));
  nano32aa1d15x5               g198(.a(new_n272), .b(new_n293), .c(new_n254), .d(new_n273), .out0(new_n294));
  oai012aa1n12x5               g199(.a(new_n294), .b(new_n197), .c(new_n194), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n293), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[26] ), .b(\b[25] ), .c(new_n290), .carry(new_n297));
  aoai13aa1n04x5               g202(.a(new_n297), .b(new_n296), .c(new_n282), .d(new_n278), .o1(new_n298));
  xorc02aa1n12x5               g203(.a(\a[27] ), .b(\b[26] ), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n298), .c(new_n219), .d(new_n294), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n297), .o1(new_n301));
  aoi112aa1n02x5               g206(.a(new_n299), .b(new_n301), .c(new_n279), .d(new_n293), .o1(new_n302));
  aobi12aa1n02x7               g207(.a(new_n300), .b(new_n302), .c(new_n295), .out0(\s[27] ));
  xorc02aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .out0(new_n304));
  norp02aa1n02x5               g209(.a(\b[26] ), .b(\a[27] ), .o1(new_n305));
  norp02aa1n02x5               g210(.a(new_n304), .b(new_n305), .o1(new_n306));
  tech160nm_fiaoi012aa1n04x5   g211(.a(new_n301), .b(new_n279), .c(new_n293), .o1(new_n307));
  inv000aa1n03x5               g212(.a(new_n305), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n299), .o1(new_n309));
  aoai13aa1n02x7               g214(.a(new_n308), .b(new_n309), .c(new_n307), .d(new_n295), .o1(new_n310));
  aoi022aa1n03x5               g215(.a(new_n310), .b(new_n304), .c(new_n300), .d(new_n306), .o1(\s[28] ));
  and002aa1n02x5               g216(.a(new_n304), .b(new_n299), .o(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n298), .c(new_n219), .d(new_n294), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n312), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[28] ), .b(\b[27] ), .c(new_n308), .carry(new_n315));
  aoai13aa1n04x5               g220(.a(new_n315), .b(new_n314), .c(new_n307), .d(new_n295), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  norb02aa1n02x5               g222(.a(new_n315), .b(new_n317), .out0(new_n318));
  aoi022aa1n02x7               g223(.a(new_n316), .b(new_n317), .c(new_n313), .d(new_n318), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g225(.a(new_n309), .b(new_n304), .c(new_n317), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n298), .c(new_n219), .d(new_n294), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n321), .o1(new_n323));
  inv000aa1d42x5               g228(.a(\b[28] ), .o1(new_n324));
  inv000aa1d42x5               g229(.a(\a[29] ), .o1(new_n325));
  oaib12aa1n02x5               g230(.a(new_n315), .b(\b[28] ), .c(new_n325), .out0(new_n326));
  oaib12aa1n02x5               g231(.a(new_n326), .b(new_n324), .c(\a[29] ), .out0(new_n327));
  aoai13aa1n02x7               g232(.a(new_n327), .b(new_n323), .c(new_n307), .d(new_n295), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[30] ), .b(\b[29] ), .out0(new_n329));
  oaoi13aa1n02x5               g234(.a(new_n329), .b(new_n326), .c(new_n325), .d(new_n324), .o1(new_n330));
  aoi022aa1n03x5               g235(.a(new_n328), .b(new_n329), .c(new_n322), .d(new_n330), .o1(\s[30] ));
  nanb02aa1n02x5               g236(.a(\b[30] ), .b(\a[31] ), .out0(new_n332));
  nanb02aa1n02x5               g237(.a(\a[31] ), .b(\b[30] ), .out0(new_n333));
  nanp02aa1n02x5               g238(.a(new_n333), .b(new_n332), .o1(new_n334));
  nano32aa1n03x7               g239(.a(new_n309), .b(new_n329), .c(new_n304), .d(new_n317), .out0(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n298), .c(new_n219), .d(new_n294), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n335), .o1(new_n337));
  norp02aa1n02x5               g242(.a(\b[29] ), .b(\a[30] ), .o1(new_n338));
  aoi022aa1n02x5               g243(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n339));
  aoi012aa1n02x5               g244(.a(new_n338), .b(new_n326), .c(new_n339), .o1(new_n340));
  aoai13aa1n02x7               g245(.a(new_n340), .b(new_n337), .c(new_n307), .d(new_n295), .o1(new_n341));
  oai112aa1n02x5               g246(.a(new_n332), .b(new_n333), .c(\b[29] ), .d(\a[30] ), .o1(new_n342));
  aoi012aa1n02x5               g247(.a(new_n342), .b(new_n326), .c(new_n339), .o1(new_n343));
  aoi022aa1n03x5               g248(.a(new_n341), .b(new_n334), .c(new_n336), .d(new_n343), .o1(\s[31] ));
  inv000aa1d42x5               g249(.a(new_n102), .o1(new_n345));
  aboi22aa1n03x5               g250(.a(new_n104), .b(new_n103), .c(new_n345), .d(new_n99), .out0(new_n346));
  norp02aa1n02x5               g251(.a(new_n346), .b(new_n105), .o1(\s[3] ));
  xorc02aa1n02x5               g252(.a(\a[4] ), .b(\b[3] ), .out0(new_n348));
  norp02aa1n02x5               g253(.a(new_n348), .b(new_n104), .o1(new_n349));
  aboi22aa1n03x5               g254(.a(new_n105), .b(new_n349), .c(new_n149), .d(new_n348), .out0(\s[4] ));
  and002aa1n02x5               g255(.a(\b[4] ), .b(\a[5] ), .o(new_n351));
  aoi112aa1n02x5               g256(.a(new_n351), .b(new_n115), .c(\a[4] ), .d(\b[3] ), .o1(new_n352));
  xnrc02aa1n02x5               g257(.a(\b[4] ), .b(\a[5] ), .out0(new_n353));
  and002aa1n02x5               g258(.a(\b[3] ), .b(\a[4] ), .o(new_n354));
  oabi12aa1n02x5               g259(.a(new_n354), .b(new_n105), .c(new_n106), .out0(new_n355));
  aoi022aa1n02x5               g260(.a(new_n355), .b(new_n353), .c(new_n149), .d(new_n352), .o1(\s[5] ));
  norb02aa1n02x5               g261(.a(new_n114), .b(new_n113), .out0(new_n357));
  aoai13aa1n02x5               g262(.a(new_n357), .b(new_n115), .c(new_n149), .d(new_n352), .o1(new_n358));
  aoi112aa1n02x5               g263(.a(new_n115), .b(new_n357), .c(new_n149), .d(new_n352), .o1(new_n359));
  norb02aa1n02x5               g264(.a(new_n358), .b(new_n359), .out0(\s[6] ));
  oai012aa1n02x5               g265(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n361));
  nand23aa1n03x5               g266(.a(new_n149), .b(new_n352), .c(new_n357), .o1(new_n362));
  xnbna2aa1n03x5               g267(.a(new_n121), .b(new_n362), .c(new_n361), .out0(\s[7] ));
  inv000aa1d42x5               g268(.a(new_n110), .o1(new_n364));
  aob012aa1n02x5               g269(.a(new_n121), .b(new_n362), .c(new_n361), .out0(new_n365));
  norb02aa1n02x5               g270(.a(new_n107), .b(new_n108), .out0(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n366), .b(new_n365), .c(new_n364), .out0(\s[8] ));
  aoi113aa1n02x5               g272(.a(new_n123), .b(new_n131), .c(new_n119), .d(new_n121), .e(new_n120), .o1(new_n368));
  aoi022aa1n02x5               g273(.a(new_n130), .b(new_n131), .c(new_n118), .d(new_n368), .o1(\s[9] ));
endmodule


