// Benchmark "adder" written by ABC on Thu Jul 18 09:56:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n324,
    new_n325, new_n326, new_n327, new_n330, new_n332, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[3] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[4] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[2] ), .o1(new_n99));
  aboi22aa1n03x5               g004(.a(\b[3] ), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n100));
  xnrc02aa1n02x5               g005(.a(\b[2] ), .b(\a[3] ), .out0(new_n101));
  nanp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor042aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  tech160nm_fioai012aa1n03p5x5 g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  oai012aa1n12x5               g010(.a(new_n100), .b(new_n101), .c(new_n105), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[7] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[6] ), .o1(new_n109));
  nand02aa1d04x5               g014(.a(new_n109), .b(new_n108), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nanp03aa1n02x5               g016(.a(new_n110), .b(new_n107), .c(new_n111), .o1(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .out0(new_n113));
  nor022aa1n16x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nanp02aa1n03x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor022aa1n08x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nona23aa1n02x4               g022(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n118));
  nor043aa1n06x5               g023(.a(new_n118), .b(new_n113), .c(new_n112), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[8] ), .o1(new_n120));
  nanb02aa1n02x5               g025(.a(\b[7] ), .b(new_n120), .out0(new_n121));
  oaih12aa1n06x5               g026(.a(new_n115), .b(new_n116), .c(new_n114), .o1(new_n122));
  aob012aa1n02x5               g027(.a(new_n107), .b(\b[7] ), .c(\a[8] ), .out0(new_n123));
  aoai13aa1n12x5               g028(.a(new_n121), .b(new_n123), .c(new_n122), .d(new_n110), .o1(new_n124));
  aoi012aa1d18x5               g029(.a(new_n124), .b(new_n119), .c(new_n106), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[9] ), .b(\b[8] ), .c(new_n125), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  tech160nm_finand02aa1n05x5   g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  and002aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o(new_n129));
  xnrc02aa1n12x5               g034(.a(\b[8] ), .b(\a[9] ), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  nor022aa1n04x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  norb02aa1n03x5               g037(.a(new_n128), .b(new_n132), .out0(new_n133));
  aoai13aa1n03x5               g038(.a(new_n133), .b(new_n129), .c(new_n125), .d(new_n131), .o1(new_n134));
  xnrc02aa1n02x5               g039(.a(\b[10] ), .b(\a[11] ), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n134), .c(new_n128), .out0(\s[11] ));
  orn002aa1n02x5               g041(.a(\a[11] ), .b(\b[10] ), .o(new_n137));
  xorc02aa1n12x5               g042(.a(\a[11] ), .b(\b[10] ), .out0(new_n138));
  nanp03aa1n03x5               g043(.a(new_n134), .b(new_n128), .c(new_n138), .o1(new_n139));
  xorc02aa1n02x5               g044(.a(\a[12] ), .b(\b[11] ), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n139), .c(new_n137), .out0(\s[12] ));
  xnrc02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .out0(new_n142));
  nano23aa1n02x5               g047(.a(new_n130), .b(new_n142), .c(new_n138), .d(new_n133), .out0(new_n143));
  aoai13aa1n06x5               g048(.a(new_n143), .b(new_n124), .c(new_n119), .d(new_n106), .o1(new_n144));
  norp02aa1n02x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  inv000aa1n02x5               g050(.a(new_n145), .o1(new_n146));
  tech160nm_fiao0012aa1n02p5x5 g051(.a(new_n137), .b(\a[12] ), .c(\b[11] ), .o(new_n147));
  norp02aa1n02x5               g052(.a(\b[8] ), .b(\a[9] ), .o1(new_n148));
  oai012aa1n02x5               g053(.a(new_n128), .b(new_n132), .c(new_n148), .o1(new_n149));
  norp03aa1n02x5               g054(.a(new_n135), .b(new_n142), .c(new_n149), .o1(new_n150));
  nano22aa1n02x4               g055(.a(new_n150), .b(new_n147), .c(new_n146), .out0(new_n151));
  xorc02aa1n12x5               g056(.a(\a[13] ), .b(\b[12] ), .out0(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n144), .c(new_n151), .out0(\s[13] ));
  nona23aa1n02x4               g058(.a(new_n138), .b(new_n133), .c(new_n142), .d(new_n130), .out0(new_n154));
  norp02aa1n02x5               g059(.a(new_n125), .b(new_n154), .o1(new_n155));
  nanb03aa1n02x5               g060(.a(new_n149), .b(new_n138), .c(new_n140), .out0(new_n156));
  nand03aa1n02x5               g061(.a(new_n156), .b(new_n146), .c(new_n147), .o1(new_n157));
  norp02aa1n02x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  oaoi13aa1n03x5               g063(.a(new_n158), .b(new_n152), .c(new_n155), .d(new_n157), .o1(new_n159));
  xnrb03aa1n02x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nanp02aa1n02x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nor002aa1n04x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nanb02aa1n12x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n152), .o1(new_n165));
  oai022aa1d24x5               g070(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n04x5               g072(.a(new_n167), .b(new_n165), .c(new_n144), .d(new_n151), .o1(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n164), .b(new_n168), .c(new_n161), .out0(\s[15] ));
  nano22aa1n02x4               g074(.a(new_n163), .b(new_n161), .c(new_n162), .out0(new_n170));
  tech160nm_fixorc02aa1n04x5   g075(.a(\a[16] ), .b(\b[15] ), .out0(new_n171));
  aoi112aa1n02x5               g076(.a(new_n171), .b(new_n163), .c(new_n168), .d(new_n170), .o1(new_n172));
  aoai13aa1n02x5               g077(.a(new_n171), .b(new_n163), .c(new_n168), .d(new_n170), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(\s[16] ));
  xnrc02aa1n02x5               g079(.a(\b[13] ), .b(\a[14] ), .out0(new_n175));
  nona23aa1n06x5               g080(.a(new_n171), .b(new_n152), .c(new_n175), .d(new_n164), .out0(new_n176));
  nor042aa1n03x5               g081(.a(new_n154), .b(new_n176), .o1(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n124), .c(new_n106), .d(new_n119), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nano23aa1n09x5               g084(.a(new_n164), .b(new_n175), .c(new_n171), .d(new_n152), .out0(new_n180));
  aoai13aa1n06x5               g085(.a(new_n162), .b(new_n163), .c(new_n166), .d(new_n161), .o1(new_n181));
  oai012aa1n02x5               g086(.a(new_n181), .b(\b[15] ), .c(\a[16] ), .o1(new_n182));
  aoi022aa1n12x5               g087(.a(new_n157), .b(new_n180), .c(new_n179), .d(new_n182), .o1(new_n183));
  xorc02aa1n12x5               g088(.a(\a[17] ), .b(\b[16] ), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n178), .c(new_n183), .out0(\s[17] ));
  nano22aa1n02x4               g090(.a(new_n125), .b(new_n180), .c(new_n143), .out0(new_n186));
  nanp02aa1n02x5               g091(.a(new_n182), .b(new_n179), .o1(new_n187));
  tech160nm_fioai012aa1n04x5   g092(.a(new_n187), .b(new_n151), .c(new_n176), .o1(new_n188));
  norp02aa1n02x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  oaoi13aa1n03x5               g094(.a(new_n189), .b(new_n184), .c(new_n186), .d(new_n188), .o1(new_n190));
  xnrb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n02x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nand42aa1n04x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  inv040aa1d32x5               g098(.a(\a[19] ), .o1(new_n194));
  inv040aa1d30x5               g099(.a(\b[18] ), .o1(new_n195));
  nand02aa1d08x5               g100(.a(new_n195), .b(new_n194), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n184), .o1(new_n197));
  oai022aa1d24x5               g102(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n197), .c(new_n178), .d(new_n183), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n200), .b(new_n192), .c(new_n193), .d(new_n196), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(new_n180), .b(new_n143), .o1(new_n202));
  oai012aa1n18x5               g107(.a(new_n183), .b(new_n202), .c(new_n125), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n196), .o1(new_n204));
  nano22aa1n02x4               g109(.a(new_n204), .b(new_n192), .c(new_n193), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n198), .c(new_n203), .d(new_n184), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n09x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand42aa1n06x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  tech160nm_fiaoi012aa1n05x5   g117(.a(new_n212), .b(new_n206), .c(new_n196), .o1(new_n213));
  aoi112aa1n03x4               g118(.a(new_n211), .b(new_n204), .c(new_n200), .d(new_n205), .o1(new_n214));
  nor042aa1n03x5               g119(.a(new_n213), .b(new_n214), .o1(\s[20] ));
  xnrc02aa1n02x5               g120(.a(\b[17] ), .b(\a[18] ), .out0(new_n216));
  nanb03aa1n12x5               g121(.a(new_n209), .b(new_n210), .c(new_n193), .out0(new_n217));
  nano23aa1n06x5               g122(.a(new_n217), .b(new_n216), .c(new_n184), .d(new_n196), .out0(new_n218));
  inv020aa1n02x5               g123(.a(new_n218), .o1(new_n219));
  nand23aa1n04x5               g124(.a(new_n198), .b(new_n196), .c(new_n192), .o1(new_n220));
  aoai13aa1n12x5               g125(.a(new_n210), .b(new_n209), .c(new_n194), .d(new_n195), .o1(new_n221));
  oai012aa1d24x5               g126(.a(new_n221), .b(new_n220), .c(new_n217), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n04x5               g128(.a(new_n223), .b(new_n219), .c(new_n178), .d(new_n183), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  xnrc02aa1n12x5               g133(.a(\b[21] ), .b(\a[22] ), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoi112aa1n02x5               g135(.a(new_n226), .b(new_n230), .c(new_n224), .d(new_n228), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n226), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n228), .b(new_n222), .c(new_n203), .d(new_n218), .o1(new_n233));
  tech160nm_fiaoi012aa1n02p5x5 g138(.a(new_n229), .b(new_n233), .c(new_n232), .o1(new_n234));
  norp02aa1n02x5               g139(.a(new_n234), .b(new_n231), .o1(\s[22] ));
  nor022aa1n08x5               g140(.a(new_n229), .b(new_n227), .o1(new_n236));
  nand22aa1n12x5               g141(.a(new_n218), .b(new_n236), .o1(new_n237));
  oaoi03aa1n09x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n232), .o1(new_n238));
  aoi012aa1n09x5               g143(.a(new_n238), .b(new_n222), .c(new_n236), .o1(new_n239));
  aoai13aa1n04x5               g144(.a(new_n239), .b(new_n237), .c(new_n178), .d(new_n183), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n04x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  and002aa1n06x5               g147(.a(\b[22] ), .b(\a[23] ), .o(new_n243));
  nor002aa1n02x5               g148(.a(new_n243), .b(new_n242), .o1(new_n244));
  tech160nm_fixorc02aa1n03p5x5 g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoi112aa1n03x4               g150(.a(new_n242), .b(new_n245), .c(new_n240), .d(new_n244), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n242), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n237), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n239), .o1(new_n249));
  aoai13aa1n03x5               g154(.a(new_n244), .b(new_n249), .c(new_n203), .d(new_n248), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n245), .o1(new_n251));
  tech160nm_fiaoi012aa1n02p5x5 g156(.a(new_n251), .b(new_n250), .c(new_n247), .o1(new_n252));
  nor002aa1n02x5               g157(.a(new_n252), .b(new_n246), .o1(\s[24] ));
  inv000aa1d42x5               g158(.a(new_n124), .o1(new_n254));
  aob012aa1n06x5               g159(.a(new_n254), .b(new_n119), .c(new_n106), .out0(new_n255));
  nano32aa1n06x5               g160(.a(new_n219), .b(new_n245), .c(new_n236), .d(new_n244), .out0(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n188), .c(new_n255), .d(new_n177), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n243), .o1(new_n258));
  aoai13aa1n09x5               g163(.a(new_n258), .b(new_n238), .c(new_n222), .d(new_n236), .o1(new_n259));
  oab012aa1n09x5               g164(.a(new_n242), .b(\a[24] ), .c(\b[23] ), .out0(new_n260));
  aoi022aa1n06x5               g165(.a(new_n259), .b(new_n260), .c(\b[23] ), .d(\a[24] ), .o1(new_n261));
  inv000aa1n06x5               g166(.a(new_n261), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[24] ), .b(\a[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n262), .c(new_n257), .out0(\s[25] ));
  orn002aa1n02x5               g170(.a(\a[25] ), .b(\b[24] ), .o(new_n266));
  aoai13aa1n06x5               g171(.a(new_n264), .b(new_n261), .c(new_n203), .d(new_n256), .o1(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  aoi012aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n266), .o1(new_n269));
  tech160nm_fiaoi012aa1n05x5   g174(.a(new_n263), .b(new_n262), .c(new_n257), .o1(new_n270));
  nano22aa1n03x5               g175(.a(new_n270), .b(new_n266), .c(new_n268), .out0(new_n271));
  nor002aa1n02x5               g176(.a(new_n269), .b(new_n271), .o1(\s[26] ));
  and002aa1n02x5               g177(.a(\b[23] ), .b(\a[24] ), .o(new_n273));
  nor043aa1d12x5               g178(.a(new_n268), .b(new_n263), .c(new_n273), .o1(new_n274));
  nano32aa1d12x5               g179(.a(new_n237), .b(new_n274), .c(new_n244), .d(new_n245), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n188), .c(new_n255), .d(new_n177), .o1(new_n276));
  nano22aa1n02x4               g181(.a(new_n209), .b(new_n193), .c(new_n210), .out0(new_n277));
  oai012aa1n02x5               g182(.a(new_n192), .b(\b[18] ), .c(\a[19] ), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n198), .b(new_n278), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n221), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n236), .b(new_n280), .c(new_n279), .d(new_n277), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n238), .o1(new_n282));
  aoai13aa1n02x5               g187(.a(new_n260), .b(new_n243), .c(new_n281), .d(new_n282), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .c(new_n266), .carry(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n283), .c(new_n274), .out0(new_n285));
  xorc02aa1n02x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n276), .out0(\s[27] ));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv040aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  aobi12aa1n02x7               g194(.a(new_n286), .b(new_n285), .c(new_n276), .out0(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  nano22aa1n03x5               g196(.a(new_n290), .b(new_n289), .c(new_n291), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n274), .o1(new_n293));
  aoai13aa1n12x5               g198(.a(new_n284), .b(new_n293), .c(new_n259), .d(new_n260), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n286), .b(new_n294), .c(new_n203), .d(new_n275), .o1(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n291), .b(new_n295), .c(new_n289), .o1(new_n296));
  norp02aa1n03x5               g201(.a(new_n296), .b(new_n292), .o1(\s[28] ));
  norb02aa1n02x5               g202(.a(new_n286), .b(new_n291), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n294), .c(new_n203), .d(new_n275), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[28] ), .b(\a[29] ), .out0(new_n301));
  tech160nm_fiaoi012aa1n02p5x5 g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  aobi12aa1n02x7               g207(.a(new_n298), .b(new_n285), .c(new_n276), .out0(new_n303));
  nano22aa1n03x5               g208(.a(new_n303), .b(new_n300), .c(new_n301), .out0(new_n304));
  norp02aa1n03x5               g209(.a(new_n302), .b(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g211(.a(new_n286), .b(new_n301), .c(new_n291), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n294), .c(new_n203), .d(new_n275), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[29] ), .b(\a[30] ), .out0(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n310), .b(new_n308), .c(new_n309), .o1(new_n311));
  aobi12aa1n02x7               g216(.a(new_n307), .b(new_n285), .c(new_n276), .out0(new_n312));
  nano22aa1n03x5               g217(.a(new_n312), .b(new_n309), .c(new_n310), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[30] ));
  norb02aa1n02x5               g219(.a(new_n307), .b(new_n310), .out0(new_n315));
  aoai13aa1n02x5               g220(.a(new_n315), .b(new_n294), .c(new_n203), .d(new_n275), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n318), .b(new_n316), .c(new_n317), .o1(new_n319));
  aobi12aa1n02x7               g224(.a(new_n315), .b(new_n285), .c(new_n276), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n320), .b(new_n317), .c(new_n318), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[31] ));
  xorb03aa1n02x5               g227(.a(new_n105), .b(\b[2] ), .c(new_n97), .out0(\s[3] ));
  and002aa1n02x5               g228(.a(new_n106), .b(new_n111), .o(new_n324));
  norp02aa1n02x5               g229(.a(new_n101), .b(new_n105), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[4] ), .b(\b[3] ), .out0(new_n326));
  aoi112aa1n02x5               g231(.a(new_n325), .b(new_n326), .c(new_n97), .d(new_n99), .o1(new_n327));
  oaoi13aa1n02x5               g232(.a(new_n327), .b(new_n324), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g233(.a(new_n324), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi013aa1n02x4               g234(.a(new_n116), .b(new_n106), .c(new_n111), .d(new_n117), .o1(new_n330));
  xnrb03aa1n02x5               g235(.a(new_n330), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g236(.a(\a[6] ), .b(\b[5] ), .c(new_n330), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g238(.a(new_n108), .b(new_n109), .c(new_n332), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[7] ), .c(new_n120), .out0(\s[8] ));
  xnrc02aa1n02x5               g240(.a(new_n125), .b(new_n131), .out0(\s[9] ));
endmodule


