// Benchmark "adder" written by ABC on Thu Jul 18 01:04:50 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n340, new_n341, new_n343, new_n345, new_n346, new_n347,
    new_n348, new_n351;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n06x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aoi012aa1n09x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  inv040aa1d32x5               g008(.a(\a[4] ), .o1(new_n104));
  inv000aa1d42x5               g009(.a(\b[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nand42aa1n03x5               g012(.a(new_n106), .b(new_n107), .o1(new_n108));
  inv040aa1d32x5               g013(.a(\a[3] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(new_n111), .b(new_n112), .o1(new_n113));
  nor003aa1n03x5               g018(.a(new_n103), .b(new_n108), .c(new_n113), .o1(new_n114));
  nor042aa1n09x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  oaoi03aa1n09x5               g020(.a(new_n104), .b(new_n105), .c(new_n115), .o1(new_n116));
  inv000aa1n02x5               g021(.a(new_n116), .o1(new_n117));
  nor022aa1n16x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nand42aa1n08x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor002aa1n16x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nona23aa1n06x5               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  nor042aa1n04x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  nanp02aa1n04x5               g028(.a(\b[7] ), .b(\a[8] ), .o1(new_n124));
  nor042aa1n04x5               g029(.a(\b[6] ), .b(\a[7] ), .o1(new_n125));
  nanp02aa1n04x5               g030(.a(\b[6] ), .b(\a[7] ), .o1(new_n126));
  nona23aa1n02x4               g031(.a(new_n126), .b(new_n124), .c(new_n123), .d(new_n125), .out0(new_n127));
  nor002aa1n02x5               g032(.a(new_n127), .b(new_n122), .o1(new_n128));
  tech160nm_fioai012aa1n05x5   g033(.a(new_n128), .b(new_n114), .c(new_n117), .o1(new_n129));
  nano23aa1n09x5               g034(.a(new_n123), .b(new_n125), .c(new_n126), .d(new_n124), .out0(new_n130));
  oa0012aa1n12x5               g035(.a(new_n119), .b(new_n120), .c(new_n118), .o(new_n131));
  tech160nm_fiao0012aa1n02p5x5 g036(.a(new_n123), .b(new_n125), .c(new_n124), .o(new_n132));
  aoi012aa1d24x5               g037(.a(new_n132), .b(new_n130), .c(new_n131), .o1(new_n133));
  xorc02aa1n12x5               g038(.a(\a[9] ), .b(\b[8] ), .out0(new_n134));
  inv000aa1d42x5               g039(.a(new_n134), .o1(new_n135));
  aoai13aa1n02x5               g040(.a(new_n99), .b(new_n135), .c(new_n129), .d(new_n133), .o1(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xorc02aa1n02x5               g042(.a(\a[4] ), .b(\b[3] ), .out0(new_n138));
  norb02aa1n02x5               g043(.a(new_n112), .b(new_n115), .out0(new_n139));
  nanb03aa1n06x5               g044(.a(new_n103), .b(new_n138), .c(new_n139), .out0(new_n140));
  nano23aa1n02x4               g045(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n141));
  nand02aa1n02x5               g046(.a(new_n130), .b(new_n141), .o1(new_n142));
  aoai13aa1n12x5               g047(.a(new_n133), .b(new_n142), .c(new_n140), .d(new_n116), .o1(new_n143));
  nanp02aa1n03x5               g048(.a(new_n143), .b(new_n134), .o1(new_n144));
  nor002aa1d32x5               g049(.a(\b[9] ), .b(\a[10] ), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  nand42aa1n06x5               g051(.a(\b[9] ), .b(\a[10] ), .o1(new_n147));
  norb02aa1n12x5               g052(.a(new_n147), .b(new_n145), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n146), .b(new_n149), .c(new_n144), .d(new_n99), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n06x5               g056(.a(\b[10] ), .b(\a[11] ), .o1(new_n152));
  nand02aa1d04x5               g057(.a(\b[10] ), .b(\a[11] ), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  nor042aa1n04x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand02aa1n04x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n03x5               g063(.a(new_n158), .b(new_n152), .c(new_n150), .d(new_n154), .o1(new_n159));
  aoai13aa1n02x5               g064(.a(new_n154), .b(new_n145), .c(new_n136), .d(new_n147), .o1(new_n160));
  nona22aa1n02x4               g065(.a(new_n160), .b(new_n158), .c(new_n152), .out0(new_n161));
  nanp02aa1n02x5               g066(.a(new_n159), .b(new_n161), .o1(\s[12] ));
  nona23aa1n09x5               g067(.a(new_n156), .b(new_n153), .c(new_n152), .d(new_n155), .out0(new_n163));
  nano22aa1n12x5               g068(.a(new_n163), .b(new_n134), .c(new_n148), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nano23aa1n09x5               g070(.a(new_n152), .b(new_n155), .c(new_n156), .d(new_n153), .out0(new_n166));
  aoai13aa1n09x5               g071(.a(new_n147), .b(new_n145), .c(new_n97), .d(new_n98), .o1(new_n167));
  inv000aa1n02x5               g072(.a(new_n167), .o1(new_n168));
  tech160nm_fiaoi012aa1n03p5x5 g073(.a(new_n155), .b(new_n152), .c(new_n156), .o1(new_n169));
  aobi12aa1n12x5               g074(.a(new_n169), .b(new_n166), .c(new_n168), .out0(new_n170));
  aoai13aa1n03x5               g075(.a(new_n170), .b(new_n165), .c(new_n129), .d(new_n133), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d24x5               g077(.a(\b[12] ), .b(\a[13] ), .o1(new_n173));
  nanp02aa1n02x5               g078(.a(\b[12] ), .b(\a[13] ), .o1(new_n174));
  aoi012aa1n02x5               g079(.a(new_n173), .b(new_n171), .c(new_n174), .o1(new_n175));
  xnrb03aa1n03x5               g080(.a(new_n175), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  tech160nm_fioai012aa1n03p5x5 g081(.a(new_n169), .b(new_n163), .c(new_n167), .o1(new_n177));
  nor002aa1d32x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nand02aa1n04x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nona23aa1n03x5               g084(.a(new_n179), .b(new_n174), .c(new_n173), .d(new_n178), .out0(new_n180));
  inv040aa1n03x5               g085(.a(new_n180), .o1(new_n181));
  aoai13aa1n03x5               g086(.a(new_n181), .b(new_n177), .c(new_n143), .d(new_n164), .o1(new_n182));
  oai012aa1n12x5               g087(.a(new_n179), .b(new_n178), .c(new_n173), .o1(new_n183));
  norp02aa1n04x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  nand42aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n182), .c(new_n183), .out0(\s[15] ));
  nanp02aa1n03x5               g092(.a(new_n182), .b(new_n183), .o1(new_n188));
  norp02aa1n04x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  nand42aa1n02x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nanb02aa1n02x5               g095(.a(new_n189), .b(new_n190), .out0(new_n191));
  aoai13aa1n03x5               g096(.a(new_n191), .b(new_n184), .c(new_n188), .d(new_n186), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n183), .o1(new_n193));
  aoai13aa1n02x5               g098(.a(new_n186), .b(new_n193), .c(new_n171), .d(new_n181), .o1(new_n194));
  nona22aa1n02x4               g099(.a(new_n194), .b(new_n191), .c(new_n184), .out0(new_n195));
  nanp02aa1n03x5               g100(.a(new_n192), .b(new_n195), .o1(\s[16] ));
  nona23aa1n09x5               g101(.a(new_n190), .b(new_n185), .c(new_n184), .d(new_n189), .out0(new_n197));
  nor002aa1n02x5               g102(.a(new_n197), .b(new_n180), .o1(new_n198));
  nand42aa1n02x5               g103(.a(new_n164), .b(new_n198), .o1(new_n199));
  aoi012aa1n02x5               g104(.a(new_n189), .b(new_n184), .c(new_n190), .o1(new_n200));
  tech160nm_fioai012aa1n04x5   g105(.a(new_n200), .b(new_n197), .c(new_n183), .o1(new_n201));
  tech160nm_fiaoi012aa1n03p5x5 g106(.a(new_n201), .b(new_n177), .c(new_n198), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n129), .d(new_n133), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d28x5               g109(.a(\a[17] ), .o1(new_n205));
  inv040aa1d32x5               g110(.a(\b[16] ), .o1(new_n206));
  oaoi03aa1n03x5               g111(.a(new_n205), .b(new_n206), .c(new_n203), .o1(new_n207));
  xnrb03aa1n03x5               g112(.a(new_n207), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanb02aa1n12x5               g113(.a(new_n197), .b(new_n181), .out0(new_n209));
  nano32aa1n03x7               g114(.a(new_n209), .b(new_n166), .c(new_n148), .d(new_n134), .out0(new_n210));
  oabi12aa1n18x5               g115(.a(new_n201), .b(new_n209), .c(new_n170), .out0(new_n211));
  nor002aa1n02x5               g116(.a(\b[16] ), .b(\a[17] ), .o1(new_n212));
  nand42aa1n03x5               g117(.a(\b[16] ), .b(\a[17] ), .o1(new_n213));
  nor002aa1d32x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  nand42aa1d28x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  nano23aa1n06x5               g120(.a(new_n212), .b(new_n214), .c(new_n215), .d(new_n213), .out0(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n211), .c(new_n143), .d(new_n210), .o1(new_n217));
  aoai13aa1n12x5               g122(.a(new_n215), .b(new_n214), .c(new_n205), .d(new_n206), .o1(new_n218));
  xorc02aa1n12x5               g123(.a(\a[19] ), .b(\b[18] ), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n218), .out0(\s[19] ));
  xnrc02aa1n02x5               g125(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g126(.a(new_n217), .b(new_n218), .o1(new_n222));
  norp02aa1n02x5               g127(.a(\b[18] ), .b(\a[19] ), .o1(new_n223));
  tech160nm_fixnrc02aa1n04x5   g128(.a(\b[19] ), .b(\a[20] ), .out0(new_n224));
  aoai13aa1n03x5               g129(.a(new_n224), .b(new_n223), .c(new_n222), .d(new_n219), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n218), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n219), .b(new_n226), .c(new_n203), .d(new_n216), .o1(new_n227));
  nona22aa1n02x4               g132(.a(new_n227), .b(new_n224), .c(new_n223), .out0(new_n228));
  nanp02aa1n03x5               g133(.a(new_n225), .b(new_n228), .o1(\s[20] ));
  xorc02aa1n06x5               g134(.a(\a[20] ), .b(\b[19] ), .out0(new_n230));
  nand23aa1n04x5               g135(.a(new_n216), .b(new_n219), .c(new_n230), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n211), .c(new_n143), .d(new_n210), .o1(new_n233));
  tech160nm_fixnrc02aa1n02p5x5 g138(.a(\b[18] ), .b(\a[19] ), .out0(new_n234));
  orn002aa1n02x5               g139(.a(\a[19] ), .b(\b[18] ), .o(new_n235));
  oao003aa1n02x5               g140(.a(\a[20] ), .b(\b[19] ), .c(new_n235), .carry(new_n236));
  oai013aa1d12x5               g141(.a(new_n236), .b(new_n234), .c(new_n224), .d(new_n218), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  nor022aa1n08x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  nand42aa1n03x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  nanb02aa1n06x5               g145(.a(new_n239), .b(new_n240), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  xnbna2aa1n03x5               g147(.a(new_n242), .b(new_n233), .c(new_n238), .out0(\s[21] ));
  nanp02aa1n02x5               g148(.a(new_n233), .b(new_n238), .o1(new_n244));
  nor002aa1n06x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  nanp02aa1n02x5               g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  nanb02aa1n02x5               g151(.a(new_n245), .b(new_n246), .out0(new_n247));
  aoai13aa1n03x5               g152(.a(new_n247), .b(new_n239), .c(new_n244), .d(new_n242), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n242), .b(new_n237), .c(new_n203), .d(new_n232), .o1(new_n249));
  nona22aa1n02x4               g154(.a(new_n249), .b(new_n247), .c(new_n239), .out0(new_n250));
  nanp02aa1n02x5               g155(.a(new_n248), .b(new_n250), .o1(\s[22] ));
  nona23aa1n03x5               g156(.a(new_n246), .b(new_n240), .c(new_n239), .d(new_n245), .out0(new_n252));
  nano32aa1n02x4               g157(.a(new_n252), .b(new_n216), .c(new_n219), .d(new_n230), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n211), .c(new_n143), .d(new_n210), .o1(new_n254));
  inv040aa1n02x5               g159(.a(new_n252), .o1(new_n255));
  oai012aa1n03x5               g160(.a(new_n246), .b(new_n245), .c(new_n239), .o1(new_n256));
  inv020aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  tech160nm_fiaoi012aa1n04x5   g162(.a(new_n257), .b(new_n237), .c(new_n255), .o1(new_n258));
  nor042aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  norb02aa1n02x5               g165(.a(new_n260), .b(new_n259), .out0(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n254), .c(new_n258), .out0(\s[23] ));
  tech160nm_finand02aa1n03p5x5 g167(.a(new_n254), .b(new_n258), .o1(new_n263));
  nor042aa1n02x5               g168(.a(\b[23] ), .b(\a[24] ), .o1(new_n264));
  nanp02aa1n02x5               g169(.a(\b[23] ), .b(\a[24] ), .o1(new_n265));
  nanb02aa1n02x5               g170(.a(new_n264), .b(new_n265), .out0(new_n266));
  aoai13aa1n02x5               g171(.a(new_n266), .b(new_n259), .c(new_n263), .d(new_n261), .o1(new_n267));
  inv040aa1n03x5               g172(.a(new_n258), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n261), .b(new_n268), .c(new_n203), .d(new_n253), .o1(new_n269));
  nona22aa1n02x5               g174(.a(new_n269), .b(new_n266), .c(new_n259), .out0(new_n270));
  nanp02aa1n03x5               g175(.a(new_n267), .b(new_n270), .o1(\s[24] ));
  nano23aa1n03x7               g176(.a(new_n259), .b(new_n264), .c(new_n265), .d(new_n260), .out0(new_n272));
  nano22aa1n03x7               g177(.a(new_n231), .b(new_n255), .c(new_n272), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n211), .c(new_n143), .d(new_n210), .o1(new_n274));
  nanb03aa1n03x5               g179(.a(new_n218), .b(new_n230), .c(new_n219), .out0(new_n275));
  nona22aa1n03x5               g180(.a(new_n272), .b(new_n247), .c(new_n241), .out0(new_n276));
  oai012aa1n02x5               g181(.a(new_n265), .b(new_n264), .c(new_n259), .o1(new_n277));
  aobi12aa1n06x5               g182(.a(new_n277), .b(new_n272), .c(new_n257), .out0(new_n278));
  aoai13aa1n04x5               g183(.a(new_n278), .b(new_n276), .c(new_n275), .d(new_n236), .o1(new_n279));
  inv000aa1n02x5               g184(.a(new_n279), .o1(new_n280));
  tech160nm_finand02aa1n03p5x5 g185(.a(new_n274), .b(new_n280), .o1(new_n281));
  tech160nm_fixorc02aa1n03p5x5 g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  nona23aa1n02x4               g187(.a(new_n265), .b(new_n260), .c(new_n259), .d(new_n264), .out0(new_n283));
  norp02aa1n02x5               g188(.a(new_n283), .b(new_n252), .o1(new_n284));
  oai012aa1n02x5               g189(.a(new_n277), .b(new_n283), .c(new_n256), .o1(new_n285));
  aoi112aa1n02x5               g190(.a(new_n282), .b(new_n285), .c(new_n237), .d(new_n284), .o1(new_n286));
  aoi022aa1n02x5               g191(.a(new_n281), .b(new_n282), .c(new_n274), .d(new_n286), .o1(\s[25] ));
  norp02aa1n02x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[25] ), .b(\a[26] ), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n288), .c(new_n281), .d(new_n282), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n282), .b(new_n279), .c(new_n203), .d(new_n273), .o1(new_n291));
  nona22aa1n02x4               g196(.a(new_n291), .b(new_n289), .c(new_n288), .out0(new_n292));
  nanp02aa1n02x5               g197(.a(new_n290), .b(new_n292), .o1(\s[26] ));
  norb02aa1n02x5               g198(.a(new_n282), .b(new_n289), .out0(new_n294));
  nano32aa1n03x7               g199(.a(new_n231), .b(new_n294), .c(new_n255), .d(new_n272), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n211), .c(new_n143), .d(new_n210), .o1(new_n296));
  aoi112aa1n02x5               g201(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n297));
  oab012aa1n02x4               g202(.a(new_n297), .b(\a[26] ), .c(\b[25] ), .out0(new_n298));
  aobi12aa1n06x5               g203(.a(new_n298), .b(new_n279), .c(new_n294), .out0(new_n299));
  xorc02aa1n02x5               g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  xnbna2aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n299), .out0(\s[27] ));
  nand42aa1n03x5               g206(.a(new_n296), .b(new_n299), .o1(new_n302));
  norp02aa1n02x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  norp02aa1n02x5               g208(.a(\b[27] ), .b(\a[28] ), .o1(new_n304));
  nanp02aa1n02x5               g209(.a(\b[27] ), .b(\a[28] ), .o1(new_n305));
  norb02aa1n06x4               g210(.a(new_n305), .b(new_n304), .out0(new_n306));
  inv000aa1d42x5               g211(.a(new_n306), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n302), .d(new_n300), .o1(new_n308));
  aoai13aa1n06x5               g213(.a(new_n294), .b(new_n285), .c(new_n237), .d(new_n284), .o1(new_n309));
  tech160nm_finand02aa1n05x5   g214(.a(new_n309), .b(new_n298), .o1(new_n310));
  aoai13aa1n06x5               g215(.a(new_n300), .b(new_n310), .c(new_n203), .d(new_n295), .o1(new_n311));
  nona22aa1n02x5               g216(.a(new_n311), .b(new_n307), .c(new_n303), .out0(new_n312));
  nanp02aa1n03x5               g217(.a(new_n308), .b(new_n312), .o1(\s[28] ));
  norb02aa1n02x5               g218(.a(new_n300), .b(new_n307), .out0(new_n314));
  aoai13aa1n06x5               g219(.a(new_n314), .b(new_n310), .c(new_n203), .d(new_n295), .o1(new_n315));
  oai012aa1n02x5               g220(.a(new_n305), .b(new_n304), .c(new_n303), .o1(new_n316));
  tech160nm_finand02aa1n03p5x5 g221(.a(new_n315), .b(new_n316), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n316), .b(new_n318), .out0(new_n319));
  aoi022aa1n02x7               g224(.a(new_n317), .b(new_n318), .c(new_n315), .d(new_n319), .o1(\s[29] ));
  xorb03aa1n02x5               g225(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g226(.a(new_n318), .b(new_n300), .c(new_n306), .o1(new_n322));
  nanb02aa1n03x5               g227(.a(new_n322), .b(new_n302), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .carry(new_n324));
  aoai13aa1n02x7               g229(.a(new_n324), .b(new_n322), .c(new_n296), .d(new_n299), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .out0(new_n326));
  norp02aa1n02x5               g231(.a(\b[28] ), .b(\a[29] ), .o1(new_n327));
  aoi012aa1n02x5               g232(.a(new_n316), .b(\a[29] ), .c(\b[28] ), .o1(new_n328));
  norp03aa1n02x5               g233(.a(new_n328), .b(new_n326), .c(new_n327), .o1(new_n329));
  aoi022aa1n03x5               g234(.a(new_n329), .b(new_n323), .c(new_n325), .d(new_n326), .o1(\s[30] ));
  norb02aa1n02x5               g235(.a(new_n326), .b(new_n322), .out0(new_n331));
  aoai13aa1n06x5               g236(.a(new_n331), .b(new_n310), .c(new_n203), .d(new_n295), .o1(new_n332));
  oao003aa1n02x5               g237(.a(\a[30] ), .b(\b[29] ), .c(new_n324), .carry(new_n333));
  xnrc02aa1n02x5               g238(.a(\b[30] ), .b(\a[31] ), .out0(new_n334));
  tech160nm_fiaoi012aa1n03p5x5 g239(.a(new_n334), .b(new_n332), .c(new_n333), .o1(new_n335));
  aobi12aa1n02x7               g240(.a(new_n331), .b(new_n296), .c(new_n299), .out0(new_n336));
  nano22aa1n02x4               g241(.a(new_n336), .b(new_n333), .c(new_n334), .out0(new_n337));
  nor002aa1n02x5               g242(.a(new_n335), .b(new_n337), .o1(\s[31] ));
  xnbna2aa1n03x5               g243(.a(new_n103), .b(new_n112), .c(new_n111), .out0(\s[3] ));
  nanp02aa1n02x5               g244(.a(new_n108), .b(new_n111), .o1(new_n340));
  oab012aa1n02x4               g245(.a(new_n340), .b(new_n103), .c(new_n113), .out0(new_n341));
  oaoi13aa1n02x5               g246(.a(new_n341), .b(new_n106), .c(new_n114), .d(new_n117), .o1(\s[4] ));
  nanb02aa1n02x5               g247(.a(new_n120), .b(new_n121), .out0(new_n343));
  xobna2aa1n03x5               g248(.a(new_n343), .b(new_n140), .c(new_n116), .out0(\s[5] ));
  oabi12aa1n02x5               g249(.a(new_n343), .b(new_n114), .c(new_n117), .out0(new_n345));
  aoib12aa1n02x5               g250(.a(new_n120), .b(new_n119), .c(new_n118), .out0(new_n346));
  inv000aa1d42x5               g251(.a(new_n131), .o1(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n122), .c(new_n140), .d(new_n116), .o1(new_n348));
  aboi22aa1n03x5               g253(.a(new_n118), .b(new_n348), .c(new_n345), .d(new_n346), .out0(\s[6] ));
  xorb03aa1n02x5               g254(.a(new_n348), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g255(.a(new_n125), .b(new_n348), .c(new_n126), .o1(new_n351));
  xnrb03aa1n02x5               g256(.a(new_n351), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g257(.a(new_n134), .b(new_n129), .c(new_n133), .out0(\s[9] ));
endmodule


