// Benchmark "adder" written by ABC on Wed Jul 17 18:47:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n353, new_n355, new_n357, new_n359, new_n360, new_n361,
    new_n363, new_n364, new_n366, new_n367, new_n368;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[8] ), .o1(new_n97));
  nanb02aa1n03x5               g002(.a(\a[9] ), .b(new_n97), .out0(new_n98));
  nor002aa1n03x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  inv020aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aob012aa1n03x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  nor002aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand42aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n03x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor042aa1n06x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nand23aa1n04x5               g014(.a(new_n103), .b(new_n106), .c(new_n109), .o1(new_n110));
  tech160nm_fiaoi012aa1n05x5   g015(.a(new_n104), .b(new_n107), .c(new_n105), .o1(new_n111));
  nor042aa1n09x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor042aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano23aa1n03x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nor042aa1n03x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand02aa1d08x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nor042aa1d18x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nand02aa1n04x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nano23aa1n02x5               g025(.a(new_n117), .b(new_n119), .c(new_n120), .d(new_n118), .out0(new_n121));
  nand22aa1n03x5               g026(.a(new_n121), .b(new_n116), .o1(new_n122));
  norb02aa1n06x4               g027(.a(new_n118), .b(new_n117), .out0(new_n123));
  nano22aa1n03x7               g028(.a(new_n119), .b(new_n113), .c(new_n120), .out0(new_n124));
  oai022aa1n02x5               g029(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n125));
  inv040aa1n02x5               g030(.a(new_n119), .o1(new_n126));
  oaoi03aa1n09x5               g031(.a(\a[8] ), .b(\b[7] ), .c(new_n126), .o1(new_n127));
  aoi013aa1n06x4               g032(.a(new_n127), .b(new_n124), .c(new_n125), .d(new_n123), .o1(new_n128));
  aoai13aa1n12x5               g033(.a(new_n128), .b(new_n122), .c(new_n110), .d(new_n111), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  nanp02aa1n03x5               g035(.a(new_n129), .b(new_n130), .o1(new_n131));
  xorc02aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n131), .c(new_n98), .out0(\s[10] ));
  nand02aa1d12x5               g038(.a(new_n132), .b(new_n130), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n134), .o1(new_n135));
  tech160nm_fioaoi03aa1n03p5x5 g040(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n136));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanp02aa1n06x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n09x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  aoai13aa1n06x5               g044(.a(new_n139), .b(new_n136), .c(new_n129), .d(new_n135), .o1(new_n140));
  aoi112aa1n02x5               g045(.a(new_n139), .b(new_n136), .c(new_n129), .d(new_n135), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(\s[11] ));
  inv000aa1d42x5               g047(.a(new_n137), .o1(new_n143));
  tech160nm_fixorc02aa1n02p5x5 g048(.a(\a[12] ), .b(\b[11] ), .out0(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n140), .c(new_n143), .out0(\s[12] ));
  aoi012aa1n02x5               g050(.a(new_n99), .b(new_n101), .c(new_n102), .o1(new_n146));
  nona23aa1n03x5               g051(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n147));
  tech160nm_fioai012aa1n03p5x5 g052(.a(new_n111), .b(new_n147), .c(new_n146), .o1(new_n148));
  nanb02aa1n06x5               g053(.a(new_n122), .b(new_n148), .out0(new_n149));
  nano22aa1d15x5               g054(.a(new_n134), .b(new_n139), .c(new_n144), .out0(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  inv040aa1d32x5               g056(.a(\a[12] ), .o1(new_n152));
  inv000aa1d42x5               g057(.a(\b[11] ), .o1(new_n153));
  nanp02aa1n03x5               g058(.a(new_n153), .b(new_n152), .o1(new_n154));
  nand22aa1n03x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand23aa1n03x5               g060(.a(new_n154), .b(new_n138), .c(new_n155), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[9] ), .b(\a[10] ), .o1(new_n157));
  oaih22aa1d12x5               g062(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n158));
  oai112aa1n06x5               g063(.a(new_n158), .b(new_n157), .c(\b[10] ), .d(\a[11] ), .o1(new_n159));
  tech160nm_fioaoi03aa1n03p5x5 g064(.a(new_n152), .b(new_n153), .c(new_n137), .o1(new_n160));
  oai012aa1n12x5               g065(.a(new_n160), .b(new_n159), .c(new_n156), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n151), .c(new_n149), .d(new_n128), .o1(new_n163));
  nor042aa1n06x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  norb02aa1n02x7               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  aoi112aa1n02x5               g071(.a(new_n166), .b(new_n161), .c(new_n129), .d(new_n150), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n163), .c(new_n166), .o1(\s[13] ));
  nor042aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1n08x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n06x4               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  aoi112aa1n02x5               g076(.a(new_n164), .b(new_n171), .c(new_n163), .d(new_n166), .o1(new_n172));
  aoai13aa1n02x7               g077(.a(new_n171), .b(new_n164), .c(new_n163), .d(new_n165), .o1(new_n173));
  norb02aa1n02x7               g078(.a(new_n173), .b(new_n172), .out0(\s[14] ));
  nano23aa1n06x5               g079(.a(new_n164), .b(new_n169), .c(new_n170), .d(new_n165), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n161), .c(new_n129), .d(new_n150), .o1(new_n176));
  oai012aa1d24x5               g081(.a(new_n170), .b(new_n169), .c(new_n164), .o1(new_n177));
  xorc02aa1n12x5               g082(.a(\a[15] ), .b(\b[14] ), .out0(new_n178));
  xnbna2aa1n03x5               g083(.a(new_n178), .b(new_n176), .c(new_n177), .out0(\s[15] ));
  inv000aa1d42x5               g084(.a(new_n177), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n178), .b(new_n180), .c(new_n163), .d(new_n175), .o1(new_n181));
  xorc02aa1n02x5               g086(.a(\a[16] ), .b(\b[15] ), .out0(new_n182));
  inv000aa1d42x5               g087(.a(\a[15] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[14] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\a[16] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\b[15] ), .o1(new_n186));
  nanp02aa1n02x5               g091(.a(new_n186), .b(new_n185), .o1(new_n187));
  nanp02aa1n02x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  aoi022aa1n02x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .d(new_n183), .o1(new_n189));
  nor042aa1n02x5               g094(.a(\b[14] ), .b(\a[15] ), .o1(new_n190));
  inv000aa1n02x5               g095(.a(new_n190), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n178), .o1(new_n192));
  aoai13aa1n03x5               g097(.a(new_n191), .b(new_n192), .c(new_n176), .d(new_n177), .o1(new_n193));
  aoi022aa1n03x5               g098(.a(new_n193), .b(new_n182), .c(new_n181), .d(new_n189), .o1(\s[16] ));
  nanp02aa1n02x5               g099(.a(new_n154), .b(new_n155), .o1(new_n195));
  nano22aa1n02x4               g100(.a(new_n195), .b(new_n143), .c(new_n138), .out0(new_n196));
  nand23aa1n03x5               g101(.a(new_n175), .b(new_n178), .c(new_n182), .o1(new_n197));
  nano32aa1n09x5               g102(.a(new_n197), .b(new_n196), .c(new_n132), .d(new_n130), .out0(new_n198));
  nanp02aa1n02x5               g103(.a(new_n129), .b(new_n198), .o1(new_n199));
  nano32aa1n03x7               g104(.a(new_n192), .b(new_n182), .c(new_n166), .d(new_n171), .out0(new_n200));
  nand02aa1d04x5               g105(.a(new_n150), .b(new_n200), .o1(new_n201));
  oai112aa1n02x5               g106(.a(new_n187), .b(new_n188), .c(new_n184), .d(new_n183), .o1(new_n202));
  oai112aa1n03x5               g107(.a(new_n191), .b(new_n170), .c(new_n169), .d(new_n164), .o1(new_n203));
  oaoi03aa1n02x5               g108(.a(new_n185), .b(new_n186), .c(new_n190), .o1(new_n204));
  tech160nm_fioai012aa1n04x5   g109(.a(new_n204), .b(new_n203), .c(new_n202), .o1(new_n205));
  tech160nm_fiaoi012aa1n02p5x5 g110(.a(new_n205), .b(new_n200), .c(new_n161), .o1(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n201), .c(new_n149), .d(new_n128), .o1(new_n207));
  xorc02aa1n02x5               g112(.a(\a[17] ), .b(\b[16] ), .out0(new_n208));
  aoi112aa1n02x5               g113(.a(new_n205), .b(new_n208), .c(new_n200), .d(new_n161), .o1(new_n209));
  aoi022aa1n02x5               g114(.a(new_n207), .b(new_n208), .c(new_n199), .d(new_n209), .o1(\s[17] ));
  inv000aa1d42x5               g115(.a(\a[17] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(\b[16] ), .o1(new_n212));
  nand22aa1n04x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  nanb03aa1n03x5               g118(.a(new_n156), .b(new_n136), .c(new_n143), .out0(new_n214));
  inv020aa1n02x5               g119(.a(new_n205), .o1(new_n215));
  aoai13aa1n12x5               g120(.a(new_n215), .b(new_n197), .c(new_n214), .d(new_n160), .o1(new_n216));
  aoai13aa1n06x5               g121(.a(new_n208), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n217));
  nor022aa1n08x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  nand42aa1n04x5               g123(.a(\b[17] ), .b(\a[18] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  xnbna2aa1n03x5               g125(.a(new_n220), .b(new_n217), .c(new_n213), .out0(\s[18] ));
  nanp02aa1n02x5               g126(.a(\b[16] ), .b(\a[17] ), .o1(new_n222));
  nano32aa1n02x5               g127(.a(new_n218), .b(new_n213), .c(new_n219), .d(new_n222), .out0(new_n223));
  aoai13aa1n06x5               g128(.a(new_n223), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n224));
  aoai13aa1n06x5               g129(.a(new_n219), .b(new_n218), .c(new_n211), .d(new_n212), .o1(new_n225));
  xorc02aa1n12x5               g130(.a(\a[19] ), .b(\b[18] ), .out0(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n224), .c(new_n225), .out0(\s[19] ));
  xnrc02aa1n02x5               g132(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fioaoi03aa1n03p5x5 g133(.a(\a[18] ), .b(\b[17] ), .c(new_n213), .o1(new_n229));
  aoai13aa1n02x7               g134(.a(new_n226), .b(new_n229), .c(new_n207), .d(new_n223), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[20] ), .b(\b[19] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(\a[19] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\b[18] ), .o1(new_n233));
  inv040aa1d32x5               g138(.a(\a[20] ), .o1(new_n234));
  inv040aa1d28x5               g139(.a(\b[19] ), .o1(new_n235));
  nand42aa1n02x5               g140(.a(new_n235), .b(new_n234), .o1(new_n236));
  tech160nm_finand02aa1n05x5   g141(.a(\b[19] ), .b(\a[20] ), .o1(new_n237));
  aoi022aa1n02x5               g142(.a(new_n236), .b(new_n237), .c(new_n233), .d(new_n232), .o1(new_n238));
  nor002aa1n16x5               g143(.a(\b[18] ), .b(\a[19] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n226), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n241), .c(new_n224), .d(new_n225), .o1(new_n242));
  aoi022aa1n03x5               g147(.a(new_n242), .b(new_n231), .c(new_n230), .d(new_n238), .o1(\s[20] ));
  nano32aa1n02x4               g148(.a(new_n241), .b(new_n231), .c(new_n208), .d(new_n220), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n245));
  oai112aa1n06x5               g150(.a(new_n236), .b(new_n237), .c(new_n233), .d(new_n232), .o1(new_n246));
  oaoi03aa1n06x5               g151(.a(new_n234), .b(new_n235), .c(new_n239), .o1(new_n247));
  oai013aa1n09x5               g152(.a(new_n247), .b(new_n246), .c(new_n225), .d(new_n239), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  nor042aa1d18x5               g154(.a(\b[20] ), .b(\a[21] ), .o1(new_n250));
  nanp02aa1n02x5               g155(.a(\b[20] ), .b(\a[21] ), .o1(new_n251));
  norb02aa1n02x5               g156(.a(new_n251), .b(new_n250), .out0(new_n252));
  xnbna2aa1n03x5               g157(.a(new_n252), .b(new_n245), .c(new_n249), .out0(\s[21] ));
  aoai13aa1n03x5               g158(.a(new_n252), .b(new_n248), .c(new_n207), .d(new_n244), .o1(new_n254));
  nor042aa1n04x5               g159(.a(\b[21] ), .b(\a[22] ), .o1(new_n255));
  nanp02aa1n04x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  aoib12aa1n02x5               g162(.a(new_n250), .b(new_n256), .c(new_n255), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n250), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n252), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n259), .b(new_n260), .c(new_n245), .d(new_n249), .o1(new_n261));
  aoi022aa1n03x5               g166(.a(new_n261), .b(new_n257), .c(new_n254), .d(new_n258), .o1(\s[22] ));
  xroi22aa1d04x5               g167(.a(new_n232), .b(\b[18] ), .c(new_n234), .d(\b[19] ), .out0(new_n263));
  nano23aa1n06x5               g168(.a(new_n250), .b(new_n255), .c(new_n256), .d(new_n251), .out0(new_n264));
  and003aa1n02x5               g169(.a(new_n263), .b(new_n223), .c(new_n264), .o(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n266));
  oai022aa1n02x5               g171(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n267));
  aoi022aa1n02x7               g172(.a(new_n248), .b(new_n264), .c(new_n256), .d(new_n267), .o1(new_n268));
  xorc02aa1n12x5               g173(.a(\a[23] ), .b(\b[22] ), .out0(new_n269));
  xnbna2aa1n03x5               g174(.a(new_n269), .b(new_n266), .c(new_n268), .out0(\s[23] ));
  inv040aa1n03x5               g175(.a(new_n268), .o1(new_n271));
  aoai13aa1n02x7               g176(.a(new_n269), .b(new_n271), .c(new_n207), .d(new_n265), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[24] ), .b(\b[23] ), .out0(new_n273));
  inv000aa1d42x5               g178(.a(\a[23] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(\b[22] ), .o1(new_n275));
  orn002aa1n03x5               g180(.a(\a[24] ), .b(\b[23] ), .o(new_n276));
  nand02aa1n03x5               g181(.a(\b[23] ), .b(\a[24] ), .o1(new_n277));
  aoi022aa1n02x5               g182(.a(new_n276), .b(new_n277), .c(new_n275), .d(new_n274), .o1(new_n278));
  nor042aa1n02x5               g183(.a(\b[22] ), .b(\a[23] ), .o1(new_n279));
  inv000aa1n02x5               g184(.a(new_n279), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n269), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n280), .b(new_n281), .c(new_n266), .d(new_n268), .o1(new_n282));
  aoi022aa1n03x5               g187(.a(new_n282), .b(new_n273), .c(new_n272), .d(new_n278), .o1(\s[24] ));
  nand23aa1n06x5               g188(.a(new_n264), .b(new_n269), .c(new_n273), .o1(new_n284));
  nano32aa1n02x4               g189(.a(new_n284), .b(new_n223), .c(new_n226), .d(new_n231), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n286));
  oai022aa1n02x5               g191(.a(new_n232), .b(new_n233), .c(\b[19] ), .d(\a[20] ), .o1(new_n287));
  nona23aa1n06x5               g192(.a(new_n229), .b(new_n237), .c(new_n287), .d(new_n239), .out0(new_n288));
  oai112aa1n04x5               g193(.a(new_n276), .b(new_n277), .c(new_n275), .d(new_n274), .o1(new_n289));
  oai112aa1n02x7               g194(.a(new_n280), .b(new_n256), .c(new_n255), .d(new_n250), .o1(new_n290));
  aob012aa1n02x5               g195(.a(new_n276), .b(new_n279), .c(new_n277), .out0(new_n291));
  oab012aa1n09x5               g196(.a(new_n291), .b(new_n290), .c(new_n289), .out0(new_n292));
  aoai13aa1n12x5               g197(.a(new_n292), .b(new_n284), .c(new_n288), .d(new_n247), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  nanp02aa1n02x5               g199(.a(new_n286), .b(new_n294), .o1(new_n295));
  xorc02aa1n12x5               g200(.a(\a[25] ), .b(\b[24] ), .out0(new_n296));
  nanb02aa1n06x5               g201(.a(new_n284), .b(new_n248), .out0(new_n297));
  inv000aa1d42x5               g202(.a(new_n296), .o1(new_n298));
  and003aa1n02x5               g203(.a(new_n297), .b(new_n298), .c(new_n292), .o(new_n299));
  aoi022aa1n02x5               g204(.a(new_n295), .b(new_n296), .c(new_n286), .d(new_n299), .o1(\s[25] ));
  aoai13aa1n03x5               g205(.a(new_n296), .b(new_n293), .c(new_n207), .d(new_n285), .o1(new_n301));
  tech160nm_fixorc02aa1n02p5x5 g206(.a(\a[26] ), .b(\b[25] ), .out0(new_n302));
  nor042aa1n03x5               g207(.a(\b[24] ), .b(\a[25] ), .o1(new_n303));
  norp02aa1n02x5               g208(.a(new_n302), .b(new_n303), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n303), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n298), .c(new_n286), .d(new_n294), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[26] ));
  nand02aa1d04x5               g212(.a(new_n302), .b(new_n296), .o1(new_n308));
  nano23aa1n06x5               g213(.a(new_n308), .b(new_n284), .c(new_n263), .d(new_n223), .out0(new_n309));
  aoai13aa1n12x5               g214(.a(new_n309), .b(new_n216), .c(new_n129), .d(new_n198), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n308), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[26] ), .b(\b[25] ), .c(new_n305), .carry(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  aoi012aa1n12x5               g218(.a(new_n313), .b(new_n293), .c(new_n311), .o1(new_n314));
  nanp02aa1n02x5               g219(.a(new_n310), .b(new_n314), .o1(new_n315));
  xorc02aa1n12x5               g220(.a(\a[27] ), .b(\b[26] ), .out0(new_n316));
  aoi112aa1n02x5               g221(.a(new_n316), .b(new_n313), .c(new_n293), .d(new_n311), .o1(new_n317));
  aoi022aa1n02x5               g222(.a(new_n315), .b(new_n316), .c(new_n310), .d(new_n317), .o1(\s[27] ));
  aoai13aa1n04x5               g223(.a(new_n312), .b(new_n308), .c(new_n297), .d(new_n292), .o1(new_n319));
  aoai13aa1n02x5               g224(.a(new_n316), .b(new_n319), .c(new_n207), .d(new_n309), .o1(new_n320));
  tech160nm_fixorc02aa1n03p5x5 g225(.a(\a[28] ), .b(\b[27] ), .out0(new_n321));
  norp02aa1n02x5               g226(.a(\b[26] ), .b(\a[27] ), .o1(new_n322));
  norp02aa1n02x5               g227(.a(new_n321), .b(new_n322), .o1(new_n323));
  inv000aa1n03x5               g228(.a(new_n322), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n316), .o1(new_n325));
  aoai13aa1n03x5               g230(.a(new_n324), .b(new_n325), .c(new_n310), .d(new_n314), .o1(new_n326));
  aoi022aa1n03x5               g231(.a(new_n326), .b(new_n321), .c(new_n320), .d(new_n323), .o1(\s[28] ));
  and002aa1n02x5               g232(.a(new_n321), .b(new_n316), .o(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n319), .c(new_n207), .d(new_n309), .o1(new_n329));
  inv000aa1d42x5               g234(.a(new_n328), .o1(new_n330));
  oao003aa1n02x5               g235(.a(\a[28] ), .b(\b[27] ), .c(new_n324), .carry(new_n331));
  aoai13aa1n03x5               g236(.a(new_n331), .b(new_n330), .c(new_n310), .d(new_n314), .o1(new_n332));
  xorc02aa1n02x5               g237(.a(\a[29] ), .b(\b[28] ), .out0(new_n333));
  norb02aa1n02x5               g238(.a(new_n331), .b(new_n333), .out0(new_n334));
  aoi022aa1n03x5               g239(.a(new_n332), .b(new_n333), .c(new_n329), .d(new_n334), .o1(\s[29] ));
  xorb03aa1n02x5               g240(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g241(.a(new_n325), .b(new_n321), .c(new_n333), .out0(new_n337));
  aoai13aa1n02x5               g242(.a(new_n337), .b(new_n319), .c(new_n207), .d(new_n309), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n337), .o1(new_n339));
  oao003aa1n02x5               g244(.a(\a[29] ), .b(\b[28] ), .c(new_n331), .carry(new_n340));
  aoai13aa1n03x5               g245(.a(new_n340), .b(new_n339), .c(new_n310), .d(new_n314), .o1(new_n341));
  xorc02aa1n02x5               g246(.a(\a[30] ), .b(\b[29] ), .out0(new_n342));
  norb02aa1n02x5               g247(.a(new_n340), .b(new_n342), .out0(new_n343));
  aoi022aa1n03x5               g248(.a(new_n341), .b(new_n342), .c(new_n338), .d(new_n343), .o1(\s[30] ));
  nano32aa1n03x7               g249(.a(new_n325), .b(new_n342), .c(new_n321), .d(new_n333), .out0(new_n345));
  aoai13aa1n02x5               g250(.a(new_n345), .b(new_n319), .c(new_n207), .d(new_n309), .o1(new_n346));
  xorc02aa1n02x5               g251(.a(\a[31] ), .b(\b[30] ), .out0(new_n347));
  oao003aa1n02x5               g252(.a(\a[30] ), .b(\b[29] ), .c(new_n340), .carry(new_n348));
  norb02aa1n02x5               g253(.a(new_n348), .b(new_n347), .out0(new_n349));
  inv000aa1d42x5               g254(.a(new_n345), .o1(new_n350));
  aoai13aa1n03x5               g255(.a(new_n348), .b(new_n350), .c(new_n310), .d(new_n314), .o1(new_n351));
  aoi022aa1n03x5               g256(.a(new_n351), .b(new_n347), .c(new_n346), .d(new_n349), .o1(\s[31] ));
  aoi112aa1n02x5               g257(.a(new_n109), .b(new_n99), .c(new_n101), .d(new_n102), .o1(new_n353));
  aoi012aa1n02x5               g258(.a(new_n353), .b(new_n103), .c(new_n109), .o1(\s[3] ));
  aoi112aa1n02x5               g259(.a(new_n107), .b(new_n106), .c(new_n103), .d(new_n108), .o1(new_n355));
  aoib12aa1n02x5               g260(.a(new_n355), .b(new_n148), .c(new_n104), .out0(\s[4] ));
  norb02aa1n02x5               g261(.a(new_n115), .b(new_n114), .out0(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n357), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  norb02aa1n02x5               g263(.a(new_n113), .b(new_n112), .out0(new_n359));
  aoai13aa1n02x5               g264(.a(new_n359), .b(new_n114), .c(new_n148), .d(new_n115), .o1(new_n360));
  aoi112aa1n02x5               g265(.a(new_n114), .b(new_n359), .c(new_n148), .d(new_n115), .o1(new_n361));
  norb02aa1n02x5               g266(.a(new_n360), .b(new_n361), .out0(\s[6] ));
  inv000aa1d42x5               g267(.a(new_n112), .o1(new_n363));
  norb02aa1n02x5               g268(.a(new_n120), .b(new_n119), .out0(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n364), .b(new_n360), .c(new_n363), .out0(\s[7] ));
  aob012aa1n02x5               g270(.a(new_n364), .b(new_n360), .c(new_n363), .out0(new_n366));
  nanp02aa1n02x5               g271(.a(new_n366), .b(new_n126), .o1(new_n367));
  aoib12aa1n02x5               g272(.a(new_n119), .b(new_n118), .c(new_n117), .out0(new_n368));
  aoi022aa1n02x5               g273(.a(new_n367), .b(new_n123), .c(new_n366), .d(new_n368), .o1(\s[8] ));
  xnbna2aa1n03x5               g274(.a(new_n130), .b(new_n149), .c(new_n128), .out0(\s[9] ));
endmodule


