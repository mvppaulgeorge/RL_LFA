// Benchmark "adder" written by ABC on Wed Jul 17 23:40:29 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n315, new_n317, new_n318,
    new_n319, new_n320, new_n322, new_n324, new_n326, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv020aa1n10x5               g001(.a(\b[9] ), .o1(new_n97));
  nanb02aa1n12x5               g002(.a(\a[10] ), .b(new_n97), .out0(new_n98));
  nanp02aa1n09x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[8] ), .o1(new_n101));
  xnrc02aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .out0(new_n102));
  inv000aa1d42x5               g007(.a(\a[2] ), .o1(new_n103));
  inv000aa1d42x5               g008(.a(\b[1] ), .o1(new_n104));
  nanp02aa1n06x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  oao003aa1n02x5               g010(.a(new_n103), .b(new_n104), .c(new_n105), .carry(new_n106));
  nanb02aa1n02x5               g011(.a(new_n102), .b(new_n106), .out0(new_n107));
  inv000aa1d42x5               g012(.a(\a[3] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\a[4] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  aboi22aa1n03x5               g015(.a(\b[3] ), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n111));
  nor022aa1n06x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  aoi122aa1n06x5               g017(.a(new_n112), .b(\b[5] ), .c(\a[6] ), .d(\b[3] ), .e(\a[4] ), .o1(new_n113));
  xnrc02aa1n12x5               g018(.a(\b[7] ), .b(\a[8] ), .out0(new_n114));
  inv000aa1d42x5               g019(.a(new_n114), .o1(new_n115));
  nor022aa1n04x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  aoi012aa1n02x5               g021(.a(new_n116), .b(\a[5] ), .c(\b[4] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  norp02aa1n06x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nanb02aa1n06x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  norb02aa1n03x5               g025(.a(new_n117), .b(new_n120), .out0(new_n121));
  nanp03aa1n03x5               g026(.a(new_n121), .b(new_n115), .c(new_n113), .o1(new_n122));
  aoi022aa1n02x5               g027(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n123));
  oai012aa1n02x5               g028(.a(new_n123), .b(new_n116), .c(new_n112), .o1(new_n124));
  oab012aa1n02x4               g029(.a(new_n119), .b(\a[8] ), .c(\b[7] ), .out0(new_n125));
  aoi022aa1n06x5               g030(.a(new_n124), .b(new_n125), .c(\b[7] ), .d(\a[8] ), .o1(new_n126));
  inv000aa1n06x5               g031(.a(new_n126), .o1(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n122), .c(new_n107), .d(new_n111), .o1(new_n128));
  tech160nm_fioaoi03aa1n03p5x5 g033(.a(new_n100), .b(new_n101), .c(new_n128), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n98), .c(new_n99), .out0(\s[10] ));
  xorc02aa1n02x5               g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  nanp02aa1n06x5               g036(.a(new_n129), .b(new_n131), .o1(new_n132));
  nor002aa1n16x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  and002aa1n12x5               g038(.a(\b[10] ), .b(\a[11] ), .o(new_n134));
  norp02aa1n02x5               g039(.a(new_n134), .b(new_n133), .o1(new_n135));
  xobna2aa1n03x5               g040(.a(new_n135), .b(new_n132), .c(new_n99), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n133), .o1(new_n137));
  nanp03aa1n02x5               g042(.a(new_n132), .b(new_n99), .c(new_n135), .o1(new_n138));
  xorc02aa1n12x5               g043(.a(\a[12] ), .b(\b[11] ), .out0(new_n139));
  aobi12aa1n03x5               g044(.a(new_n139), .b(new_n138), .c(new_n137), .out0(new_n140));
  aoi113aa1n02x5               g045(.a(new_n139), .b(new_n133), .c(new_n132), .d(new_n135), .e(new_n99), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n140), .b(new_n141), .o1(\s[12] ));
  tech160nm_fioaoi03aa1n02p5x5 g047(.a(new_n103), .b(new_n104), .c(new_n105), .o1(new_n143));
  oai012aa1n06x5               g048(.a(new_n111), .b(new_n143), .c(new_n102), .o1(new_n144));
  nano23aa1n09x5               g049(.a(new_n120), .b(new_n114), .c(new_n113), .d(new_n117), .out0(new_n145));
  oai112aa1n06x5               g050(.a(new_n98), .b(new_n99), .c(\b[8] ), .d(\a[9] ), .o1(new_n146));
  aoi112aa1n09x5               g051(.a(new_n134), .b(new_n133), .c(\a[9] ), .d(\b[8] ), .o1(new_n147));
  nanb03aa1d24x5               g052(.a(new_n146), .b(new_n147), .c(new_n139), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n126), .c(new_n145), .d(new_n144), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  aoi022aa1n02x5               g056(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n152));
  oai022aa1n02x5               g057(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n153));
  aoai13aa1n04x5               g058(.a(new_n151), .b(new_n153), .c(new_n146), .d(new_n152), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(new_n150), .b(new_n154), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g061(.a(\a[14] ), .o1(new_n157));
  nor002aa1d32x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand42aa1n03x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  aoi012aa1n02x5               g064(.a(new_n158), .b(new_n155), .c(new_n159), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(new_n157), .out0(\s[14] ));
  inv000aa1d42x5               g066(.a(new_n158), .o1(new_n162));
  xnrc02aa1n12x5               g067(.a(\b[13] ), .b(\a[14] ), .out0(new_n163));
  nano22aa1d15x5               g068(.a(new_n163), .b(new_n162), .c(new_n159), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[13] ), .o1(new_n166));
  tech160nm_fioaoi03aa1n03p5x5 g071(.a(new_n157), .b(new_n166), .c(new_n158), .o1(new_n167));
  aoai13aa1n04x5               g072(.a(new_n167), .b(new_n165), .c(new_n150), .d(new_n154), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand02aa1n03x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nor042aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  nand42aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  aoi122aa1n02x5               g079(.a(new_n170), .b(new_n173), .c(new_n174), .d(new_n168), .e(new_n171), .o1(new_n175));
  aoi012aa1n02x5               g080(.a(new_n170), .b(new_n168), .c(new_n171), .o1(new_n176));
  nano22aa1n02x4               g081(.a(new_n176), .b(new_n173), .c(new_n174), .out0(new_n177));
  norp02aa1n02x5               g082(.a(new_n177), .b(new_n175), .o1(\s[16] ));
  nano23aa1n06x5               g083(.a(new_n170), .b(new_n172), .c(new_n174), .d(new_n171), .out0(new_n179));
  nano22aa1d15x5               g084(.a(new_n148), .b(new_n164), .c(new_n179), .out0(new_n180));
  aoai13aa1n06x5               g085(.a(new_n180), .b(new_n126), .c(new_n145), .d(new_n144), .o1(new_n181));
  nand42aa1n04x5               g086(.a(new_n164), .b(new_n179), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n170), .o1(new_n183));
  nanp02aa1n02x5               g088(.a(new_n174), .b(new_n171), .o1(new_n184));
  aoai13aa1n06x5               g089(.a(new_n173), .b(new_n184), .c(new_n167), .d(new_n183), .o1(new_n185));
  oab012aa1n12x5               g090(.a(new_n185), .b(new_n154), .c(new_n182), .out0(new_n186));
  nanp02aa1n09x5               g091(.a(new_n181), .b(new_n186), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[16] ), .o1(new_n191));
  oaoi03aa1n03x5               g096(.a(new_n190), .b(new_n191), .c(new_n187), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(new_n189), .out0(\s[18] ));
  xroi22aa1d06x4               g098(.a(new_n190), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n194));
  oai022aa1d24x5               g099(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n195));
  oaib12aa1n18x5               g100(.a(new_n195), .b(new_n189), .c(\b[17] ), .out0(new_n196));
  inv000aa1n12x5               g101(.a(new_n196), .o1(new_n197));
  nor042aa1n06x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand02aa1n08x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n201));
  aoi112aa1n02x5               g106(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n202));
  norb02aa1n02x7               g107(.a(new_n201), .b(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand02aa1d16x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  nona22aa1n02x5               g112(.a(new_n201), .b(new_n207), .c(new_n198), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n207), .o1(new_n209));
  oaoi13aa1n06x5               g114(.a(new_n209), .b(new_n201), .c(\a[19] ), .d(\b[18] ), .o1(new_n210));
  norb02aa1n03x4               g115(.a(new_n208), .b(new_n210), .out0(\s[20] ));
  nano23aa1n09x5               g116(.a(new_n198), .b(new_n205), .c(new_n206), .d(new_n199), .out0(new_n212));
  nanp02aa1n02x5               g117(.a(new_n194), .b(new_n212), .o1(new_n213));
  nona23aa1n09x5               g118(.a(new_n206), .b(new_n199), .c(new_n198), .d(new_n205), .out0(new_n214));
  aoi012aa1n09x5               g119(.a(new_n205), .b(new_n198), .c(new_n206), .o1(new_n215));
  oai012aa1n18x5               g120(.a(new_n215), .b(new_n214), .c(new_n196), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n04x5               g122(.a(new_n217), .b(new_n213), .c(new_n181), .d(new_n186), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  xorc02aa1n02x5               g125(.a(\a[21] ), .b(\b[20] ), .out0(new_n221));
  xorc02aa1n02x5               g126(.a(\a[22] ), .b(\b[21] ), .out0(new_n222));
  aoi112aa1n02x5               g127(.a(new_n220), .b(new_n222), .c(new_n218), .d(new_n221), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n222), .b(new_n220), .c(new_n218), .d(new_n221), .o1(new_n224));
  norb02aa1n02x7               g129(.a(new_n224), .b(new_n223), .out0(\s[22] ));
  inv000aa1d42x5               g130(.a(\a[21] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  nanp03aa1n02x5               g133(.a(new_n228), .b(new_n194), .c(new_n212), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\b[21] ), .o1(new_n230));
  oaoi03aa1n09x5               g135(.a(new_n227), .b(new_n230), .c(new_n220), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n216), .c(new_n228), .o1(new_n233));
  aoai13aa1n04x5               g138(.a(new_n233), .b(new_n229), .c(new_n181), .d(new_n186), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  tech160nm_fixorc02aa1n05x5   g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  tech160nm_fixorc02aa1n05x5   g142(.a(\a[24] ), .b(\b[23] ), .out0(new_n238));
  aoi112aa1n02x5               g143(.a(new_n236), .b(new_n238), .c(new_n234), .d(new_n237), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n238), .b(new_n236), .c(new_n234), .d(new_n237), .o1(new_n240));
  norb02aa1n02x7               g145(.a(new_n240), .b(new_n239), .out0(\s[24] ));
  oabi12aa1n03x5               g146(.a(new_n185), .b(new_n154), .c(new_n182), .out0(new_n242));
  and002aa1n02x5               g147(.a(new_n238), .b(new_n237), .o(new_n243));
  inv030aa1n02x5               g148(.a(new_n243), .o1(new_n244));
  nano32aa1n02x4               g149(.a(new_n244), .b(new_n228), .c(new_n194), .d(new_n212), .out0(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n242), .c(new_n128), .d(new_n180), .o1(new_n246));
  inv020aa1n03x5               g151(.a(new_n215), .o1(new_n247));
  aoai13aa1n06x5               g152(.a(new_n228), .b(new_n247), .c(new_n212), .d(new_n197), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n249));
  oab012aa1n04x5               g154(.a(new_n249), .b(\a[24] ), .c(\b[23] ), .out0(new_n250));
  aoai13aa1n12x5               g155(.a(new_n250), .b(new_n244), .c(new_n248), .d(new_n231), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  xnrc02aa1n12x5               g157(.a(\b[24] ), .b(\a[25] ), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n246), .c(new_n252), .out0(\s[25] ));
  nor042aa1n03x5               g160(.a(\b[24] ), .b(\a[25] ), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n254), .b(new_n251), .c(new_n187), .d(new_n245), .o1(new_n258));
  xnrc02aa1n06x5               g163(.a(\b[25] ), .b(\a[26] ), .out0(new_n259));
  nand43aa1n03x5               g164(.a(new_n258), .b(new_n257), .c(new_n259), .o1(new_n260));
  tech160nm_fiaoi012aa1n03p5x5 g165(.a(new_n259), .b(new_n258), .c(new_n257), .o1(new_n261));
  norb02aa1n03x4               g166(.a(new_n260), .b(new_n261), .out0(\s[26] ));
  nor042aa1n06x5               g167(.a(new_n259), .b(new_n253), .o1(new_n263));
  nano22aa1n03x7               g168(.a(new_n229), .b(new_n243), .c(new_n263), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n242), .c(new_n128), .d(new_n180), .o1(new_n265));
  nand02aa1d08x5               g170(.a(new_n251), .b(new_n263), .o1(new_n266));
  oao003aa1n02x5               g171(.a(\a[26] ), .b(\b[25] ), .c(new_n257), .carry(new_n267));
  nor042aa1n03x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(\b[26] ), .b(\a[27] ), .o1(new_n269));
  norb02aa1n09x5               g174(.a(new_n269), .b(new_n268), .out0(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoi013aa1n06x4               g176(.a(new_n271), .b(new_n265), .c(new_n266), .d(new_n267), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n243), .b(new_n232), .c(new_n216), .d(new_n228), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n263), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n267), .b(new_n274), .c(new_n273), .d(new_n250), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(new_n275), .b(new_n270), .c(new_n187), .d(new_n264), .o1(new_n276));
  norp02aa1n02x5               g181(.a(new_n272), .b(new_n276), .o1(\s[27] ));
  inv000aa1n06x5               g182(.a(new_n268), .o1(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[27] ), .b(\a[28] ), .out0(new_n279));
  nano22aa1n03x5               g184(.a(new_n272), .b(new_n278), .c(new_n279), .out0(new_n280));
  aobi12aa1n06x5               g185(.a(new_n264), .b(new_n181), .c(new_n186), .out0(new_n281));
  oaih12aa1n02x5               g186(.a(new_n270), .b(new_n275), .c(new_n281), .o1(new_n282));
  aoi012aa1n02x7               g187(.a(new_n279), .b(new_n282), .c(new_n278), .o1(new_n283));
  norp02aa1n03x5               g188(.a(new_n283), .b(new_n280), .o1(\s[28] ));
  nano22aa1n12x5               g189(.a(new_n279), .b(new_n278), .c(new_n269), .out0(new_n285));
  oaih12aa1n02x5               g190(.a(new_n285), .b(new_n275), .c(new_n281), .o1(new_n286));
  oao003aa1n03x5               g191(.a(\a[28] ), .b(\b[27] ), .c(new_n278), .carry(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  tech160nm_fiaoi012aa1n02p5x5 g193(.a(new_n288), .b(new_n286), .c(new_n287), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n285), .o1(new_n290));
  aoi013aa1n06x4               g195(.a(new_n290), .b(new_n265), .c(new_n266), .d(new_n267), .o1(new_n291));
  nano22aa1n03x5               g196(.a(new_n291), .b(new_n287), .c(new_n288), .out0(new_n292));
  norp02aa1n03x5               g197(.a(new_n289), .b(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g199(.a(new_n288), .b(new_n279), .c(new_n269), .d(new_n278), .out0(new_n295));
  oaih12aa1n02x5               g200(.a(new_n295), .b(new_n275), .c(new_n281), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[29] ), .b(\b[28] ), .c(new_n287), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[29] ), .b(\a[30] ), .out0(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n298), .b(new_n296), .c(new_n297), .o1(new_n299));
  inv000aa1n02x5               g204(.a(new_n295), .o1(new_n300));
  aoi013aa1n02x5               g205(.a(new_n300), .b(new_n265), .c(new_n266), .d(new_n267), .o1(new_n301));
  nano22aa1n03x5               g206(.a(new_n301), .b(new_n297), .c(new_n298), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n299), .b(new_n302), .o1(\s[30] ));
  norb03aa1n02x5               g208(.a(new_n285), .b(new_n298), .c(new_n288), .out0(new_n304));
  inv000aa1n02x5               g209(.a(new_n304), .o1(new_n305));
  aoi013aa1n02x5               g210(.a(new_n305), .b(new_n265), .c(new_n266), .d(new_n267), .o1(new_n306));
  oao003aa1n03x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n297), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  nano22aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n308), .out0(new_n309));
  oaih12aa1n02x5               g214(.a(new_n304), .b(new_n275), .c(new_n281), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n308), .b(new_n310), .c(new_n307), .o1(new_n311));
  norp02aa1n03x5               g216(.a(new_n311), .b(new_n309), .o1(\s[31] ));
  xorb03aa1n02x5               g217(.a(new_n143), .b(\b[2] ), .c(new_n108), .out0(\s[3] ));
  xorc02aa1n02x5               g218(.a(\a[4] ), .b(\b[3] ), .out0(new_n314));
  aoi012aa1n02x5               g219(.a(new_n314), .b(new_n108), .c(new_n110), .o1(new_n315));
  aoi022aa1n02x5               g220(.a(new_n144), .b(new_n314), .c(new_n107), .d(new_n315), .o1(\s[4] ));
  inv000aa1d42x5               g221(.a(\b[3] ), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[5] ), .b(\b[4] ), .out0(new_n318));
  oaoi13aa1n02x5               g223(.a(new_n318), .b(new_n144), .c(new_n109), .d(new_n317), .o1(new_n319));
  oai112aa1n02x5               g224(.a(new_n144), .b(new_n318), .c(new_n317), .d(new_n109), .o1(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(\s[5] ));
  norb02aa1n06x5               g226(.a(new_n320), .b(new_n112), .out0(new_n322));
  xnrb03aa1n02x5               g227(.a(new_n322), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fioaoi03aa1n03p5x5 g228(.a(\a[6] ), .b(\b[5] ), .c(new_n322), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoai13aa1n04x5               g230(.a(new_n115), .b(new_n119), .c(new_n324), .d(new_n118), .o1(new_n326));
  aoi112aa1n02x5               g231(.a(new_n119), .b(new_n115), .c(new_n324), .d(new_n118), .o1(new_n327));
  norb02aa1n02x5               g232(.a(new_n326), .b(new_n327), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


