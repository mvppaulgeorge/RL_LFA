// Benchmark "adder" written by ABC on Wed Jul 17 22:14:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n309, new_n312,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n320;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_finand02aa1n03p5x5 g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand22aa1n12x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  oai012aa1n09x5               g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  tech160nm_fixnrc02aa1n04x5   g005(.a(\b[3] ), .b(\a[4] ), .out0(new_n101));
  nor022aa1n08x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanb02aa1n09x5               g008(.a(new_n102), .b(new_n103), .out0(new_n104));
  inv000aa1d42x5               g009(.a(\a[3] ), .o1(new_n105));
  nanb02aa1n12x5               g010(.a(\b[2] ), .b(new_n105), .out0(new_n106));
  oao003aa1n03x5               g011(.a(\a[4] ), .b(\b[3] ), .c(new_n106), .carry(new_n107));
  oai013aa1d12x5               g012(.a(new_n107), .b(new_n101), .c(new_n100), .d(new_n104), .o1(new_n108));
  nor022aa1n08x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand22aa1n04x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nor002aa1d32x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand02aa1n16x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nona23aa1d18x5               g017(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[5] ), .b(\a[6] ), .out0(new_n114));
  nor042aa1n04x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  nor043aa1n06x5               g022(.a(new_n113), .b(new_n114), .c(new_n117), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[6] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[5] ), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(new_n119), .b(new_n120), .c(new_n115), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n111), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  oabi12aa1n06x5               g028(.a(new_n123), .b(new_n113), .c(new_n121), .out0(new_n124));
  aoi012aa1n02x5               g029(.a(new_n124), .b(new_n108), .c(new_n118), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[9] ), .b(\b[8] ), .c(new_n125), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n04x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nor042aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanp02aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  aoi012aa1n12x5               g035(.a(new_n129), .b(new_n128), .c(new_n130), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  nano23aa1n06x5               g037(.a(new_n128), .b(new_n129), .c(new_n130), .d(new_n132), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n124), .c(new_n108), .d(new_n118), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(new_n134), .b(new_n131), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(\a[12] ), .o1(new_n137));
  nor002aa1d32x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand42aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  aoi012aa1n02x5               g044(.a(new_n138), .b(new_n135), .c(new_n139), .o1(new_n140));
  xorb03aa1n02x5               g045(.a(new_n140), .b(\b[11] ), .c(new_n137), .out0(\s[12] ));
  nor002aa1d32x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand22aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nona23aa1d18x5               g048(.a(new_n143), .b(new_n139), .c(new_n138), .d(new_n142), .out0(new_n144));
  ao0012aa1n03x7               g049(.a(new_n142), .b(new_n138), .c(new_n143), .o(new_n145));
  oabi12aa1n18x5               g050(.a(new_n145), .b(new_n144), .c(new_n131), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n133), .b(new_n144), .out0(new_n148));
  aoai13aa1n06x5               g053(.a(new_n148), .b(new_n124), .c(new_n108), .d(new_n118), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n149), .b(new_n147), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g056(.a(\a[14] ), .o1(new_n152));
  nor002aa1n03x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1d28x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n03x5               g059(.a(new_n153), .b(new_n150), .c(new_n154), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(new_n152), .out0(\s[14] ));
  nor022aa1n08x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand42aa1n08x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nona23aa1n02x4               g063(.a(new_n158), .b(new_n154), .c(new_n153), .d(new_n157), .out0(new_n159));
  nano23aa1n03x7               g064(.a(new_n153), .b(new_n157), .c(new_n158), .d(new_n154), .out0(new_n160));
  aoi012aa1n02x5               g065(.a(new_n157), .b(new_n153), .c(new_n158), .o1(new_n161));
  aobi12aa1n02x5               g066(.a(new_n161), .b(new_n146), .c(new_n160), .out0(new_n162));
  tech160nm_fioai012aa1n04x5   g067(.a(new_n162), .b(new_n149), .c(new_n159), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand42aa1n20x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nor042aa1n02x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nand42aa1n08x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  nanb02aa1n02x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n165), .b(new_n169), .c(new_n163), .d(new_n166), .o1(new_n171));
  nanb02aa1n03x5               g076(.a(new_n171), .b(new_n170), .out0(\s[16] ));
  nano23aa1n03x7               g077(.a(new_n138), .b(new_n142), .c(new_n143), .d(new_n139), .out0(new_n173));
  nano23aa1n03x7               g078(.a(new_n165), .b(new_n167), .c(new_n168), .d(new_n166), .out0(new_n174));
  nand22aa1n03x5               g079(.a(new_n174), .b(new_n160), .o1(new_n175));
  nano22aa1n03x7               g080(.a(new_n175), .b(new_n133), .c(new_n173), .out0(new_n176));
  aoai13aa1n12x5               g081(.a(new_n176), .b(new_n124), .c(new_n108), .d(new_n118), .o1(new_n177));
  aoi012aa1n02x5               g082(.a(new_n167), .b(new_n165), .c(new_n168), .o1(new_n178));
  oaib12aa1n02x5               g083(.a(new_n178), .b(new_n161), .c(new_n174), .out0(new_n179));
  aoib12aa1n12x5               g084(.a(new_n179), .b(new_n146), .c(new_n175), .out0(new_n180));
  xorc02aa1n12x5               g085(.a(\a[17] ), .b(\b[16] ), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n177), .c(new_n180), .out0(\s[17] ));
  nanp02aa1n06x5               g087(.a(new_n177), .b(new_n180), .o1(new_n183));
  nor042aa1n04x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  aoi012aa1n06x5               g089(.a(new_n184), .b(new_n183), .c(new_n181), .o1(new_n185));
  inv040aa1d32x5               g090(.a(\a[18] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[17] ), .o1(new_n187));
  nanp02aa1n04x5               g092(.a(new_n187), .b(new_n186), .o1(new_n188));
  nand22aa1n04x5               g093(.a(\b[17] ), .b(\a[18] ), .o1(new_n189));
  xnbna2aa1n03x5               g094(.a(new_n185), .b(new_n189), .c(new_n188), .out0(\s[18] ));
  oaoi03aa1n02x5               g095(.a(new_n186), .b(new_n187), .c(new_n184), .o1(new_n191));
  inv000aa1n06x5               g096(.a(new_n181), .o1(new_n192));
  nano22aa1n12x5               g097(.a(new_n192), .b(new_n188), .c(new_n189), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n191), .b(new_n194), .c(new_n177), .d(new_n180), .o1(new_n195));
  xorb03aa1n03x5               g100(.a(new_n195), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand42aa1n04x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nor042aa1d18x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nand42aa1d28x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  norb02aa1n12x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n198), .c(new_n195), .d(new_n199), .o1(new_n204));
  norb02aa1n06x4               g109(.a(new_n199), .b(new_n198), .out0(new_n205));
  nand22aa1n03x5               g110(.a(new_n195), .b(new_n205), .o1(new_n206));
  nona22aa1n03x5               g111(.a(new_n206), .b(new_n203), .c(new_n198), .out0(new_n207));
  nanp02aa1n03x5               g112(.a(new_n207), .b(new_n204), .o1(\s[20] ));
  aob012aa1n03x5               g113(.a(new_n188), .b(new_n184), .c(new_n189), .out0(new_n209));
  nano23aa1n06x5               g114(.a(new_n198), .b(new_n200), .c(new_n201), .d(new_n199), .out0(new_n210));
  aoi012aa1d18x5               g115(.a(new_n200), .b(new_n198), .c(new_n201), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoi012aa1n02x5               g117(.a(new_n212), .b(new_n210), .c(new_n209), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(new_n193), .b(new_n210), .o1(new_n214));
  aoai13aa1n06x5               g119(.a(new_n213), .b(new_n214), .c(new_n177), .d(new_n180), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  nand42aa1d28x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  nor022aa1n16x5               g124(.a(\b[21] ), .b(\a[22] ), .o1(new_n220));
  nand02aa1d28x5               g125(.a(\b[21] ), .b(\a[22] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n217), .c(new_n215), .d(new_n219), .o1(new_n224));
  nand02aa1n03x5               g129(.a(new_n215), .b(new_n219), .o1(new_n225));
  nona22aa1n02x5               g130(.a(new_n225), .b(new_n223), .c(new_n217), .out0(new_n226));
  nanp02aa1n03x5               g131(.a(new_n226), .b(new_n224), .o1(\s[22] ));
  nano23aa1d15x5               g132(.a(new_n217), .b(new_n220), .c(new_n221), .d(new_n218), .out0(new_n228));
  nanp03aa1n02x5               g133(.a(new_n193), .b(new_n210), .c(new_n228), .o1(new_n229));
  nano22aa1n02x4               g134(.a(new_n191), .b(new_n205), .c(new_n202), .out0(new_n230));
  ao0012aa1n03x7               g135(.a(new_n220), .b(new_n217), .c(new_n221), .o(new_n231));
  oaoi13aa1n02x5               g136(.a(new_n231), .b(new_n228), .c(new_n230), .d(new_n212), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n229), .c(new_n177), .d(new_n180), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n09x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  nand02aa1d24x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  nor042aa1n06x5               g142(.a(\b[23] ), .b(\a[24] ), .o1(new_n238));
  nand02aa1d24x5               g143(.a(\b[23] ), .b(\a[24] ), .o1(new_n239));
  nanb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n235), .c(new_n233), .d(new_n237), .o1(new_n241));
  nand22aa1n03x5               g146(.a(new_n233), .b(new_n237), .o1(new_n242));
  nona22aa1n03x5               g147(.a(new_n242), .b(new_n240), .c(new_n235), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n243), .b(new_n241), .o1(\s[24] ));
  nand03aa1n04x5               g149(.a(new_n209), .b(new_n205), .c(new_n202), .o1(new_n245));
  nano23aa1d15x5               g150(.a(new_n235), .b(new_n238), .c(new_n239), .d(new_n236), .out0(new_n246));
  nand22aa1n09x5               g151(.a(new_n246), .b(new_n228), .o1(new_n247));
  tech160nm_fiao0012aa1n02p5x5 g152(.a(new_n238), .b(new_n235), .c(new_n239), .o(new_n248));
  aoi012aa1n12x5               g153(.a(new_n248), .b(new_n246), .c(new_n231), .o1(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n247), .c(new_n245), .d(new_n211), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  nanb03aa1n02x5               g156(.a(new_n247), .b(new_n193), .c(new_n210), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n251), .b(new_n252), .c(new_n177), .d(new_n180), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g159(.a(\b[24] ), .b(\a[25] ), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[25] ), .b(\b[24] ), .out0(new_n256));
  xnrc02aa1n02x5               g161(.a(\b[25] ), .b(\a[26] ), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n255), .c(new_n253), .d(new_n256), .o1(new_n258));
  nand02aa1n04x5               g163(.a(new_n253), .b(new_n256), .o1(new_n259));
  nona22aa1n02x5               g164(.a(new_n259), .b(new_n257), .c(new_n255), .out0(new_n260));
  nanp02aa1n03x5               g165(.a(new_n260), .b(new_n258), .o1(\s[26] ));
  inv000aa1d42x5               g166(.a(new_n247), .o1(new_n262));
  norb02aa1n02x7               g167(.a(new_n256), .b(new_n257), .out0(new_n263));
  nanb03aa1n03x5               g168(.a(new_n214), .b(new_n263), .c(new_n262), .out0(new_n264));
  inv000aa1d42x5               g169(.a(\a[26] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(\b[25] ), .o1(new_n266));
  oaoi03aa1n02x5               g171(.a(new_n265), .b(new_n266), .c(new_n255), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  tech160nm_fiaoi012aa1n05x5   g173(.a(new_n268), .b(new_n250), .c(new_n263), .o1(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n264), .c(new_n177), .d(new_n180), .o1(new_n270));
  xorb03aa1n03x5               g175(.a(new_n270), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[27] ), .b(\b[26] ), .out0(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[27] ), .b(\a[28] ), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n275));
  nano22aa1n03x7               g180(.a(new_n214), .b(new_n262), .c(new_n263), .out0(new_n276));
  nanp02aa1n06x5               g181(.a(new_n250), .b(new_n263), .o1(new_n277));
  nanp02aa1n06x5               g182(.a(new_n277), .b(new_n267), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n273), .b(new_n278), .c(new_n183), .d(new_n276), .o1(new_n279));
  nona22aa1n02x4               g184(.a(new_n279), .b(new_n274), .c(new_n272), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n275), .b(new_n280), .o1(\s[28] ));
  inv000aa1d42x5               g186(.a(\a[28] ), .o1(new_n282));
  inv000aa1d42x5               g187(.a(\b[27] ), .o1(new_n283));
  oaoi03aa1n09x5               g188(.a(new_n282), .b(new_n283), .c(new_n272), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  norb02aa1n02x5               g190(.a(new_n273), .b(new_n274), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n278), .c(new_n183), .d(new_n276), .o1(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  nona22aa1n03x5               g193(.a(new_n287), .b(new_n288), .c(new_n285), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n288), .b(new_n285), .c(new_n270), .d(new_n286), .o1(new_n290));
  nanp02aa1n03x5               g195(.a(new_n290), .b(new_n289), .o1(\s[29] ));
  xorb03aa1n02x5               g196(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  tech160nm_fioaoi03aa1n03p5x5 g197(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .o1(new_n293));
  norb03aa1n02x5               g198(.a(new_n273), .b(new_n288), .c(new_n274), .out0(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n293), .c(new_n270), .d(new_n294), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n294), .b(new_n278), .c(new_n183), .d(new_n276), .o1(new_n297));
  nona22aa1n02x4               g202(.a(new_n297), .b(new_n295), .c(new_n293), .out0(new_n298));
  nanp02aa1n03x5               g203(.a(new_n296), .b(new_n298), .o1(\s[30] ));
  norb02aa1n02x5               g204(.a(new_n294), .b(new_n295), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n278), .c(new_n183), .d(new_n276), .o1(new_n301));
  nanb02aa1n02x5               g206(.a(new_n295), .b(new_n293), .out0(new_n302));
  oai012aa1n02x5               g207(.a(new_n302), .b(\b[29] ), .c(\a[30] ), .o1(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  nona22aa1n03x5               g209(.a(new_n301), .b(new_n303), .c(new_n304), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n304), .b(new_n303), .c(new_n270), .d(new_n300), .o1(new_n306));
  nanp02aa1n03x5               g211(.a(new_n306), .b(new_n305), .o1(\s[31] ));
  xnbna2aa1n03x5               g212(.a(new_n100), .b(new_n103), .c(new_n106), .out0(\s[3] ));
  oaoi03aa1n02x5               g213(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n309));
  xorb03aa1n02x5               g214(.a(new_n309), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g215(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g216(.a(new_n116), .b(new_n108), .c(new_n115), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[5] ), .c(new_n119), .out0(\s[6] ));
  inv000aa1d42x5               g218(.a(new_n112), .o1(new_n314));
  and002aa1n02x5               g219(.a(\b[5] ), .b(\a[6] ), .o(new_n315));
  nanb02aa1n02x5               g220(.a(new_n114), .b(new_n312), .out0(new_n316));
  nona32aa1n02x4               g221(.a(new_n316), .b(new_n315), .c(new_n314), .d(new_n111), .out0(new_n317));
  aboi22aa1n03x5               g222(.a(new_n315), .b(new_n316), .c(new_n122), .d(new_n112), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n317), .b(new_n318), .out0(\s[7] ));
  norb02aa1n02x5               g224(.a(new_n110), .b(new_n109), .out0(new_n320));
  xnbna2aa1n03x5               g225(.a(new_n320), .b(new_n317), .c(new_n122), .out0(\s[8] ));
  xnrb03aa1n02x5               g226(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


