// Benchmark "adder" written by ABC on Thu Jul 18 02:44:56 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n325, new_n326,
    new_n328, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  nanp02aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n09x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nor002aa1n03x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oai012aa1n06x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  nor022aa1n16x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand22aa1n09x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n09x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .d(new_n102), .out0(new_n106));
  tech160nm_fiaoi012aa1n03p5x5 g011(.a(new_n105), .b(new_n102), .c(new_n104), .o1(new_n107));
  oai012aa1n12x5               g012(.a(new_n107), .b(new_n106), .c(new_n101), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\a[6] ), .o1(new_n110));
  inv040aa1d28x5               g015(.a(\b[5] ), .o1(new_n111));
  nor022aa1n12x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  aoi012aa1n02x5               g017(.a(new_n112), .b(new_n110), .c(new_n111), .o1(new_n113));
  norp02aa1n24x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand22aa1n09x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand22aa1n12x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  norp02aa1n24x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nona23aa1n09x5               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nand42aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano32aa1n03x7               g024(.a(new_n118), .b(new_n113), .c(new_n109), .d(new_n119), .out0(new_n120));
  tech160nm_fioaoi03aa1n02p5x5 g025(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n121));
  ao0012aa1n03x7               g026(.a(new_n117), .b(new_n114), .c(new_n116), .o(new_n122));
  oabi12aa1n06x5               g027(.a(new_n122), .b(new_n118), .c(new_n121), .out0(new_n123));
  nor042aa1d18x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nand42aa1n16x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n127));
  nor042aa1d18x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n06x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n97), .out0(\s[10] ));
  nor042aa1d18x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand02aa1d12x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanb02aa1n02x5               g038(.a(new_n132), .b(new_n133), .out0(new_n134));
  nona22aa1n02x4               g039(.a(new_n127), .b(new_n128), .c(new_n124), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n134), .b(new_n135), .c(new_n129), .out0(\s[11] ));
  aoi013aa1n02x4               g041(.a(new_n132), .b(new_n135), .c(new_n133), .d(new_n129), .o1(new_n137));
  xnrb03aa1n03x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norb03aa1n03x5               g043(.a(new_n125), .b(new_n124), .c(new_n132), .out0(new_n139));
  nor002aa1d24x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand02aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nano22aa1n03x7               g046(.a(new_n140), .b(new_n133), .c(new_n141), .out0(new_n142));
  nand03aa1n04x5               g047(.a(new_n142), .b(new_n139), .c(new_n130), .o1(new_n143));
  inv000aa1n02x5               g048(.a(new_n143), .o1(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n145));
  nanb03aa1n12x5               g050(.a(new_n140), .b(new_n141), .c(new_n133), .out0(new_n146));
  inv040aa1n09x5               g051(.a(new_n132), .o1(new_n147));
  oai112aa1n06x5               g052(.a(new_n147), .b(new_n129), .c(new_n128), .d(new_n124), .o1(new_n148));
  aoi012aa1d18x5               g053(.a(new_n140), .b(new_n132), .c(new_n141), .o1(new_n149));
  oai012aa1n18x5               g054(.a(new_n149), .b(new_n148), .c(new_n146), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  nor042aa1d18x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1d28x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  xnbna2aa1n03x5               g059(.a(new_n154), .b(new_n145), .c(new_n151), .out0(\s[13] ));
  inv000aa1d42x5               g060(.a(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(\b[12] ), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(new_n145), .b(new_n151), .o1(new_n158));
  oaoi03aa1n02x5               g063(.a(new_n156), .b(new_n157), .c(new_n158), .o1(new_n159));
  xnrb03aa1n02x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1d18x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand42aa1d28x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nano23aa1d15x5               g067(.a(new_n152), .b(new_n161), .c(new_n162), .d(new_n153), .out0(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  oa0012aa1n02x5               g069(.a(new_n162), .b(new_n161), .c(new_n152), .o(new_n165));
  inv040aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  aoai13aa1n04x5               g071(.a(new_n166), .b(new_n164), .c(new_n145), .d(new_n151), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n09x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand02aa1d24x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nor042aa1n09x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nand02aa1d28x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n169), .c(new_n167), .d(new_n170), .o1(new_n174));
  aoi112aa1n02x5               g079(.a(new_n169), .b(new_n173), .c(new_n167), .d(new_n170), .o1(new_n175));
  norb02aa1n03x4               g080(.a(new_n174), .b(new_n175), .out0(\s[16] ));
  nano23aa1d15x5               g081(.a(new_n169), .b(new_n171), .c(new_n172), .d(new_n170), .out0(new_n177));
  nano22aa1d15x5               g082(.a(new_n143), .b(new_n163), .c(new_n177), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n179));
  aoai13aa1n06x5               g084(.a(new_n177), .b(new_n165), .c(new_n150), .d(new_n163), .o1(new_n180));
  aoi012aa1d18x5               g085(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n181));
  nand23aa1n06x5               g086(.a(new_n179), .b(new_n180), .c(new_n181), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g088(.a(\a[18] ), .o1(new_n184));
  inv030aa1d32x5               g089(.a(\a[17] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\b[16] ), .o1(new_n186));
  oaoi03aa1n03x5               g091(.a(new_n185), .b(new_n186), .c(new_n182), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[17] ), .c(new_n184), .out0(\s[18] ));
  inv040aa1n09x5               g093(.a(new_n123), .o1(new_n189));
  aob012aa1d18x5               g094(.a(new_n189), .b(new_n108), .c(new_n120), .out0(new_n190));
  inv000aa1d42x5               g095(.a(new_n177), .o1(new_n191));
  oai012aa1n03x5               g096(.a(new_n129), .b(\b[10] ), .c(\a[11] ), .o1(new_n192));
  oab012aa1n03x5               g097(.a(new_n192), .b(new_n124), .c(new_n128), .out0(new_n193));
  inv020aa1n02x5               g098(.a(new_n149), .o1(new_n194));
  aoai13aa1n04x5               g099(.a(new_n163), .b(new_n194), .c(new_n193), .d(new_n142), .o1(new_n195));
  aoai13aa1n12x5               g100(.a(new_n181), .b(new_n191), .c(new_n195), .d(new_n166), .o1(new_n196));
  xroi22aa1d06x4               g101(.a(new_n185), .b(\b[16] ), .c(new_n184), .d(\b[17] ), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n196), .c(new_n190), .d(new_n178), .o1(new_n198));
  inv000aa1d42x5               g103(.a(\b[17] ), .o1(new_n199));
  oai022aa1d18x5               g104(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n200));
  oa0012aa1n02x5               g105(.a(new_n200), .b(new_n199), .c(new_n184), .o(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  xnrc02aa1n12x5               g107(.a(\b[18] ), .b(\a[19] ), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n198), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g111(.a(\a[19] ), .o1(new_n207));
  inv040aa1d32x5               g112(.a(\b[18] ), .o1(new_n208));
  nand42aa1n02x5               g113(.a(new_n208), .b(new_n207), .o1(new_n209));
  aoai13aa1n03x5               g114(.a(new_n204), .b(new_n201), .c(new_n182), .d(new_n197), .o1(new_n210));
  tech160nm_fixnrc02aa1n04x5   g115(.a(\b[19] ), .b(\a[20] ), .out0(new_n211));
  tech160nm_fiaoi012aa1n02p5x5 g116(.a(new_n211), .b(new_n210), .c(new_n209), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n203), .b(new_n198), .c(new_n202), .o1(new_n213));
  nano22aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n211), .out0(new_n214));
  norp02aa1n03x5               g119(.a(new_n212), .b(new_n214), .o1(\s[20] ));
  nona22aa1d18x5               g120(.a(new_n197), .b(new_n203), .c(new_n211), .out0(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n196), .c(new_n190), .d(new_n178), .o1(new_n218));
  inv000aa1d42x5               g123(.a(\b[19] ), .o1(new_n219));
  oai122aa1n12x5               g124(.a(new_n200), .b(new_n207), .c(new_n208), .d(new_n184), .e(new_n199), .o1(new_n220));
  oai112aa1n06x5               g125(.a(new_n220), .b(new_n209), .c(\b[19] ), .d(\a[20] ), .o1(new_n221));
  oaib12aa1n12x5               g126(.a(new_n221), .b(new_n219), .c(\a[20] ), .out0(new_n222));
  xorc02aa1n12x5               g127(.a(\a[21] ), .b(\b[20] ), .out0(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n218), .c(new_n222), .out0(\s[21] ));
  orn002aa1n03x5               g129(.a(\a[21] ), .b(\b[20] ), .o(new_n225));
  inv000aa1d42x5               g130(.a(new_n222), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n223), .b(new_n226), .c(new_n182), .d(new_n217), .o1(new_n227));
  xorc02aa1n12x5               g132(.a(\a[22] ), .b(\b[21] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  tech160nm_fiaoi012aa1n02p5x5 g134(.a(new_n229), .b(new_n227), .c(new_n225), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n223), .o1(new_n231));
  tech160nm_fiaoi012aa1n03p5x5 g136(.a(new_n231), .b(new_n218), .c(new_n222), .o1(new_n232));
  nano22aa1n03x5               g137(.a(new_n232), .b(new_n225), .c(new_n229), .out0(new_n233));
  nor002aa1n02x5               g138(.a(new_n230), .b(new_n233), .o1(\s[22] ));
  xnrc02aa1n12x5               g139(.a(\b[22] ), .b(\a[23] ), .out0(new_n235));
  nand02aa1d08x5               g140(.a(new_n228), .b(new_n223), .o1(new_n236));
  nor042aa1n03x5               g141(.a(new_n216), .b(new_n236), .o1(new_n237));
  oaoi03aa1n03x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .o1(new_n238));
  oabi12aa1n06x5               g143(.a(new_n238), .b(new_n222), .c(new_n236), .out0(new_n239));
  aoai13aa1n02x5               g144(.a(new_n235), .b(new_n239), .c(new_n182), .d(new_n237), .o1(new_n240));
  norp02aa1n02x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  and002aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o(new_n242));
  aoai13aa1n06x5               g147(.a(new_n237), .b(new_n196), .c(new_n190), .d(new_n178), .o1(new_n243));
  nona32aa1n02x5               g148(.a(new_n243), .b(new_n239), .c(new_n242), .d(new_n241), .out0(new_n244));
  nanp02aa1n02x5               g149(.a(new_n240), .b(new_n244), .o1(\s[23] ));
  aoi112aa1n03x5               g150(.a(new_n235), .b(new_n239), .c(new_n182), .d(new_n237), .o1(new_n246));
  xorc02aa1n12x5               g151(.a(\a[24] ), .b(\b[23] ), .out0(new_n247));
  oai012aa1n03x5               g152(.a(new_n247), .b(new_n246), .c(new_n242), .o1(new_n248));
  nona22aa1n03x5               g153(.a(new_n244), .b(new_n247), .c(new_n242), .out0(new_n249));
  nanp02aa1n03x5               g154(.a(new_n248), .b(new_n249), .o1(\s[24] ));
  inv040aa1n03x5               g155(.a(new_n236), .o1(new_n251));
  norb02aa1n12x5               g156(.a(new_n247), .b(new_n235), .out0(new_n252));
  nano22aa1n03x7               g157(.a(new_n216), .b(new_n251), .c(new_n252), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n196), .c(new_n190), .d(new_n178), .o1(new_n254));
  and002aa1n02x5               g159(.a(\b[19] ), .b(\a[20] ), .o(new_n255));
  nona23aa1n09x5               g160(.a(new_n221), .b(new_n252), .c(new_n236), .d(new_n255), .out0(new_n256));
  aob012aa1n02x5               g161(.a(new_n241), .b(\b[23] ), .c(\a[24] ), .out0(new_n257));
  oai012aa1n02x5               g162(.a(new_n257), .b(\b[23] ), .c(\a[24] ), .o1(new_n258));
  aoi012aa1n12x5               g163(.a(new_n258), .b(new_n252), .c(new_n238), .o1(new_n259));
  nand02aa1d04x5               g164(.a(new_n256), .b(new_n259), .o1(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  xnrc02aa1n12x5               g166(.a(\b[24] ), .b(\a[25] ), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  xnbna2aa1n03x5               g168(.a(new_n263), .b(new_n254), .c(new_n261), .out0(\s[25] ));
  nor042aa1n09x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n263), .b(new_n260), .c(new_n182), .d(new_n253), .o1(new_n267));
  xnrc02aa1n12x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  tech160nm_fiaoi012aa1n02p5x5 g173(.a(new_n268), .b(new_n267), .c(new_n266), .o1(new_n269));
  tech160nm_fiaoi012aa1n02p5x5 g174(.a(new_n262), .b(new_n254), .c(new_n261), .o1(new_n270));
  nano22aa1n03x5               g175(.a(new_n270), .b(new_n266), .c(new_n268), .out0(new_n271));
  norp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[26] ));
  nor042aa1n09x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  nanp02aa1n02x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  nanb02aa1n06x5               g179(.a(new_n273), .b(new_n274), .out0(new_n275));
  nor042aa1n12x5               g180(.a(new_n268), .b(new_n262), .o1(new_n276));
  nano32aa1d12x5               g181(.a(new_n216), .b(new_n276), .c(new_n251), .d(new_n252), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n196), .c(new_n190), .d(new_n178), .o1(new_n278));
  oao003aa1n09x5               g183(.a(\a[26] ), .b(\b[25] ), .c(new_n266), .carry(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoi012aa1n09x5               g185(.a(new_n280), .b(new_n260), .c(new_n276), .o1(new_n281));
  xobna2aa1n03x5               g186(.a(new_n275), .b(new_n278), .c(new_n281), .out0(\s[27] ));
  inv000aa1d42x5               g187(.a(new_n273), .o1(new_n283));
  xnrc02aa1n12x5               g188(.a(\b[27] ), .b(\a[28] ), .out0(new_n284));
  aoi022aa1n02x7               g189(.a(new_n278), .b(new_n281), .c(\b[26] ), .d(\a[27] ), .o1(new_n285));
  nano22aa1n03x5               g190(.a(new_n285), .b(new_n283), .c(new_n284), .out0(new_n286));
  inv000aa1d42x5               g191(.a(new_n276), .o1(new_n287));
  aoai13aa1n06x5               g192(.a(new_n279), .b(new_n287), .c(new_n256), .d(new_n259), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n274), .b(new_n288), .c(new_n182), .d(new_n277), .o1(new_n289));
  tech160nm_fiaoi012aa1n03p5x5 g194(.a(new_n284), .b(new_n289), .c(new_n283), .o1(new_n290));
  norp02aa1n03x5               g195(.a(new_n290), .b(new_n286), .o1(\s[28] ));
  nor042aa1n04x5               g196(.a(new_n284), .b(new_n275), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n288), .c(new_n182), .d(new_n277), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n283), .carry(new_n294));
  xnrc02aa1n12x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n292), .o1(new_n297));
  tech160nm_fiaoi012aa1n03p5x5 g202(.a(new_n297), .b(new_n278), .c(new_n281), .o1(new_n298));
  nano22aa1n03x7               g203(.a(new_n298), .b(new_n294), .c(new_n295), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n296), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nor043aa1n03x5               g206(.a(new_n295), .b(new_n284), .c(new_n275), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n288), .c(new_n182), .d(new_n277), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[29] ), .b(\a[30] ), .out0(new_n305));
  tech160nm_fiaoi012aa1n02p5x5 g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n302), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n307), .b(new_n278), .c(new_n281), .o1(new_n308));
  nano22aa1n03x5               g213(.a(new_n308), .b(new_n304), .c(new_n305), .out0(new_n309));
  norp02aa1n03x5               g214(.a(new_n306), .b(new_n309), .o1(\s[30] ));
  xnrc02aa1n02x5               g215(.a(\b[30] ), .b(\a[31] ), .out0(new_n311));
  norb03aa1n09x5               g216(.a(new_n292), .b(new_n305), .c(new_n295), .out0(new_n312));
  inv000aa1n02x5               g217(.a(new_n312), .o1(new_n313));
  tech160nm_fiaoi012aa1n03p5x5 g218(.a(new_n313), .b(new_n278), .c(new_n281), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n304), .carry(new_n315));
  nano22aa1n03x7               g220(.a(new_n314), .b(new_n311), .c(new_n315), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n312), .b(new_n288), .c(new_n182), .d(new_n277), .o1(new_n317));
  tech160nm_fiaoi012aa1n02p5x5 g222(.a(new_n311), .b(new_n317), .c(new_n315), .o1(new_n318));
  norp02aa1n03x5               g223(.a(new_n318), .b(new_n316), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n101), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g228(.a(new_n119), .b(new_n112), .out0(new_n324));
  oai112aa1n02x5               g229(.a(new_n107), .b(new_n324), .c(new_n106), .d(new_n101), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[6] ), .b(\b[5] ), .out0(new_n326));
  xobna2aa1n03x5               g231(.a(new_n326), .b(new_n325), .c(new_n119), .out0(\s[6] ));
  norp02aa1n02x5               g232(.a(\b[5] ), .b(\a[6] ), .o1(new_n328));
  aoi013aa1n02x4               g233(.a(new_n328), .b(new_n325), .c(new_n119), .d(new_n109), .o1(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g235(.a(\a[7] ), .b(\b[6] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g237(.a(new_n190), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


