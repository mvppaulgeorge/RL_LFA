// Benchmark "adder" written by ABC on Wed Jul 17 17:30:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n355, new_n357, new_n358, new_n360,
    new_n361, new_n364, new_n366, new_n367, new_n368, new_n370;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n12x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nor002aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  tech160nm_finand02aa1n03p5x5 g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  norb03aa1n03x5               g006(.a(new_n101), .b(new_n99), .c(new_n100), .out0(new_n102));
  norp02aa1n12x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  aoi022aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .c(\a[3] ), .d(\b[2] ), .o1(new_n105));
  nona23aa1n06x5               g010(.a(new_n105), .b(new_n101), .c(new_n103), .d(new_n104), .out0(new_n106));
  aob012aa1n02x5               g011(.a(new_n104), .b(\b[3] ), .c(\a[4] ), .out0(new_n107));
  norb02aa1n06x4               g012(.a(new_n107), .b(new_n103), .out0(new_n108));
  tech160nm_fioai012aa1n03p5x5 g013(.a(new_n108), .b(new_n106), .c(new_n102), .o1(new_n109));
  xnrc02aa1n12x5               g014(.a(\b[6] ), .b(\a[7] ), .out0(new_n110));
  nor022aa1n06x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  norb02aa1n02x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nor002aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand42aa1n08x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  norb02aa1n03x4               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  tech160nm_fixorc02aa1n02p5x5 g021(.a(\a[8] ), .b(\b[7] ), .out0(new_n117));
  nano32aa1n03x7               g022(.a(new_n110), .b(new_n117), .c(new_n113), .d(new_n116), .out0(new_n118));
  aoi022aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n119));
  tech160nm_fioai012aa1n04x5   g024(.a(new_n119), .b(new_n114), .c(new_n111), .o1(new_n120));
  oa0022aa1n06x5               g025(.a(\a[8] ), .b(\b[7] ), .c(\a[7] ), .d(\b[6] ), .o(new_n121));
  aoi022aa1d18x5               g026(.a(new_n120), .b(new_n121), .c(\b[7] ), .d(\a[8] ), .o1(new_n122));
  nand42aa1n03x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  norb02aa1n02x5               g028(.a(new_n123), .b(new_n97), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n122), .c(new_n118), .d(new_n109), .o1(new_n125));
  nor042aa1n04x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand02aa1n06x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  inv030aa1n04x5               g034(.a(new_n102), .o1(new_n130));
  nanb02aa1n06x5               g035(.a(new_n106), .b(new_n130), .out0(new_n131));
  nanb02aa1n02x5               g036(.a(new_n111), .b(new_n112), .out0(new_n132));
  nona23aa1n06x5               g037(.a(new_n117), .b(new_n116), .c(new_n110), .d(new_n132), .out0(new_n133));
  inv040aa1n06x5               g038(.a(new_n122), .o1(new_n134));
  aoai13aa1n12x5               g039(.a(new_n134), .b(new_n133), .c(new_n131), .d(new_n108), .o1(new_n135));
  aoai13aa1n06x5               g040(.a(new_n128), .b(new_n97), .c(new_n135), .d(new_n124), .o1(new_n136));
  oaoi03aa1n02x5               g041(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  nand42aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  inv000aa1d42x5               g044(.a(\b[10] ), .o1(new_n140));
  nanb02aa1d24x5               g045(.a(\a[11] ), .b(new_n140), .out0(new_n141));
  nand22aa1n03x5               g046(.a(new_n141), .b(new_n139), .o1(new_n142));
  xobna2aa1n03x5               g047(.a(new_n142), .b(new_n136), .c(new_n138), .out0(\s[11] ));
  oaoi13aa1n02x5               g048(.a(new_n142), .b(new_n127), .c(new_n97), .d(new_n126), .o1(new_n144));
  aoi022aa1n02x5               g049(.a(new_n136), .b(new_n144), .c(\b[10] ), .d(\a[11] ), .o1(new_n145));
  norp02aa1n02x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  and002aa1n12x5               g051(.a(\b[11] ), .b(\a[12] ), .o(new_n147));
  norp02aa1n02x5               g052(.a(new_n147), .b(new_n146), .o1(new_n148));
  aoi012aa1n02x5               g053(.a(new_n148), .b(\a[11] ), .c(\b[10] ), .o1(new_n149));
  aob012aa1n02x5               g054(.a(new_n149), .b(new_n136), .c(new_n144), .out0(new_n150));
  oaib12aa1n02x5               g055(.a(new_n150), .b(new_n145), .c(new_n148), .out0(\s[12] ));
  nano23aa1n06x5               g056(.a(new_n97), .b(new_n126), .c(new_n127), .d(new_n123), .out0(new_n152));
  nona32aa1d18x5               g057(.a(new_n152), .b(new_n142), .c(new_n147), .d(new_n146), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n122), .c(new_n118), .d(new_n109), .o1(new_n155));
  oai022aa1n02x5               g060(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n156));
  nor002aa1n02x5               g061(.a(new_n156), .b(new_n147), .o1(new_n157));
  oai112aa1n04x5               g062(.a(new_n127), .b(new_n139), .c(new_n126), .d(new_n97), .o1(new_n158));
  oaoi03aa1n02x5               g063(.a(\a[12] ), .b(\b[11] ), .c(new_n141), .o1(new_n159));
  inv000aa1n02x5               g064(.a(new_n159), .o1(new_n160));
  oaib12aa1n06x5               g065(.a(new_n160), .b(new_n158), .c(new_n157), .out0(new_n161));
  nanb02aa1n03x5               g066(.a(new_n161), .b(new_n155), .out0(new_n162));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nor022aa1n06x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  nand42aa1n02x5               g070(.a(new_n139), .b(new_n127), .o1(new_n166));
  oab012aa1n06x5               g071(.a(new_n166), .b(new_n97), .c(new_n126), .out0(new_n167));
  aoi112aa1n02x5               g072(.a(new_n159), .b(new_n165), .c(new_n167), .d(new_n157), .o1(new_n168));
  aoi022aa1n02x5               g073(.a(new_n162), .b(new_n165), .c(new_n155), .d(new_n168), .o1(\s[13] ));
  nor042aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  aoi112aa1n02x5               g077(.a(new_n164), .b(new_n172), .c(new_n162), .d(new_n165), .o1(new_n173));
  aoai13aa1n02x5               g078(.a(new_n172), .b(new_n164), .c(new_n162), .d(new_n163), .o1(new_n174));
  norb02aa1n03x4               g079(.a(new_n174), .b(new_n173), .out0(\s[14] ));
  nano23aa1n06x5               g080(.a(new_n170), .b(new_n164), .c(new_n171), .d(new_n163), .out0(new_n176));
  aoai13aa1n03x5               g081(.a(new_n176), .b(new_n161), .c(new_n135), .d(new_n154), .o1(new_n177));
  tech160nm_fioai012aa1n04x5   g082(.a(new_n171), .b(new_n170), .c(new_n164), .o1(new_n178));
  xnrc02aa1n12x5               g083(.a(\b[14] ), .b(\a[15] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n177), .c(new_n178), .out0(\s[15] ));
  inv000aa1n02x5               g086(.a(new_n178), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n180), .b(new_n182), .c(new_n162), .d(new_n176), .o1(new_n183));
  xorc02aa1n02x5               g088(.a(\a[16] ), .b(\b[15] ), .out0(new_n184));
  nor042aa1n04x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[16] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[15] ), .o1(new_n187));
  nanp02aa1n02x5               g092(.a(new_n187), .b(new_n186), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  aoi012aa1n02x5               g094(.a(new_n185), .b(new_n188), .c(new_n189), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n185), .o1(new_n191));
  aoai13aa1n02x5               g096(.a(new_n191), .b(new_n179), .c(new_n177), .d(new_n178), .o1(new_n192));
  aoi022aa1n02x5               g097(.a(new_n192), .b(new_n184), .c(new_n183), .d(new_n190), .o1(\s[16] ));
  norp02aa1n12x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  and002aa1n06x5               g099(.a(\b[16] ), .b(\a[17] ), .o(new_n195));
  nano22aa1d15x5               g100(.a(new_n179), .b(new_n188), .c(new_n189), .out0(new_n196));
  nano22aa1d15x5               g101(.a(new_n153), .b(new_n176), .c(new_n196), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n122), .c(new_n109), .d(new_n118), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n196), .o1(new_n199));
  aoai13aa1n06x5               g104(.a(new_n176), .b(new_n159), .c(new_n167), .d(new_n157), .o1(new_n200));
  oaoi03aa1n02x5               g105(.a(new_n186), .b(new_n187), .c(new_n185), .o1(new_n201));
  aoai13aa1n04x5               g106(.a(new_n201), .b(new_n199), .c(new_n200), .d(new_n178), .o1(new_n202));
  obai22aa1n02x7               g107(.a(new_n198), .b(new_n202), .c(new_n194), .d(new_n195), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n196), .b(new_n182), .c(new_n161), .d(new_n176), .o1(new_n204));
  oai022aa1n02x5               g109(.a(\a[16] ), .b(\b[15] ), .c(\b[16] ), .d(\a[17] ), .o1(new_n205));
  aoi112aa1n02x5               g110(.a(new_n205), .b(new_n195), .c(new_n185), .d(new_n189), .o1(new_n206));
  nanp03aa1n02x5               g111(.a(new_n198), .b(new_n204), .c(new_n206), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n203), .b(new_n207), .o1(\s[17] ));
  inv000aa1d42x5               g113(.a(new_n195), .o1(new_n209));
  nor022aa1n08x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nand02aa1n06x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nanb02aa1n06x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n207), .c(new_n209), .out0(\s[18] ));
  nor043aa1n06x5               g118(.a(new_n212), .b(new_n195), .c(new_n194), .o1(new_n214));
  aoai13aa1n06x5               g119(.a(new_n214), .b(new_n202), .c(new_n135), .d(new_n197), .o1(new_n215));
  oa0012aa1n02x5               g120(.a(new_n211), .b(new_n210), .c(new_n194), .o(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  nanp02aa1n04x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nor042aa1d18x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  norb02aa1n09x5               g124(.a(new_n218), .b(new_n219), .out0(new_n220));
  xnbna2aa1n03x5               g125(.a(new_n220), .b(new_n215), .c(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand23aa1n06x5               g127(.a(new_n198), .b(new_n204), .c(new_n201), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n220), .b(new_n216), .c(new_n223), .d(new_n214), .o1(new_n224));
  nor002aa1d32x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand02aa1d10x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n09x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  inv030aa1n04x5               g132(.a(new_n225), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n219), .b(new_n228), .c(new_n226), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n219), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n220), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n230), .b(new_n231), .c(new_n215), .d(new_n217), .o1(new_n232));
  aoi022aa1n03x5               g137(.a(new_n232), .b(new_n227), .c(new_n224), .d(new_n229), .o1(\s[20] ));
  nand23aa1d12x5               g138(.a(new_n214), .b(new_n220), .c(new_n227), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n202), .c(new_n135), .d(new_n197), .o1(new_n236));
  oai112aa1n06x5               g141(.a(new_n228), .b(new_n226), .c(\b[18] ), .d(\a[19] ), .o1(new_n237));
  oai112aa1n06x5               g142(.a(new_n211), .b(new_n218), .c(new_n210), .d(new_n194), .o1(new_n238));
  aoi012aa1n12x5               g143(.a(new_n225), .b(new_n219), .c(new_n226), .o1(new_n239));
  oai012aa1n18x5               g144(.a(new_n239), .b(new_n238), .c(new_n237), .o1(new_n240));
  nand42aa1n02x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  nor002aa1n20x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  norb02aa1n06x5               g147(.a(new_n241), .b(new_n242), .out0(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n240), .c(new_n223), .d(new_n235), .o1(new_n244));
  norb03aa1n09x5               g149(.a(new_n226), .b(new_n219), .c(new_n225), .out0(new_n245));
  nand42aa1n03x5               g150(.a(new_n218), .b(new_n211), .o1(new_n246));
  oab012aa1n06x5               g151(.a(new_n246), .b(new_n194), .c(new_n210), .out0(new_n247));
  inv020aa1n03x5               g152(.a(new_n239), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n248), .b(new_n243), .c(new_n247), .d(new_n245), .o1(new_n249));
  aobi12aa1n03x7               g154(.a(new_n244), .b(new_n249), .c(new_n236), .out0(\s[21] ));
  nor042aa1n04x5               g155(.a(\b[21] ), .b(\a[22] ), .o1(new_n251));
  nand02aa1n08x5               g156(.a(\b[21] ), .b(\a[22] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  norp02aa1n02x5               g158(.a(new_n253), .b(new_n242), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n240), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n242), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n243), .o1(new_n257));
  aoai13aa1n02x5               g162(.a(new_n256), .b(new_n257), .c(new_n236), .d(new_n255), .o1(new_n258));
  aoi022aa1n02x7               g163(.a(new_n258), .b(new_n253), .c(new_n244), .d(new_n254), .o1(\s[22] ));
  nano22aa1n02x4               g164(.a(new_n234), .b(new_n243), .c(new_n253), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n202), .c(new_n135), .d(new_n197), .o1(new_n261));
  nano23aa1n09x5               g166(.a(new_n251), .b(new_n242), .c(new_n252), .d(new_n241), .out0(new_n262));
  aoi012aa1d24x5               g167(.a(new_n251), .b(new_n242), .c(new_n252), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aoi012aa1n02x5               g169(.a(new_n264), .b(new_n240), .c(new_n262), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(new_n261), .b(new_n265), .o1(new_n266));
  nor042aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .o1(new_n267));
  and002aa1n12x5               g172(.a(\b[22] ), .b(\a[23] ), .o(new_n268));
  nor042aa1n04x5               g173(.a(new_n268), .b(new_n267), .o1(new_n269));
  aoi112aa1n02x5               g174(.a(new_n269), .b(new_n264), .c(new_n240), .d(new_n262), .o1(new_n270));
  aoi022aa1n02x5               g175(.a(new_n266), .b(new_n269), .c(new_n261), .d(new_n270), .o1(\s[23] ));
  aoai13aa1n06x5               g176(.a(new_n262), .b(new_n248), .c(new_n247), .d(new_n245), .o1(new_n272));
  aoi112aa1n02x5               g177(.a(new_n251), .b(new_n267), .c(new_n242), .d(new_n252), .o1(new_n273));
  nanp02aa1n02x5               g178(.a(new_n272), .b(new_n273), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n274), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[24] ), .b(\b[23] ), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n268), .c(new_n261), .d(new_n275), .o1(new_n277));
  orn002aa1n02x5               g182(.a(new_n276), .b(new_n268), .o(new_n278));
  aoai13aa1n03x5               g183(.a(new_n277), .b(new_n278), .c(new_n275), .d(new_n261), .o1(\s[24] ));
  nano32aa1n02x5               g184(.a(new_n234), .b(new_n276), .c(new_n262), .d(new_n269), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n202), .c(new_n135), .d(new_n197), .o1(new_n281));
  and002aa1n06x5               g186(.a(new_n276), .b(new_n269), .o(new_n282));
  inv030aa1n02x5               g187(.a(new_n282), .o1(new_n283));
  orn002aa1n02x5               g188(.a(\a[23] ), .b(\b[22] ), .o(new_n284));
  oao003aa1n02x5               g189(.a(\a[24] ), .b(\b[23] ), .c(new_n284), .carry(new_n285));
  aoai13aa1n12x5               g190(.a(new_n285), .b(new_n283), .c(new_n272), .d(new_n263), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[25] ), .b(\b[24] ), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n287), .b(new_n286), .c(new_n223), .d(new_n280), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n282), .b(new_n264), .c(new_n240), .d(new_n262), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n287), .o1(new_n290));
  and003aa1n02x5               g195(.a(new_n289), .b(new_n290), .c(new_n285), .o(new_n291));
  aobi12aa1n03x7               g196(.a(new_n288), .b(new_n291), .c(new_n281), .out0(\s[25] ));
  xorc02aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .out0(new_n293));
  nor042aa1n03x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  norp02aa1n02x5               g199(.a(new_n293), .b(new_n294), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n286), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n294), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n290), .c(new_n281), .d(new_n296), .o1(new_n298));
  aoi022aa1n02x7               g203(.a(new_n298), .b(new_n293), .c(new_n288), .d(new_n295), .o1(\s[26] ));
  and002aa1n12x5               g204(.a(new_n293), .b(new_n287), .o(new_n300));
  nano23aa1n06x5               g205(.a(new_n283), .b(new_n234), .c(new_n300), .d(new_n262), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n202), .c(new_n135), .d(new_n197), .o1(new_n302));
  nor042aa1n04x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  and002aa1n12x5               g208(.a(\b[26] ), .b(\a[27] ), .o(new_n304));
  nor042aa1n03x5               g209(.a(new_n304), .b(new_n303), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[26] ), .b(\b[25] ), .c(new_n297), .carry(new_n306));
  inv000aa1d42x5               g211(.a(new_n306), .o1(new_n307));
  aoi112aa1n02x5               g212(.a(new_n307), .b(new_n305), .c(new_n286), .d(new_n300), .o1(new_n308));
  aoi012aa1n12x5               g213(.a(new_n307), .b(new_n286), .c(new_n300), .o1(new_n309));
  nanp02aa1n02x5               g214(.a(new_n302), .b(new_n309), .o1(new_n310));
  aoi022aa1n02x5               g215(.a(new_n310), .b(new_n305), .c(new_n302), .d(new_n308), .o1(\s[27] ));
  inv000aa1d42x5               g216(.a(new_n304), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n300), .o1(new_n313));
  aoai13aa1n04x5               g218(.a(new_n306), .b(new_n313), .c(new_n289), .d(new_n285), .o1(new_n314));
  aoai13aa1n02x5               g219(.a(new_n312), .b(new_n314), .c(new_n223), .d(new_n301), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .out0(new_n316));
  norp02aa1n02x5               g221(.a(new_n316), .b(new_n303), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n303), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n304), .c(new_n302), .d(new_n309), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n319), .b(new_n316), .c(new_n315), .d(new_n317), .o1(\s[28] ));
  and002aa1n03x5               g225(.a(new_n316), .b(new_n305), .o(new_n321));
  aoai13aa1n02x5               g226(.a(new_n321), .b(new_n314), .c(new_n223), .d(new_n301), .o1(new_n322));
  inv020aa1n02x5               g227(.a(new_n321), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[28] ), .b(\b[27] ), .c(new_n318), .carry(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n323), .c(new_n302), .d(new_n309), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n324), .b(new_n326), .out0(new_n327));
  aoi022aa1n03x5               g232(.a(new_n325), .b(new_n326), .c(new_n322), .d(new_n327), .o1(\s[29] ));
  xorb03aa1n02x5               g233(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g234(.a(new_n316), .b(new_n326), .c(new_n305), .o(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n314), .c(new_n223), .d(new_n301), .o1(new_n331));
  inv000aa1d42x5               g236(.a(new_n330), .o1(new_n332));
  inv000aa1d42x5               g237(.a(\b[28] ), .o1(new_n333));
  inv000aa1d42x5               g238(.a(\a[29] ), .o1(new_n334));
  oaib12aa1n02x5               g239(.a(new_n324), .b(\b[28] ), .c(new_n334), .out0(new_n335));
  oaib12aa1n02x5               g240(.a(new_n335), .b(new_n333), .c(\a[29] ), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n332), .c(new_n302), .d(new_n309), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[30] ), .b(\b[29] ), .out0(new_n338));
  oaoi13aa1n02x5               g243(.a(new_n338), .b(new_n335), .c(new_n334), .d(new_n333), .o1(new_n339));
  aoi022aa1n03x5               g244(.a(new_n337), .b(new_n338), .c(new_n331), .d(new_n339), .o1(\s[30] ));
  nanb02aa1n02x5               g245(.a(\b[30] ), .b(\a[31] ), .out0(new_n341));
  nanb02aa1n02x5               g246(.a(\a[31] ), .b(\b[30] ), .out0(new_n342));
  nanp02aa1n02x5               g247(.a(new_n342), .b(new_n341), .o1(new_n343));
  nano22aa1d24x5               g248(.a(new_n323), .b(new_n326), .c(new_n338), .out0(new_n344));
  aoai13aa1n02x5               g249(.a(new_n344), .b(new_n314), .c(new_n223), .d(new_n301), .o1(new_n345));
  inv000aa1d42x5               g250(.a(new_n344), .o1(new_n346));
  norp02aa1n02x5               g251(.a(\b[29] ), .b(\a[30] ), .o1(new_n347));
  aoi022aa1n02x5               g252(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n348));
  aoi012aa1n02x5               g253(.a(new_n347), .b(new_n335), .c(new_n348), .o1(new_n349));
  aoai13aa1n03x5               g254(.a(new_n349), .b(new_n346), .c(new_n302), .d(new_n309), .o1(new_n350));
  oai112aa1n02x5               g255(.a(new_n341), .b(new_n342), .c(\b[29] ), .d(\a[30] ), .o1(new_n351));
  aoi012aa1n02x5               g256(.a(new_n351), .b(new_n335), .c(new_n348), .o1(new_n352));
  aoi022aa1n03x5               g257(.a(new_n350), .b(new_n343), .c(new_n345), .d(new_n352), .o1(\s[31] ));
  nanp02aa1n02x5               g258(.a(\b[2] ), .b(\a[3] ), .o1(new_n354));
  norb02aa1n02x5               g259(.a(new_n354), .b(new_n104), .out0(new_n355));
  xobna2aa1n03x5               g260(.a(new_n355), .b(new_n130), .c(new_n101), .out0(\s[3] ));
  aoai13aa1n02x5               g261(.a(new_n355), .b(new_n102), .c(\a[2] ), .d(\b[1] ), .o1(new_n357));
  xnrc02aa1n02x5               g262(.a(\b[3] ), .b(\a[4] ), .out0(new_n358));
  xnbna2aa1n03x5               g263(.a(new_n358), .b(new_n357), .c(new_n354), .out0(\s[4] ));
  nona23aa1n02x4               g264(.a(new_n107), .b(new_n115), .c(new_n114), .d(new_n103), .out0(new_n360));
  oabi12aa1n02x5               g265(.a(new_n360), .b(new_n102), .c(new_n106), .out0(new_n361));
  aoai13aa1n02x5               g266(.a(new_n361), .b(new_n116), .c(new_n131), .d(new_n108), .o1(\s[5] ));
  xnbna2aa1n03x5               g267(.a(new_n132), .b(new_n361), .c(new_n115), .out0(\s[6] ));
  aob012aa1n02x5               g268(.a(new_n113), .b(new_n361), .c(new_n115), .out0(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n110), .b(new_n364), .c(new_n112), .out0(\s[7] ));
  aoi012aa1n02x5               g270(.a(new_n110), .b(new_n364), .c(new_n112), .o1(new_n366));
  aoai13aa1n02x5               g271(.a(new_n117), .b(new_n366), .c(\b[6] ), .d(\a[7] ), .o1(new_n367));
  aoi012aa1n02x5               g272(.a(new_n117), .b(\a[7] ), .c(\b[6] ), .o1(new_n368));
  oaib12aa1n02x5               g273(.a(new_n367), .b(new_n366), .c(new_n368), .out0(\s[8] ));
  aoi112aa1n02x5               g274(.a(new_n122), .b(new_n124), .c(new_n118), .d(new_n109), .o1(new_n370));
  aoi012aa1n02x5               g275(.a(new_n370), .b(new_n135), .c(new_n124), .o1(\s[9] ));
endmodule


