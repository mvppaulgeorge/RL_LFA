// Benchmark "adder" written by ABC on Wed Jul 17 18:07:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n302, new_n305,
    new_n307, new_n308, new_n310, new_n312;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nand02aa1d04x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  nor022aa1n06x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nona23aa1n09x5               g008(.a(new_n103), .b(new_n101), .c(new_n100), .d(new_n102), .out0(new_n104));
  norp02aa1n12x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nand02aa1d06x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nand02aa1n04x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nona23aa1d18x5               g013(.a(new_n108), .b(new_n106), .c(new_n105), .d(new_n107), .out0(new_n109));
  nor042aa1n04x5               g014(.a(new_n109), .b(new_n104), .o1(new_n110));
  and002aa1n02x5               g015(.a(\b[3] ), .b(\a[4] ), .o(new_n111));
  oa0022aa1n02x5               g016(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n112));
  inv040aa1d32x5               g017(.a(\a[3] ), .o1(new_n113));
  inv040aa1d28x5               g018(.a(\b[2] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(new_n114), .b(new_n113), .o1(new_n115));
  nand42aa1n03x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nand02aa1n02x5               g021(.a(new_n115), .b(new_n116), .o1(new_n117));
  nand42aa1n04x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  nor042aa1d18x5               g023(.a(\b[1] ), .b(\a[2] ), .o1(new_n119));
  nand42aa1n16x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  oai012aa1n12x5               g025(.a(new_n118), .b(new_n119), .c(new_n120), .o1(new_n121));
  oaoi13aa1n12x5               g026(.a(new_n111), .b(new_n112), .c(new_n121), .d(new_n117), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n100), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n102), .b(new_n101), .o1(new_n124));
  aoi012aa1n06x5               g029(.a(new_n105), .b(new_n107), .c(new_n106), .o1(new_n125));
  oai112aa1n06x5               g030(.a(new_n123), .b(new_n124), .c(new_n104), .d(new_n125), .o1(new_n126));
  tech160nm_fixorc02aa1n03p5x5 g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n97), .b(new_n128), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g034(.a(new_n97), .o1(new_n130));
  aoi112aa1n03x5               g035(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n131));
  oab012aa1n06x5               g036(.a(new_n131), .b(\a[10] ), .c(\b[9] ), .out0(new_n132));
  aoai13aa1n04x5               g037(.a(new_n132), .b(new_n130), .c(new_n128), .d(new_n99), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand02aa1n06x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nor002aa1n06x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand02aa1n06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  aoi112aa1n02x5               g044(.a(new_n139), .b(new_n135), .c(new_n133), .d(new_n136), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n139), .b(new_n135), .c(new_n133), .d(new_n136), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(\s[12] ));
  nona23aa1n09x5               g047(.a(new_n138), .b(new_n136), .c(new_n135), .d(new_n137), .out0(new_n143));
  nano22aa1n02x4               g048(.a(new_n143), .b(new_n97), .c(new_n127), .out0(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n145));
  aoi012aa1n06x5               g050(.a(new_n137), .b(new_n135), .c(new_n138), .o1(new_n146));
  oai012aa1d24x5               g051(.a(new_n146), .b(new_n143), .c(new_n132), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n145), .b(new_n148), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n04x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  tech160nm_finand02aa1n03p5x5 g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  aoi012aa1n02x5               g057(.a(new_n151), .b(new_n149), .c(new_n152), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nanp02aa1n04x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nona23aa1n03x5               g061(.a(new_n156), .b(new_n152), .c(new_n151), .d(new_n155), .out0(new_n157));
  tech160nm_fiaoi012aa1n05x5   g062(.a(new_n155), .b(new_n151), .c(new_n156), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n157), .c(new_n145), .d(new_n148), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n03x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  tech160nm_fixorc02aa1n02p5x5 g066(.a(\a[15] ), .b(\b[14] ), .out0(new_n162));
  xorc02aa1n02x5               g067(.a(\a[16] ), .b(\b[15] ), .out0(new_n163));
  aoi112aa1n02x5               g068(.a(new_n163), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n164));
  aoai13aa1n02x7               g069(.a(new_n163), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n165));
  norb02aa1n03x4               g070(.a(new_n165), .b(new_n164), .out0(\s[16] ));
  nano23aa1n02x5               g071(.a(new_n135), .b(new_n137), .c(new_n138), .d(new_n136), .out0(new_n167));
  nano23aa1n02x4               g072(.a(new_n151), .b(new_n155), .c(new_n156), .d(new_n152), .out0(new_n168));
  nanp03aa1n02x5               g073(.a(new_n168), .b(new_n162), .c(new_n163), .o1(new_n169));
  nano32aa1n03x7               g074(.a(new_n169), .b(new_n167), .c(new_n127), .d(new_n97), .out0(new_n170));
  aoai13aa1n12x5               g075(.a(new_n170), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n171));
  xnrc02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .out0(new_n172));
  xnrc02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .out0(new_n173));
  nor043aa1n02x5               g078(.a(new_n157), .b(new_n173), .c(new_n172), .o1(new_n174));
  aob012aa1n02x5               g079(.a(new_n161), .b(\b[15] ), .c(\a[16] ), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  nanb03aa1n03x5               g081(.a(new_n158), .b(new_n163), .c(new_n162), .out0(new_n177));
  tech160nm_fioai012aa1n04x5   g082(.a(new_n177), .b(\b[15] ), .c(\a[16] ), .o1(new_n178));
  aoi112aa1n09x5               g083(.a(new_n178), .b(new_n176), .c(new_n147), .d(new_n174), .o1(new_n179));
  nand02aa1d08x5               g084(.a(new_n171), .b(new_n179), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g086(.a(\a[18] ), .o1(new_n182));
  inv040aa1d30x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(new_n183), .b(new_n184), .c(new_n180), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n182), .out0(\s[18] ));
  xroi22aa1d06x4               g091(.a(new_n183), .b(\b[16] ), .c(new_n182), .d(\b[17] ), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  norp02aa1n02x5               g093(.a(\b[17] ), .b(\a[18] ), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(\b[17] ), .b(\a[18] ), .o1(new_n190));
  aoi013aa1n06x4               g095(.a(new_n189), .b(new_n190), .c(new_n183), .d(new_n184), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n188), .c(new_n171), .d(new_n179), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g098(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n06x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand42aa1n06x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nor022aa1n06x5               g101(.a(\b[19] ), .b(\a[20] ), .o1(new_n197));
  nand42aa1n06x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  aoi112aa1n02x5               g104(.a(new_n195), .b(new_n199), .c(new_n192), .d(new_n196), .o1(new_n200));
  aoai13aa1n03x5               g105(.a(new_n199), .b(new_n195), .c(new_n192), .d(new_n196), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(\s[20] ));
  nano23aa1n03x5               g107(.a(new_n195), .b(new_n197), .c(new_n198), .d(new_n196), .out0(new_n203));
  nand02aa1n02x5               g108(.a(new_n187), .b(new_n203), .o1(new_n204));
  nona23aa1n03x5               g109(.a(new_n198), .b(new_n196), .c(new_n195), .d(new_n197), .out0(new_n205));
  tech160nm_fioai012aa1n04x5   g110(.a(new_n198), .b(new_n197), .c(new_n195), .o1(new_n206));
  oai012aa1n12x5               g111(.a(new_n206), .b(new_n205), .c(new_n191), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n204), .c(new_n171), .d(new_n179), .o1(new_n209));
  xorb03aa1n02x5               g114(.a(new_n209), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g115(.a(\b[20] ), .b(\a[21] ), .o1(new_n211));
  xorc02aa1n02x5               g116(.a(\a[21] ), .b(\b[20] ), .out0(new_n212));
  xorc02aa1n02x5               g117(.a(\a[22] ), .b(\b[21] ), .out0(new_n213));
  aoi112aa1n03x5               g118(.a(new_n211), .b(new_n213), .c(new_n209), .d(new_n212), .o1(new_n214));
  aoai13aa1n03x5               g119(.a(new_n213), .b(new_n211), .c(new_n209), .d(new_n212), .o1(new_n215));
  norb02aa1n02x7               g120(.a(new_n215), .b(new_n214), .out0(\s[22] ));
  inv000aa1d42x5               g121(.a(\a[21] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\a[22] ), .o1(new_n218));
  xroi22aa1d06x4               g123(.a(new_n217), .b(\b[20] ), .c(new_n218), .d(\b[21] ), .out0(new_n219));
  nanp03aa1n02x5               g124(.a(new_n219), .b(new_n187), .c(new_n203), .o1(new_n220));
  inv000aa1d42x5               g125(.a(\b[21] ), .o1(new_n221));
  oao003aa1n02x5               g126(.a(new_n218), .b(new_n221), .c(new_n211), .carry(new_n222));
  aoi012aa1n02x5               g127(.a(new_n222), .b(new_n207), .c(new_n219), .o1(new_n223));
  aoai13aa1n06x5               g128(.a(new_n223), .b(new_n220), .c(new_n171), .d(new_n179), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g130(.a(\b[22] ), .b(\a[23] ), .o1(new_n226));
  xorc02aa1n02x5               g131(.a(\a[23] ), .b(\b[22] ), .out0(new_n227));
  xorc02aa1n02x5               g132(.a(\a[24] ), .b(\b[23] ), .out0(new_n228));
  aoi112aa1n02x5               g133(.a(new_n226), .b(new_n228), .c(new_n224), .d(new_n227), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n228), .b(new_n226), .c(new_n224), .d(new_n227), .o1(new_n230));
  norb02aa1n02x7               g135(.a(new_n230), .b(new_n229), .out0(\s[24] ));
  inv000aa1d42x5               g136(.a(\a[23] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\a[24] ), .o1(new_n233));
  xroi22aa1d06x4               g138(.a(new_n232), .b(\b[22] ), .c(new_n233), .d(\b[23] ), .out0(new_n234));
  nano22aa1n02x5               g139(.a(new_n204), .b(new_n219), .c(new_n234), .out0(new_n235));
  nona22aa1n02x4               g140(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(new_n236));
  oaib12aa1n02x5               g141(.a(new_n236), .b(\b[17] ), .c(new_n182), .out0(new_n237));
  inv040aa1n03x5               g142(.a(new_n206), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n219), .b(new_n238), .c(new_n203), .d(new_n237), .o1(new_n239));
  inv040aa1n02x5               g144(.a(new_n222), .o1(new_n240));
  inv000aa1n02x5               g145(.a(new_n234), .o1(new_n241));
  oai022aa1n02x5               g146(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n242));
  oaib12aa1n02x5               g147(.a(new_n242), .b(new_n233), .c(\b[23] ), .out0(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n241), .c(new_n239), .d(new_n240), .o1(new_n244));
  xorc02aa1n02x5               g149(.a(\a[25] ), .b(\b[24] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n244), .c(new_n180), .d(new_n235), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n245), .b(new_n244), .c(new_n180), .d(new_n235), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[26] ), .b(\b[25] ), .out0(new_n250));
  nona22aa1n02x5               g155(.a(new_n246), .b(new_n250), .c(new_n249), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n249), .o1(new_n252));
  aobi12aa1n06x5               g157(.a(new_n250), .b(new_n246), .c(new_n252), .out0(new_n253));
  norb02aa1n03x4               g158(.a(new_n251), .b(new_n253), .out0(\s[26] ));
  inv000aa1d42x5               g159(.a(\a[25] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(\a[26] ), .o1(new_n256));
  xroi22aa1d06x4               g161(.a(new_n255), .b(\b[24] ), .c(new_n256), .d(\b[25] ), .out0(new_n257));
  nano32aa1n03x7               g162(.a(new_n204), .b(new_n257), .c(new_n219), .d(new_n234), .out0(new_n258));
  nand02aa1d06x5               g163(.a(new_n180), .b(new_n258), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .c(new_n252), .carry(new_n260));
  aobi12aa1n06x5               g165(.a(new_n260), .b(new_n244), .c(new_n257), .out0(new_n261));
  xorc02aa1n02x5               g166(.a(\a[27] ), .b(\b[26] ), .out0(new_n262));
  xnbna2aa1n03x5               g167(.a(new_n262), .b(new_n261), .c(new_n259), .out0(\s[27] ));
  norp02aa1n02x5               g168(.a(\b[26] ), .b(\a[27] ), .o1(new_n264));
  inv040aa1n03x5               g169(.a(new_n264), .o1(new_n265));
  aobi12aa1n06x5               g170(.a(new_n262), .b(new_n261), .c(new_n259), .out0(new_n266));
  xnrc02aa1n02x5               g171(.a(\b[27] ), .b(\a[28] ), .out0(new_n267));
  nano22aa1n03x7               g172(.a(new_n266), .b(new_n265), .c(new_n267), .out0(new_n268));
  aobi12aa1n06x5               g173(.a(new_n258), .b(new_n171), .c(new_n179), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n234), .b(new_n222), .c(new_n207), .d(new_n219), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n257), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n260), .b(new_n271), .c(new_n270), .d(new_n243), .o1(new_n272));
  oaih12aa1n02x5               g177(.a(new_n262), .b(new_n272), .c(new_n269), .o1(new_n273));
  tech160nm_fiaoi012aa1n02p5x5 g178(.a(new_n267), .b(new_n273), .c(new_n265), .o1(new_n274));
  nor002aa1n02x5               g179(.a(new_n274), .b(new_n268), .o1(\s[28] ));
  norb02aa1n02x5               g180(.a(new_n262), .b(new_n267), .out0(new_n276));
  aobi12aa1n02x7               g181(.a(new_n276), .b(new_n261), .c(new_n259), .out0(new_n277));
  oao003aa1n02x5               g182(.a(\a[28] ), .b(\b[27] ), .c(new_n265), .carry(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[28] ), .b(\a[29] ), .out0(new_n279));
  nano22aa1n03x5               g184(.a(new_n277), .b(new_n278), .c(new_n279), .out0(new_n280));
  oai012aa1n02x7               g185(.a(new_n276), .b(new_n272), .c(new_n269), .o1(new_n281));
  tech160nm_fiaoi012aa1n02p5x5 g186(.a(new_n279), .b(new_n281), .c(new_n278), .o1(new_n282));
  norp02aa1n03x5               g187(.a(new_n282), .b(new_n280), .o1(\s[29] ));
  xorb03aa1n02x5               g188(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g189(.a(new_n262), .b(new_n279), .c(new_n267), .out0(new_n285));
  aobi12aa1n02x7               g190(.a(new_n285), .b(new_n261), .c(new_n259), .out0(new_n286));
  oao003aa1n02x5               g191(.a(\a[29] ), .b(\b[28] ), .c(new_n278), .carry(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[29] ), .b(\a[30] ), .out0(new_n288));
  nano22aa1n03x5               g193(.a(new_n286), .b(new_n287), .c(new_n288), .out0(new_n289));
  oaih12aa1n02x5               g194(.a(new_n285), .b(new_n272), .c(new_n269), .o1(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n288), .b(new_n290), .c(new_n287), .o1(new_n291));
  norp02aa1n03x5               g196(.a(new_n291), .b(new_n289), .o1(\s[30] ));
  norb02aa1n02x5               g197(.a(new_n285), .b(new_n288), .out0(new_n293));
  aobi12aa1n02x7               g198(.a(new_n293), .b(new_n261), .c(new_n259), .out0(new_n294));
  oao003aa1n02x5               g199(.a(\a[30] ), .b(\b[29] ), .c(new_n287), .carry(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[30] ), .b(\a[31] ), .out0(new_n296));
  nano22aa1n03x5               g201(.a(new_n294), .b(new_n295), .c(new_n296), .out0(new_n297));
  oai012aa1n02x5               g202(.a(new_n293), .b(new_n272), .c(new_n269), .o1(new_n298));
  aoi012aa1n03x5               g203(.a(new_n296), .b(new_n298), .c(new_n295), .o1(new_n299));
  norp02aa1n03x5               g204(.a(new_n299), .b(new_n297), .o1(\s[31] ));
  xnbna2aa1n03x5               g205(.a(new_n121), .b(new_n115), .c(new_n116), .out0(\s[3] ));
  oaoi03aa1n02x5               g206(.a(\a[3] ), .b(\b[2] ), .c(new_n121), .o1(new_n302));
  xorb03aa1n02x5               g207(.a(new_n302), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g208(.a(new_n122), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g209(.a(new_n107), .b(new_n122), .c(new_n108), .o1(new_n305));
  xnrb03aa1n02x5               g210(.a(new_n305), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g211(.a(new_n109), .o1(new_n307));
  aobi12aa1n02x5               g212(.a(new_n125), .b(new_n122), .c(new_n307), .out0(new_n308));
  xnrb03aa1n02x5               g213(.a(new_n308), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g214(.a(\a[7] ), .b(\b[6] ), .c(new_n308), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  aoi112aa1n02x5               g216(.a(new_n126), .b(new_n127), .c(new_n122), .d(new_n110), .o1(new_n312));
  norb02aa1n02x5               g217(.a(new_n128), .b(new_n312), .out0(\s[9] ));
endmodule


