// Benchmark "adder" written by ABC on Thu Jul 18 08:57:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n128, new_n129, new_n130, new_n131, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n287, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n307, new_n309, new_n311,
    new_n313, new_n315, new_n317;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nand42aa1n02x5               g003(.a(\b[8] ), .b(\a[9] ), .o1(new_n99));
  nor002aa1n03x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nand42aa1n08x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nand42aa1n06x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nano23aa1n09x5               g008(.a(new_n100), .b(new_n102), .c(new_n103), .d(new_n101), .out0(new_n104));
  nor042aa1n02x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nanp02aa1n12x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor042aa1n03x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  ao0012aa1n03x7               g012(.a(new_n105), .b(new_n107), .c(new_n106), .o(new_n108));
  ao0012aa1n03x5               g013(.a(new_n100), .b(new_n102), .c(new_n101), .o(new_n109));
  aoi012aa1n12x5               g014(.a(new_n109), .b(new_n104), .c(new_n108), .o1(new_n110));
  xorc02aa1n12x5               g015(.a(\a[4] ), .b(\b[3] ), .out0(new_n111));
  nor002aa1n03x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanp02aa1n12x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  norb02aa1n03x5               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  nor042aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  aoi022aa1n06x5               g020(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n116));
  oai112aa1n06x5               g021(.a(new_n111), .b(new_n114), .c(new_n115), .d(new_n116), .o1(new_n117));
  aoi112aa1n02x7               g022(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n118));
  oab012aa1n04x5               g023(.a(new_n118), .b(\a[4] ), .c(\b[3] ), .out0(new_n119));
  nand42aa1n03x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nano23aa1n03x5               g025(.a(new_n105), .b(new_n107), .c(new_n120), .d(new_n106), .out0(new_n121));
  nanp02aa1n03x5               g026(.a(new_n121), .b(new_n104), .o1(new_n122));
  aoai13aa1n12x5               g027(.a(new_n110), .b(new_n122), .c(new_n117), .d(new_n119), .o1(new_n123));
  tech160nm_fiaoi012aa1n05x5   g028(.a(new_n98), .b(new_n123), .c(new_n99), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  oaoi03aa1n09x5               g030(.a(\a[10] ), .b(\b[9] ), .c(new_n124), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n02x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  nor042aa1n02x5               g035(.a(\b[11] ), .b(\a[12] ), .o1(new_n131));
  nand42aa1n02x5               g036(.a(\b[11] ), .b(\a[12] ), .o1(new_n132));
  nanb02aa1n02x5               g037(.a(new_n131), .b(new_n132), .out0(new_n133));
  aoai13aa1n03x5               g038(.a(new_n133), .b(new_n128), .c(new_n126), .d(new_n130), .o1(new_n134));
  nand22aa1n03x5               g039(.a(new_n126), .b(new_n130), .o1(new_n135));
  nona22aa1n02x4               g040(.a(new_n135), .b(new_n133), .c(new_n128), .out0(new_n136));
  nanp02aa1n03x5               g041(.a(new_n136), .b(new_n134), .o1(\s[12] ));
  nano23aa1n06x5               g042(.a(new_n128), .b(new_n131), .c(new_n132), .d(new_n129), .out0(new_n138));
  orn002aa1n02x5               g043(.a(\a[9] ), .b(\b[8] ), .o(new_n139));
  oaoi03aa1n02x5               g044(.a(\a[10] ), .b(\b[9] ), .c(new_n139), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n131), .b(new_n128), .c(new_n132), .o1(new_n141));
  aobi12aa1n06x5               g046(.a(new_n141), .b(new_n138), .c(new_n140), .out0(new_n142));
  xorc02aa1n02x5               g047(.a(\a[10] ), .b(\b[9] ), .out0(new_n143));
  norb02aa1n02x5               g048(.a(new_n99), .b(new_n98), .out0(new_n144));
  nanp03aa1n02x5               g049(.a(new_n138), .b(new_n143), .c(new_n144), .o1(new_n145));
  nanb02aa1n06x5               g050(.a(new_n145), .b(new_n123), .out0(new_n146));
  nand22aa1n03x5               g051(.a(new_n146), .b(new_n142), .o1(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nand02aa1n08x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  tech160nm_fiaoi012aa1n05x5   g055(.a(new_n149), .b(new_n147), .c(new_n150), .o1(new_n151));
  xnrb03aa1n03x5               g056(.a(new_n151), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nand42aa1n04x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nano23aa1d15x5               g059(.a(new_n149), .b(new_n153), .c(new_n154), .d(new_n150), .out0(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n153), .b(new_n149), .c(new_n154), .o1(new_n157));
  aoai13aa1n04x5               g062(.a(new_n157), .b(new_n156), .c(new_n146), .d(new_n142), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  nor022aa1n04x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nand42aa1n02x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  aoai13aa1n03x5               g070(.a(new_n165), .b(new_n160), .c(new_n158), .d(new_n162), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(new_n158), .b(new_n162), .o1(new_n167));
  nona22aa1n02x4               g072(.a(new_n167), .b(new_n165), .c(new_n160), .out0(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n166), .o1(\s[16] ));
  nano23aa1n06x5               g074(.a(new_n160), .b(new_n163), .c(new_n164), .d(new_n161), .out0(new_n170));
  oa0012aa1n02x5               g075(.a(new_n154), .b(new_n153), .c(new_n149), .o(new_n171));
  tech160nm_fiao0012aa1n02p5x5 g076(.a(new_n163), .b(new_n160), .c(new_n164), .o(new_n172));
  tech160nm_fiaoi012aa1n04x5   g077(.a(new_n172), .b(new_n170), .c(new_n171), .o1(new_n173));
  inv000aa1n02x5               g078(.a(new_n173), .o1(new_n174));
  nand22aa1n06x5               g079(.a(new_n170), .b(new_n155), .o1(new_n175));
  oab012aa1n12x5               g080(.a(new_n174), .b(new_n142), .c(new_n175), .out0(new_n176));
  nano32aa1d12x5               g081(.a(new_n175), .b(new_n138), .c(new_n144), .d(new_n143), .out0(new_n177));
  nand42aa1n10x5               g082(.a(new_n123), .b(new_n177), .o1(new_n178));
  nanp02aa1n06x5               g083(.a(new_n178), .b(new_n176), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g085(.a(\a[18] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n03x5               g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  oai012aa1n06x5               g090(.a(new_n173), .b(new_n142), .c(new_n175), .o1(new_n186));
  xroi22aa1d04x5               g091(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n187));
  aoai13aa1n06x5               g092(.a(new_n187), .b(new_n186), .c(new_n123), .d(new_n177), .o1(new_n188));
  nor042aa1n02x5               g093(.a(\b[17] ), .b(\a[18] ), .o1(new_n189));
  aoi112aa1n09x5               g094(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n190));
  nor042aa1n04x5               g095(.a(new_n190), .b(new_n189), .o1(new_n191));
  norp02aa1n24x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nand42aa1n10x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  norb02aa1n06x5               g098(.a(new_n193), .b(new_n192), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n188), .c(new_n191), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n03p5x5 g101(.a(new_n188), .b(new_n191), .o1(new_n197));
  nor002aa1d32x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nand02aa1d28x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  norb02aa1d21x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n201), .b(new_n192), .c(new_n197), .d(new_n193), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(new_n197), .b(new_n194), .o1(new_n203));
  nona22aa1n03x5               g108(.a(new_n203), .b(new_n201), .c(new_n192), .out0(new_n204));
  nanp02aa1n02x5               g109(.a(new_n204), .b(new_n202), .o1(\s[20] ));
  nona23aa1n09x5               g110(.a(new_n199), .b(new_n193), .c(new_n192), .d(new_n198), .out0(new_n206));
  aoi012aa1n06x5               g111(.a(new_n198), .b(new_n192), .c(new_n199), .o1(new_n207));
  oai012aa1n12x5               g112(.a(new_n207), .b(new_n206), .c(new_n191), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n206), .b(new_n187), .out0(new_n210));
  aoai13aa1n06x5               g115(.a(new_n209), .b(new_n210), .c(new_n178), .d(new_n176), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n08x5               g117(.a(\b[20] ), .b(\a[21] ), .o1(new_n213));
  xorc02aa1n12x5               g118(.a(\a[21] ), .b(\b[20] ), .out0(new_n214));
  tech160nm_fixnrc02aa1n05x5   g119(.a(\b[21] ), .b(\a[22] ), .out0(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n213), .c(new_n211), .d(new_n214), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(new_n211), .b(new_n214), .o1(new_n217));
  nona22aa1n02x4               g122(.a(new_n217), .b(new_n215), .c(new_n213), .out0(new_n218));
  nanp02aa1n03x5               g123(.a(new_n218), .b(new_n216), .o1(\s[22] ));
  oai112aa1n06x5               g124(.a(new_n194), .b(new_n200), .c(new_n190), .d(new_n189), .o1(new_n220));
  nanb02aa1n12x5               g125(.a(new_n215), .b(new_n214), .out0(new_n221));
  inv000aa1d42x5               g126(.a(\a[22] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\b[21] ), .o1(new_n223));
  oaoi03aa1n12x5               g128(.a(new_n222), .b(new_n223), .c(new_n213), .o1(new_n224));
  aoai13aa1n12x5               g129(.a(new_n224), .b(new_n221), .c(new_n220), .d(new_n207), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  nona23aa1n09x5               g131(.a(new_n187), .b(new_n214), .c(new_n215), .d(new_n206), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n226), .b(new_n227), .c(new_n178), .d(new_n176), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g134(.a(\b[22] ), .b(\a[23] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[23] ), .b(\b[22] ), .out0(new_n231));
  xorc02aa1n12x5               g136(.a(\a[24] ), .b(\b[23] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n03x5               g138(.a(new_n233), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(new_n228), .b(new_n231), .o1(new_n235));
  nona22aa1n02x4               g140(.a(new_n235), .b(new_n233), .c(new_n230), .out0(new_n236));
  nanp02aa1n03x5               g141(.a(new_n236), .b(new_n234), .o1(\s[24] ));
  norb02aa1n02x5               g142(.a(new_n214), .b(new_n215), .out0(new_n238));
  and002aa1n02x5               g143(.a(new_n232), .b(new_n231), .o(new_n239));
  nano22aa1n03x5               g144(.a(new_n210), .b(new_n239), .c(new_n238), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n186), .c(new_n123), .d(new_n177), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n224), .o1(new_n242));
  aoai13aa1n06x5               g147(.a(new_n239), .b(new_n242), .c(new_n208), .d(new_n238), .o1(new_n243));
  inv000aa1d42x5               g148(.a(\a[24] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(\b[23] ), .o1(new_n245));
  oaoi03aa1n12x5               g150(.a(new_n244), .b(new_n245), .c(new_n230), .o1(new_n246));
  nanp02aa1n03x5               g151(.a(new_n243), .b(new_n246), .o1(new_n247));
  nanb02aa1n03x5               g152(.a(new_n247), .b(new_n241), .out0(new_n248));
  xorb03aa1n02x5               g153(.a(new_n248), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g154(.a(\b[24] ), .b(\a[25] ), .o1(new_n250));
  tech160nm_fixorc02aa1n02p5x5 g155(.a(\a[25] ), .b(\b[24] ), .out0(new_n251));
  xorc02aa1n12x5               g156(.a(\a[26] ), .b(\b[25] ), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n250), .c(new_n248), .d(new_n251), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n251), .b(new_n247), .c(new_n179), .d(new_n240), .o1(new_n255));
  nona22aa1n02x5               g160(.a(new_n255), .b(new_n253), .c(new_n250), .out0(new_n256));
  nanp02aa1n03x5               g161(.a(new_n254), .b(new_n256), .o1(\s[26] ));
  inv000aa1d42x5               g162(.a(new_n246), .o1(new_n258));
  and002aa1n18x5               g163(.a(new_n252), .b(new_n251), .o(new_n259));
  aoai13aa1n09x5               g164(.a(new_n259), .b(new_n258), .c(new_n225), .d(new_n239), .o1(new_n260));
  aoi112aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n261));
  oab012aa1n02x4               g166(.a(new_n261), .b(\a[26] ), .c(\b[25] ), .out0(new_n262));
  nano22aa1n03x7               g167(.a(new_n227), .b(new_n239), .c(new_n259), .out0(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n186), .c(new_n123), .d(new_n177), .o1(new_n264));
  nand23aa1n04x5               g169(.a(new_n264), .b(new_n260), .c(new_n262), .o1(new_n265));
  xorb03aa1n02x5               g170(.a(new_n265), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor002aa1n02x5               g171(.a(\b[26] ), .b(\a[27] ), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[27] ), .b(\b[26] ), .out0(new_n268));
  xnrc02aa1n02x5               g173(.a(\b[27] ), .b(\a[28] ), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n267), .c(new_n265), .d(new_n268), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n259), .o1(new_n271));
  aoai13aa1n04x5               g176(.a(new_n262), .b(new_n271), .c(new_n243), .d(new_n246), .o1(new_n272));
  aobi12aa1n09x5               g177(.a(new_n263), .b(new_n178), .c(new_n176), .out0(new_n273));
  oai012aa1n02x7               g178(.a(new_n268), .b(new_n272), .c(new_n273), .o1(new_n274));
  nona22aa1n02x5               g179(.a(new_n274), .b(new_n269), .c(new_n267), .out0(new_n275));
  nanp02aa1n03x5               g180(.a(new_n275), .b(new_n270), .o1(\s[28] ));
  norb02aa1n02x5               g181(.a(new_n268), .b(new_n269), .out0(new_n277));
  oai012aa1n03x5               g182(.a(new_n277), .b(new_n272), .c(new_n273), .o1(new_n278));
  aob012aa1n02x5               g183(.a(new_n267), .b(\b[27] ), .c(\a[28] ), .out0(new_n279));
  tech160nm_fioai012aa1n03p5x5 g184(.a(new_n279), .b(\b[27] ), .c(\a[28] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(\b[28] ), .b(\a[29] ), .o1(new_n281));
  and002aa1n02x5               g186(.a(\b[28] ), .b(\a[29] ), .o(new_n282));
  nona32aa1n03x5               g187(.a(new_n278), .b(new_n282), .c(new_n281), .d(new_n280), .out0(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[28] ), .b(\a[29] ), .out0(new_n284));
  aoai13aa1n02x7               g189(.a(new_n284), .b(new_n280), .c(new_n265), .d(new_n277), .o1(new_n285));
  nanp02aa1n03x5               g190(.a(new_n285), .b(new_n283), .o1(\s[29] ));
  nanp02aa1n02x5               g191(.a(\b[0] ), .b(\a[1] ), .o1(new_n287));
  xorb03aa1n02x5               g192(.a(new_n287), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g193(.a(new_n268), .b(new_n284), .c(new_n269), .out0(new_n289));
  inv000aa1d42x5               g194(.a(new_n282), .o1(new_n290));
  tech160nm_fiao0012aa1n02p5x5 g195(.a(new_n281), .b(new_n280), .c(new_n290), .o(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[29] ), .b(\a[30] ), .out0(new_n292));
  aoai13aa1n02x7               g197(.a(new_n292), .b(new_n291), .c(new_n265), .d(new_n289), .o1(new_n293));
  oaih12aa1n02x5               g198(.a(new_n289), .b(new_n272), .c(new_n273), .o1(new_n294));
  norp02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .o1(new_n295));
  and002aa1n02x5               g200(.a(\b[29] ), .b(\a[30] ), .o(new_n296));
  nona32aa1n02x5               g201(.a(new_n294), .b(new_n296), .c(new_n295), .d(new_n291), .out0(new_n297));
  nanp02aa1n03x5               g202(.a(new_n293), .b(new_n297), .o1(\s[30] ));
  norb02aa1n02x5               g203(.a(new_n291), .b(new_n292), .out0(new_n299));
  norb02aa1n02x5               g204(.a(new_n289), .b(new_n292), .out0(new_n300));
  oaih12aa1n02x5               g205(.a(new_n300), .b(new_n272), .c(new_n273), .o1(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[30] ), .b(\a[31] ), .out0(new_n302));
  nona32aa1n03x5               g207(.a(new_n301), .b(new_n302), .c(new_n299), .d(new_n295), .out0(new_n303));
  oabi12aa1n02x5               g208(.a(new_n299), .b(\a[30] ), .c(\b[29] ), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n302), .b(new_n304), .c(new_n265), .d(new_n300), .o1(new_n305));
  nanp02aa1n03x5               g210(.a(new_n305), .b(new_n303), .o1(\s[31] ));
  norp02aa1n02x5               g211(.a(new_n116), .b(new_n115), .o1(new_n307));
  xnrb03aa1n02x5               g212(.a(new_n307), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi13aa1n02x5               g213(.a(new_n112), .b(new_n113), .c(new_n116), .d(new_n115), .o1(new_n309));
  xnrc02aa1n02x5               g214(.a(new_n309), .b(new_n111), .out0(\s[4] ));
  nanp02aa1n02x5               g215(.a(new_n117), .b(new_n119), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g217(.a(new_n107), .b(new_n311), .c(new_n120), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g219(.a(new_n108), .b(new_n311), .c(new_n121), .o(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g221(.a(new_n102), .b(new_n315), .c(new_n103), .o1(new_n317));
  xnrb03aa1n02x5               g222(.a(new_n317), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g223(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


