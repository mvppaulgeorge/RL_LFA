// Benchmark "adder" written by ABC on Wed Jul 17 20:36:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n339, new_n340, new_n342, new_n343, new_n344, new_n346, new_n347,
    new_n349, new_n350, new_n351, new_n352, new_n354, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[4] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[3] ), .o1(new_n99));
  nor042aa1n03x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  tech160nm_fiaoi012aa1n03p5x5 g005(.a(new_n100), .b(new_n98), .c(new_n99), .o1(new_n101));
  nand02aa1d12x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  norb02aa1n02x5               g007(.a(new_n102), .b(new_n100), .out0(new_n103));
  tech160nm_finand02aa1n03p5x5 g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nor042aa1n04x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand22aa1n12x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  oai112aa1n03x5               g011(.a(new_n103), .b(new_n104), .c(new_n105), .d(new_n106), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  aoi122aa1n06x5               g013(.a(new_n108), .b(\b[6] ), .c(\a[7] ), .d(\b[3] ), .e(\a[4] ), .o1(new_n109));
  nand42aa1d28x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  tech160nm_fioai012aa1n03p5x5 g015(.a(new_n110), .b(\b[6] ), .c(\a[7] ), .o1(new_n111));
  oai022aa1d18x5               g016(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n112));
  aoi022aa1n02x7               g017(.a(\b[7] ), .b(\a[8] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n109), .b(new_n113), .c(new_n112), .d(new_n111), .out0(new_n114));
  inv000aa1d42x5               g019(.a(\a[7] ), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\b[6] ), .o1(new_n116));
  nand02aa1n04x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  aoai13aa1n06x5               g022(.a(new_n117), .b(new_n108), .c(new_n115), .d(new_n116), .o1(new_n118));
  nand22aa1n03x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano22aa1n02x4               g024(.a(new_n108), .b(new_n119), .c(new_n117), .out0(new_n120));
  nor042aa1n04x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nor002aa1n16x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  oab012aa1n03x5               g027(.a(new_n111), .b(new_n121), .c(new_n122), .out0(new_n123));
  aobi12aa1n06x5               g028(.a(new_n118), .b(new_n123), .c(new_n120), .out0(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n114), .c(new_n101), .d(new_n107), .o1(new_n125));
  nanp02aa1n04x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  nor042aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand22aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n03x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  aoai13aa1n06x5               g034(.a(new_n129), .b(new_n97), .c(new_n125), .d(new_n126), .o1(new_n130));
  norb02aa1n03x5               g035(.a(new_n126), .b(new_n97), .out0(new_n131));
  aoi112aa1n02x5               g036(.a(new_n129), .b(new_n97), .c(new_n125), .d(new_n131), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n130), .b(new_n132), .out0(\s[10] ));
  inv040aa1n08x5               g038(.a(new_n97), .o1(new_n134));
  oaoi03aa1n12x5               g039(.a(\a[10] ), .b(\b[9] ), .c(new_n134), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nor042aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand02aa1n06x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n130), .c(new_n136), .out0(\s[11] ));
  aobi12aa1n06x5               g045(.a(new_n139), .b(new_n130), .c(new_n136), .out0(new_n141));
  nor042aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1n08x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  inv020aa1n02x5               g048(.a(new_n143), .o1(new_n144));
  oai022aa1n03x5               g049(.a(new_n141), .b(new_n137), .c(new_n144), .d(new_n142), .o1(new_n145));
  norb03aa1n02x5               g050(.a(new_n143), .b(new_n137), .c(new_n142), .out0(new_n146));
  oaib12aa1n03x5               g051(.a(new_n145), .b(new_n141), .c(new_n146), .out0(\s[12] ));
  inv000aa1d42x5               g052(.a(\b[2] ), .o1(new_n148));
  nanb02aa1n03x5               g053(.a(\a[3] ), .b(new_n148), .out0(new_n149));
  nanp02aa1n02x5               g054(.a(new_n149), .b(new_n102), .o1(new_n150));
  tech160nm_fioai012aa1n04x5   g055(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n151));
  tech160nm_fioai012aa1n05x5   g056(.a(new_n101), .b(new_n151), .c(new_n150), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n108), .o1(new_n153));
  aoi022aa1n02x5               g058(.a(\b[6] ), .b(\a[7] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n154));
  nor022aa1n16x5               g059(.a(\b[6] ), .b(\a[7] ), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n155), .b(\a[6] ), .c(\b[5] ), .o1(new_n156));
  nona22aa1n02x4               g061(.a(new_n113), .b(new_n122), .c(new_n121), .out0(new_n157));
  nano32aa1n03x7               g062(.a(new_n157), .b(new_n156), .c(new_n154), .d(new_n153), .out0(new_n158));
  nanb03aa1n03x5               g063(.a(new_n108), .b(new_n117), .c(new_n119), .out0(new_n159));
  oai112aa1n02x5               g064(.a(new_n112), .b(new_n110), .c(\b[6] ), .d(\a[7] ), .o1(new_n160));
  oai012aa1n06x5               g065(.a(new_n118), .b(new_n160), .c(new_n159), .o1(new_n161));
  nona23aa1n03x5               g066(.a(new_n143), .b(new_n138), .c(new_n137), .d(new_n142), .out0(new_n162));
  nano22aa1n03x7               g067(.a(new_n162), .b(new_n131), .c(new_n129), .out0(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n161), .c(new_n158), .d(new_n152), .o1(new_n164));
  nanb03aa1n03x5               g069(.a(new_n142), .b(new_n143), .c(new_n138), .out0(new_n165));
  oai122aa1n02x7               g070(.a(new_n128), .b(new_n127), .c(new_n97), .d(\b[10] ), .e(\a[11] ), .o1(new_n166));
  oaih12aa1n06x5               g071(.a(new_n143), .b(new_n142), .c(new_n137), .o1(new_n167));
  tech160nm_fioai012aa1n04x5   g072(.a(new_n167), .b(new_n166), .c(new_n165), .o1(new_n168));
  nanb02aa1n02x5               g073(.a(new_n168), .b(new_n164), .out0(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n16x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[12] ), .b(\a[13] ), .o1(new_n173));
  nanp03aa1n02x5               g078(.a(new_n169), .b(new_n172), .c(new_n173), .o1(new_n174));
  nor002aa1n04x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nand02aa1n06x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  oaih22aa1d12x5               g082(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n178));
  nanb03aa1n02x5               g083(.a(new_n178), .b(new_n174), .c(new_n176), .out0(new_n179));
  aoai13aa1n02x5               g084(.a(new_n179), .b(new_n177), .c(new_n172), .d(new_n174), .o1(\s[14] ));
  nano23aa1n06x5               g085(.a(new_n171), .b(new_n175), .c(new_n176), .d(new_n173), .out0(new_n181));
  aoai13aa1n03x5               g086(.a(new_n181), .b(new_n168), .c(new_n125), .d(new_n163), .o1(new_n182));
  oai012aa1n02x5               g087(.a(new_n176), .b(new_n175), .c(new_n171), .o1(new_n183));
  nor002aa1n06x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  nand42aa1n03x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nanb02aa1n06x5               g090(.a(new_n184), .b(new_n185), .out0(new_n186));
  xobna2aa1n03x5               g091(.a(new_n186), .b(new_n182), .c(new_n183), .out0(\s[15] ));
  aoi012aa1n02x7               g092(.a(new_n186), .b(new_n182), .c(new_n183), .o1(new_n188));
  inv040aa1d32x5               g093(.a(\a[16] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[15] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n190), .b(new_n189), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(\b[15] ), .b(\a[16] ), .o1(new_n192));
  nanp02aa1n03x5               g097(.a(new_n191), .b(new_n192), .o1(new_n193));
  oai012aa1n03x5               g098(.a(new_n193), .b(new_n188), .c(new_n184), .o1(new_n194));
  nano22aa1n02x4               g099(.a(new_n184), .b(new_n191), .c(new_n192), .out0(new_n195));
  oaib12aa1n03x5               g100(.a(new_n194), .b(new_n188), .c(new_n195), .out0(\s[16] ));
  aoi012aa1n06x5               g101(.a(new_n161), .b(new_n158), .c(new_n152), .o1(new_n197));
  nona23aa1n03x5               g102(.a(new_n176), .b(new_n173), .c(new_n171), .d(new_n175), .out0(new_n198));
  nor043aa1n03x5               g103(.a(new_n198), .b(new_n186), .c(new_n193), .o1(new_n199));
  nand02aa1n02x5               g104(.a(new_n199), .b(new_n163), .o1(new_n200));
  nanp03aa1n02x5               g105(.a(new_n191), .b(new_n185), .c(new_n192), .o1(new_n201));
  oai112aa1n02x5               g106(.a(new_n178), .b(new_n176), .c(\b[14] ), .d(\a[15] ), .o1(new_n202));
  oao003aa1n03x5               g107(.a(new_n189), .b(new_n190), .c(new_n184), .carry(new_n203));
  oabi12aa1n02x5               g108(.a(new_n203), .b(new_n201), .c(new_n202), .out0(new_n204));
  aoi012aa1n02x7               g109(.a(new_n204), .b(new_n168), .c(new_n199), .o1(new_n205));
  oai012aa1n09x5               g110(.a(new_n205), .b(new_n197), .c(new_n200), .o1(new_n206));
  xorb03aa1n02x5               g111(.a(new_n206), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  inv040aa1n08x5               g113(.a(new_n208), .o1(new_n209));
  nano23aa1n02x4               g114(.a(new_n137), .b(new_n142), .c(new_n143), .d(new_n138), .out0(new_n210));
  nona22aa1n03x5               g115(.a(new_n181), .b(new_n186), .c(new_n193), .out0(new_n211));
  nano32aa1n03x7               g116(.a(new_n211), .b(new_n210), .c(new_n129), .d(new_n131), .out0(new_n212));
  oai012aa1n02x5               g117(.a(new_n138), .b(\b[11] ), .c(\a[12] ), .o1(new_n213));
  nona32aa1n06x5               g118(.a(new_n135), .b(new_n213), .c(new_n144), .d(new_n137), .out0(new_n214));
  oab012aa1n02x4               g119(.a(new_n203), .b(new_n202), .c(new_n201), .out0(new_n215));
  aoai13aa1n04x5               g120(.a(new_n215), .b(new_n211), .c(new_n214), .d(new_n167), .o1(new_n216));
  xorc02aa1n12x5               g121(.a(\a[17] ), .b(\b[16] ), .out0(new_n217));
  aoai13aa1n02x5               g122(.a(new_n217), .b(new_n216), .c(new_n125), .d(new_n212), .o1(new_n218));
  xorc02aa1n12x5               g123(.a(\a[18] ), .b(\b[17] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(\a[18] ), .o1(new_n220));
  inv000aa1d42x5               g125(.a(\b[17] ), .o1(new_n221));
  aoi012aa1n02x5               g126(.a(new_n208), .b(new_n220), .c(new_n221), .o1(new_n222));
  oai112aa1n02x5               g127(.a(new_n218), .b(new_n222), .c(new_n221), .d(new_n220), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n223), .b(new_n219), .c(new_n209), .d(new_n218), .o1(\s[18] ));
  and002aa1n02x5               g129(.a(new_n219), .b(new_n217), .o(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n216), .c(new_n125), .d(new_n212), .o1(new_n226));
  oaoi03aa1n12x5               g131(.a(\a[18] ), .b(\b[17] ), .c(new_n209), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  nor002aa1n06x5               g133(.a(\b[18] ), .b(\a[19] ), .o1(new_n229));
  nanp02aa1n06x5               g134(.a(\b[18] ), .b(\a[19] ), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  xnbna2aa1n03x5               g136(.a(new_n231), .b(new_n226), .c(new_n228), .out0(\s[19] ));
  xnrc02aa1n02x5               g137(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aobi12aa1n06x5               g138(.a(new_n231), .b(new_n226), .c(new_n228), .out0(new_n234));
  xorc02aa1n02x5               g139(.a(\a[20] ), .b(\b[19] ), .out0(new_n235));
  oabi12aa1n03x5               g140(.a(new_n235), .b(new_n234), .c(new_n229), .out0(new_n236));
  inv040aa1d32x5               g141(.a(\a[20] ), .o1(new_n237));
  inv030aa1d32x5               g142(.a(\b[19] ), .o1(new_n238));
  nand02aa1n04x5               g143(.a(new_n238), .b(new_n237), .o1(new_n239));
  and002aa1n12x5               g144(.a(\b[19] ), .b(\a[20] ), .o(new_n240));
  norb03aa1n02x5               g145(.a(new_n239), .b(new_n229), .c(new_n240), .out0(new_n241));
  oaib12aa1n02x5               g146(.a(new_n236), .b(new_n234), .c(new_n241), .out0(\s[20] ));
  nano23aa1n06x5               g147(.a(new_n229), .b(new_n240), .c(new_n239), .d(new_n230), .out0(new_n243));
  nand23aa1d12x5               g148(.a(new_n243), .b(new_n217), .c(new_n219), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  oai012aa1n02x5               g150(.a(new_n230), .b(\b[19] ), .c(\a[20] ), .o1(new_n246));
  nona32aa1n06x5               g151(.a(new_n227), .b(new_n246), .c(new_n240), .d(new_n229), .out0(new_n247));
  oaoi03aa1n03x5               g152(.a(new_n237), .b(new_n238), .c(new_n229), .o1(new_n248));
  nanp02aa1n02x5               g153(.a(new_n247), .b(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[21] ), .b(\b[20] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(new_n206), .d(new_n245), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(new_n250), .b(new_n249), .c(new_n206), .d(new_n245), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(\s[21] ));
  norp02aa1n02x5               g158(.a(\b[20] ), .b(\a[21] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  xorc02aa1n02x5               g160(.a(\a[22] ), .b(\b[21] ), .out0(new_n256));
  nanp02aa1n02x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  oai022aa1n02x5               g162(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n258));
  nanb03aa1n03x5               g163(.a(new_n258), .b(new_n251), .c(new_n257), .out0(new_n259));
  aoai13aa1n02x5               g164(.a(new_n259), .b(new_n256), .c(new_n251), .d(new_n255), .o1(\s[22] ));
  nanp02aa1n02x5               g165(.a(new_n256), .b(new_n250), .o1(new_n261));
  nano32aa1n02x4               g166(.a(new_n261), .b(new_n243), .c(new_n219), .d(new_n217), .out0(new_n262));
  nanp02aa1n02x5               g167(.a(new_n258), .b(new_n257), .o1(new_n263));
  aoai13aa1n12x5               g168(.a(new_n263), .b(new_n261), .c(new_n247), .d(new_n248), .o1(new_n264));
  xorc02aa1n02x5               g169(.a(\a[23] ), .b(\b[22] ), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n264), .c(new_n206), .d(new_n262), .o1(new_n266));
  aoi112aa1n02x5               g171(.a(new_n265), .b(new_n264), .c(new_n206), .d(new_n262), .o1(new_n267));
  norb02aa1n02x5               g172(.a(new_n266), .b(new_n267), .out0(\s[23] ));
  nor042aa1n06x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[24] ), .b(\b[23] ), .out0(new_n271));
  nand42aa1n03x5               g176(.a(\b[23] ), .b(\a[24] ), .o1(new_n272));
  oab012aa1n02x4               g177(.a(new_n269), .b(\a[24] ), .c(\b[23] ), .out0(new_n273));
  nanp03aa1n03x5               g178(.a(new_n266), .b(new_n272), .c(new_n273), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n271), .c(new_n270), .d(new_n266), .o1(\s[24] ));
  nand42aa1n03x5               g180(.a(\b[22] ), .b(\a[23] ), .o1(new_n276));
  norp02aa1n02x5               g181(.a(\b[23] ), .b(\a[24] ), .o1(new_n277));
  nano23aa1n06x5               g182(.a(new_n269), .b(new_n277), .c(new_n272), .d(new_n276), .out0(new_n278));
  nano32aa1n02x5               g183(.a(new_n244), .b(new_n278), .c(new_n250), .d(new_n256), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n216), .c(new_n125), .d(new_n212), .o1(new_n280));
  oaoi03aa1n02x5               g185(.a(\a[24] ), .b(\b[23] ), .c(new_n270), .o1(new_n281));
  aoi012aa1n02x7               g186(.a(new_n281), .b(new_n264), .c(new_n278), .o1(new_n282));
  xorc02aa1n12x5               g187(.a(\a[25] ), .b(\b[24] ), .out0(new_n283));
  xnbna2aa1n03x5               g188(.a(new_n283), .b(new_n280), .c(new_n282), .out0(\s[25] ));
  norp02aa1n02x5               g189(.a(\b[24] ), .b(\a[25] ), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  aob012aa1n03x5               g191(.a(new_n283), .b(new_n280), .c(new_n282), .out0(new_n287));
  xorc02aa1n02x5               g192(.a(\a[26] ), .b(\b[25] ), .out0(new_n288));
  nanp02aa1n02x5               g193(.a(\b[25] ), .b(\a[26] ), .o1(new_n289));
  oai022aa1n02x5               g194(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n290));
  norb02aa1n02x5               g195(.a(new_n289), .b(new_n290), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n287), .b(new_n291), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n288), .c(new_n286), .d(new_n287), .o1(\s[26] ));
  and002aa1n02x5               g198(.a(new_n288), .b(new_n283), .o(new_n294));
  aoai13aa1n09x5               g199(.a(new_n294), .b(new_n281), .c(new_n264), .d(new_n278), .o1(new_n295));
  nand03aa1n02x5               g200(.a(new_n278), .b(new_n250), .c(new_n256), .o1(new_n296));
  norb03aa1n06x5               g201(.a(new_n294), .b(new_n244), .c(new_n296), .out0(new_n297));
  aoai13aa1n04x5               g202(.a(new_n297), .b(new_n216), .c(new_n125), .d(new_n212), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n290), .b(new_n289), .o1(new_n299));
  nanp03aa1d12x5               g204(.a(new_n295), .b(new_n298), .c(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  aoi122aa1n02x5               g206(.a(new_n301), .b(new_n289), .c(new_n290), .d(new_n206), .e(new_n297), .o1(new_n302));
  aoi022aa1n02x5               g207(.a(new_n302), .b(new_n295), .c(new_n300), .d(new_n301), .o1(\s[27] ));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  norp02aa1n02x5               g209(.a(\b[27] ), .b(\a[28] ), .o1(new_n305));
  nanp02aa1n02x5               g210(.a(\b[27] ), .b(\a[28] ), .o1(new_n306));
  nanb02aa1n02x5               g211(.a(new_n305), .b(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n304), .c(new_n300), .d(new_n301), .o1(new_n308));
  aoi022aa1n06x5               g213(.a(new_n206), .b(new_n297), .c(new_n289), .d(new_n290), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n301), .o1(new_n310));
  norb03aa1n02x5               g215(.a(new_n306), .b(new_n304), .c(new_n305), .out0(new_n311));
  aoai13aa1n02x5               g216(.a(new_n311), .b(new_n310), .c(new_n309), .d(new_n295), .o1(new_n312));
  nanp02aa1n03x5               g217(.a(new_n308), .b(new_n312), .o1(\s[28] ));
  norb02aa1n03x5               g218(.a(new_n301), .b(new_n307), .out0(new_n314));
  nand02aa1n02x5               g219(.a(new_n300), .b(new_n314), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n314), .o1(new_n316));
  aoi012aa1n02x5               g221(.a(new_n305), .b(new_n304), .c(new_n306), .o1(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n316), .c(new_n309), .d(new_n295), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[29] ), .b(\b[28] ), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n317), .b(new_n319), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n315), .d(new_n320), .o1(\s[29] ));
  xorb03aa1n02x5               g226(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g227(.a(new_n307), .b(new_n301), .c(new_n319), .out0(new_n323));
  nand02aa1n02x5               g228(.a(new_n300), .b(new_n323), .o1(new_n324));
  inv000aa1n02x5               g229(.a(new_n323), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .c(new_n317), .carry(new_n326));
  aoai13aa1n02x7               g231(.a(new_n326), .b(new_n325), .c(new_n309), .d(new_n295), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .out0(new_n328));
  norb02aa1n02x5               g233(.a(new_n326), .b(new_n328), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n324), .d(new_n329), .o1(\s[30] ));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  nand03aa1n02x5               g236(.a(new_n314), .b(new_n319), .c(new_n328), .o1(new_n332));
  nanb02aa1n03x5               g237(.a(new_n332), .b(new_n300), .out0(new_n333));
  oao003aa1n02x5               g238(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n334));
  aoai13aa1n02x7               g239(.a(new_n334), .b(new_n332), .c(new_n309), .d(new_n295), .o1(new_n335));
  norb02aa1n02x5               g240(.a(new_n334), .b(new_n331), .out0(new_n336));
  aoi022aa1n03x5               g241(.a(new_n335), .b(new_n331), .c(new_n333), .d(new_n336), .o1(\s[31] ));
  xnbna2aa1n03x5               g242(.a(new_n151), .b(new_n149), .c(new_n102), .out0(\s[3] ));
  xorc02aa1n02x5               g243(.a(\a[4] ), .b(\b[3] ), .out0(new_n339));
  norp02aa1n02x5               g244(.a(new_n339), .b(new_n100), .o1(new_n340));
  aoi022aa1n02x5               g245(.a(new_n152), .b(new_n339), .c(new_n340), .d(new_n107), .o1(\s[4] ));
  xorc02aa1n02x5               g246(.a(\a[5] ), .b(\b[4] ), .out0(new_n342));
  oaoi13aa1n02x5               g247(.a(new_n342), .b(new_n152), .c(new_n98), .d(new_n99), .o1(new_n343));
  oai112aa1n03x5               g248(.a(new_n152), .b(new_n342), .c(new_n99), .d(new_n98), .o1(new_n344));
  norb02aa1n02x5               g249(.a(new_n344), .b(new_n343), .out0(\s[5] ));
  inv000aa1d42x5               g250(.a(new_n122), .o1(new_n346));
  norb02aa1n02x5               g251(.a(new_n110), .b(new_n121), .out0(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n347), .b(new_n344), .c(new_n346), .out0(\s[6] ));
  nanp02aa1n03x5               g253(.a(new_n344), .b(new_n346), .o1(new_n349));
  norb02aa1n02x5               g254(.a(new_n119), .b(new_n155), .out0(new_n350));
  aoai13aa1n06x5               g255(.a(new_n350), .b(new_n121), .c(new_n349), .d(new_n110), .o1(new_n351));
  aoi112aa1n02x5               g256(.a(new_n350), .b(new_n121), .c(new_n349), .d(new_n347), .o1(new_n352));
  norb02aa1n02x5               g257(.a(new_n351), .b(new_n352), .out0(\s[7] ));
  inv000aa1d42x5               g258(.a(new_n155), .o1(new_n354));
  norb02aa1n02x5               g259(.a(new_n117), .b(new_n108), .out0(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n355), .b(new_n351), .c(new_n354), .out0(\s[8] ));
  xnbna2aa1n03x5               g261(.a(new_n197), .b(new_n126), .c(new_n134), .out0(\s[9] ));
endmodule


