// Benchmark "adder" written by ABC on Thu Jul 18 02:33:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n331, new_n333, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixnrc02aa1n02p5x5 g001(.a(\b[7] ), .b(\a[8] ), .out0(new_n97));
  nor002aa1d24x5               g002(.a(\b[6] ), .b(\a[7] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nanb02aa1n02x5               g004(.a(new_n98), .b(new_n99), .out0(new_n100));
  nanp02aa1n02x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  nor022aa1n08x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  tech160nm_finor002aa1n05x5   g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  oai012aa1n02x5               g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  inv000aa1d42x5               g009(.a(new_n98), .o1(new_n105));
  oao003aa1n02x5               g010(.a(\a[8] ), .b(\b[7] ), .c(new_n105), .carry(new_n106));
  oai013aa1n03x5               g011(.a(new_n106), .b(new_n97), .c(new_n104), .d(new_n100), .o1(new_n107));
  nor022aa1n06x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor002aa1n06x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  aoi012aa1n02x5               g015(.a(new_n108), .b(new_n109), .c(new_n110), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[1] ), .b(\a[2] ), .o1(new_n112));
  nand02aa1d04x5               g017(.a(\b[0] ), .b(\a[1] ), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  tech160nm_fioai012aa1n04x5   g019(.a(new_n112), .b(new_n114), .c(new_n113), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nona23aa1n03x5               g021(.a(new_n110), .b(new_n116), .c(new_n109), .d(new_n108), .out0(new_n117));
  oai012aa1n09x5               g022(.a(new_n111), .b(new_n117), .c(new_n115), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(new_n102), .b(new_n101), .out0(new_n119));
  nanp02aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nona23aa1n02x4               g025(.a(new_n120), .b(new_n99), .c(new_n98), .d(new_n103), .out0(new_n121));
  nor043aa1n03x5               g026(.a(new_n121), .b(new_n119), .c(new_n97), .o1(new_n122));
  aoi012aa1n06x5               g027(.a(new_n107), .b(new_n118), .c(new_n122), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .c(new_n123), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1d28x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  oaih22aa1d12x5               g031(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  nor042aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanb02aa1n02x5               g033(.a(new_n128), .b(new_n126), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  nor002aa1n04x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nand42aa1n08x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  nano22aa1n03x7               g038(.a(new_n123), .b(new_n130), .c(new_n133), .out0(new_n134));
  inv040aa1d32x5               g039(.a(\a[11] ), .o1(new_n135));
  inv040aa1d32x5               g040(.a(\b[10] ), .o1(new_n136));
  nand02aa1d08x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  nand22aa1n12x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand22aa1n12x5               g043(.a(new_n137), .b(new_n138), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  aoai13aa1n06x5               g045(.a(new_n140), .b(new_n134), .c(new_n126), .d(new_n127), .o1(new_n141));
  aoi112aa1n02x5               g046(.a(new_n134), .b(new_n140), .c(new_n126), .d(new_n127), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(\s[11] ));
  inv040aa1d32x5               g048(.a(\a[12] ), .o1(new_n144));
  inv040aa1d32x5               g049(.a(\b[11] ), .o1(new_n145));
  nand02aa1n03x5               g050(.a(new_n145), .b(new_n144), .o1(new_n146));
  nand22aa1n03x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1d04x5               g052(.a(new_n146), .b(new_n147), .o1(new_n148));
  xobna2aa1n03x5               g053(.a(new_n148), .b(new_n141), .c(new_n137), .out0(\s[12] ));
  nano23aa1d15x5               g054(.a(new_n128), .b(new_n131), .c(new_n132), .d(new_n126), .out0(new_n150));
  nona22aa1d30x5               g055(.a(new_n150), .b(new_n148), .c(new_n139), .out0(new_n151));
  nor002aa1n04x5               g056(.a(\b[10] ), .b(\a[11] ), .o1(new_n152));
  nanb03aa1n06x5               g057(.a(new_n152), .b(new_n138), .c(new_n126), .out0(new_n153));
  nand23aa1n03x5               g058(.a(new_n127), .b(new_n146), .c(new_n147), .o1(new_n154));
  oaoi03aa1n02x5               g059(.a(new_n144), .b(new_n145), .c(new_n152), .o1(new_n155));
  oai012aa1n02x7               g060(.a(new_n155), .b(new_n154), .c(new_n153), .o1(new_n156));
  oabi12aa1n06x5               g061(.a(new_n156), .b(new_n123), .c(new_n151), .out0(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n02x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand22aa1n03x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n03x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand42aa1n03x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1n06x5               g069(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n165));
  oa0012aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n159), .o(new_n166));
  aoi012aa1n02x5               g071(.a(new_n166), .b(new_n156), .c(new_n165), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n151), .o1(new_n168));
  nano22aa1n03x7               g073(.a(new_n123), .b(new_n168), .c(new_n165), .out0(new_n169));
  nor042aa1n09x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand42aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  oaib12aa1n06x5               g077(.a(new_n172), .b(new_n169), .c(new_n167), .out0(new_n173));
  norb03aa1n02x5               g078(.a(new_n167), .b(new_n169), .c(new_n172), .out0(new_n174));
  norb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(\s[15] ));
  inv000aa1d42x5               g080(.a(new_n170), .o1(new_n176));
  nor042aa1n03x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand42aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n173), .c(new_n176), .out0(\s[16] ));
  nano23aa1n09x5               g085(.a(new_n170), .b(new_n177), .c(new_n178), .d(new_n171), .out0(new_n181));
  nano22aa1d15x5               g086(.a(new_n151), .b(new_n165), .c(new_n181), .out0(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n107), .c(new_n118), .d(new_n122), .o1(new_n183));
  aoai13aa1n02x7               g088(.a(new_n181), .b(new_n166), .c(new_n156), .d(new_n165), .o1(new_n184));
  aoi012aa1d18x5               g089(.a(new_n177), .b(new_n170), .c(new_n178), .o1(new_n185));
  nand23aa1n06x5               g090(.a(new_n183), .b(new_n184), .c(new_n185), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g092(.a(\a[18] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\a[17] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[16] ), .o1(new_n190));
  oaoi03aa1n03x5               g095(.a(new_n189), .b(new_n190), .c(new_n186), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[17] ), .c(new_n188), .out0(\s[18] ));
  nona23aa1n02x4               g097(.a(new_n164), .b(new_n160), .c(new_n159), .d(new_n163), .out0(new_n193));
  oaoi13aa1n06x5               g098(.a(new_n193), .b(new_n155), .c(new_n154), .d(new_n153), .o1(new_n194));
  inv000aa1n02x5               g099(.a(new_n185), .o1(new_n195));
  oaoi13aa1n04x5               g100(.a(new_n195), .b(new_n181), .c(new_n194), .d(new_n166), .o1(new_n196));
  xroi22aa1d06x4               g101(.a(new_n189), .b(\b[16] ), .c(new_n188), .d(\b[17] ), .out0(new_n197));
  inv000aa1n03x5               g102(.a(new_n197), .o1(new_n198));
  inv000aa1d42x5               g103(.a(\b[17] ), .o1(new_n199));
  oai022aa1d24x5               g104(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n200));
  oa0012aa1n02x5               g105(.a(new_n200), .b(new_n199), .c(new_n188), .o(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  aoai13aa1n02x7               g107(.a(new_n202), .b(new_n198), .c(new_n196), .d(new_n183), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[18] ), .o1(new_n207));
  nand22aa1n09x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  tech160nm_fixorc02aa1n02p5x5 g113(.a(\a[19] ), .b(\b[18] ), .out0(new_n209));
  aoai13aa1n03x5               g114(.a(new_n209), .b(new_n201), .c(new_n186), .d(new_n197), .o1(new_n210));
  xorc02aa1n12x5               g115(.a(\a[20] ), .b(\b[19] ), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n212), .b(new_n210), .c(new_n208), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n208), .o1(new_n214));
  aoi112aa1n02x5               g119(.a(new_n214), .b(new_n211), .c(new_n203), .d(new_n209), .o1(new_n215));
  nor002aa1n02x5               g120(.a(new_n213), .b(new_n215), .o1(\s[20] ));
  nano22aa1n12x5               g121(.a(new_n198), .b(new_n209), .c(new_n211), .out0(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  and002aa1n02x5               g123(.a(\b[19] ), .b(\a[20] ), .o(new_n219));
  oai122aa1n06x5               g124(.a(new_n200), .b(new_n206), .c(new_n207), .d(new_n188), .e(new_n199), .o1(new_n220));
  oai112aa1n04x5               g125(.a(new_n220), .b(new_n208), .c(\b[19] ), .d(\a[20] ), .o1(new_n221));
  norb02aa1n12x5               g126(.a(new_n221), .b(new_n219), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n04x5               g128(.a(new_n223), .b(new_n218), .c(new_n196), .d(new_n183), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nanp02aa1n06x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n226), .out0(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n222), .c(new_n186), .d(new_n217), .o1(new_n230));
  nor042aa1n09x5               g135(.a(\b[21] ), .b(\a[22] ), .o1(new_n231));
  nand42aa1n06x5               g136(.a(\b[21] ), .b(\a[22] ), .o1(new_n232));
  nanb02aa1d36x5               g137(.a(new_n231), .b(new_n232), .out0(new_n233));
  aoi012aa1n03x5               g138(.a(new_n233), .b(new_n230), .c(new_n227), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n233), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n226), .b(new_n235), .c(new_n224), .d(new_n228), .o1(new_n236));
  nor002aa1n02x5               g141(.a(new_n234), .b(new_n236), .o1(\s[22] ));
  xorc02aa1n02x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  nano23aa1n06x5               g143(.a(new_n226), .b(new_n231), .c(new_n232), .d(new_n228), .out0(new_n239));
  nand23aa1n03x5               g144(.a(new_n186), .b(new_n217), .c(new_n239), .o1(new_n240));
  tech160nm_fioai012aa1n05x5   g145(.a(new_n232), .b(new_n231), .c(new_n226), .o1(new_n241));
  aob012aa1n02x5               g146(.a(new_n241), .b(new_n222), .c(new_n239), .out0(new_n242));
  norb02aa1n06x4               g147(.a(new_n238), .b(new_n242), .out0(new_n243));
  nand42aa1n03x5               g148(.a(new_n240), .b(new_n243), .o1(new_n244));
  aoi013aa1n02x4               g149(.a(new_n242), .b(new_n186), .c(new_n217), .d(new_n239), .o1(new_n245));
  oai012aa1n02x5               g150(.a(new_n244), .b(new_n245), .c(new_n238), .o1(\s[23] ));
  and002aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .o(new_n247));
  xorc02aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .out0(new_n248));
  aoai13aa1n02x7               g153(.a(new_n248), .b(new_n247), .c(new_n240), .d(new_n243), .o1(new_n249));
  nona22aa1n03x5               g154(.a(new_n244), .b(new_n248), .c(new_n247), .out0(new_n250));
  nanp02aa1n03x5               g155(.a(new_n250), .b(new_n249), .o1(\s[24] ));
  inv000aa1d42x5               g156(.a(\a[23] ), .o1(new_n252));
  inv000aa1d42x5               g157(.a(\b[22] ), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n253), .b(new_n252), .o1(new_n254));
  tech160nm_finand02aa1n05x5   g159(.a(\b[23] ), .b(\a[24] ), .o1(new_n255));
  orn002aa1n24x5               g160(.a(\a[24] ), .b(\b[23] ), .o(new_n256));
  oai112aa1n06x5               g161(.a(new_n256), .b(new_n255), .c(new_n253), .d(new_n252), .o1(new_n257));
  nano22aa1n12x5               g162(.a(new_n257), .b(new_n239), .c(new_n254), .out0(new_n258));
  inv000aa1n06x5               g163(.a(new_n258), .o1(new_n259));
  nano32aa1n02x5               g164(.a(new_n259), .b(new_n197), .c(new_n209), .d(new_n211), .out0(new_n260));
  inv030aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  aoi112aa1n03x5               g166(.a(new_n257), .b(new_n241), .c(new_n252), .d(new_n253), .o1(new_n262));
  oaoi03aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n254), .o1(new_n263));
  nor042aa1n04x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  nano32aa1n03x7               g169(.a(new_n233), .b(new_n227), .c(new_n254), .d(new_n228), .out0(new_n265));
  nona23aa1n09x5               g170(.a(new_n221), .b(new_n265), .c(new_n257), .d(new_n219), .out0(new_n266));
  nand02aa1d10x5               g171(.a(new_n266), .b(new_n264), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n02x7               g173(.a(new_n268), .b(new_n261), .c(new_n196), .d(new_n183), .o1(new_n269));
  xorb03aa1n02x5               g174(.a(new_n269), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  inv040aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  aoai13aa1n03x5               g178(.a(new_n273), .b(new_n267), .c(new_n186), .d(new_n260), .o1(new_n274));
  xorc02aa1n12x5               g179(.a(\a[26] ), .b(\b[25] ), .out0(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  tech160nm_fiaoi012aa1n02p5x5 g181(.a(new_n276), .b(new_n274), .c(new_n272), .o1(new_n277));
  aoi112aa1n02x5               g182(.a(new_n271), .b(new_n275), .c(new_n269), .d(new_n273), .o1(new_n278));
  nor002aa1n02x5               g183(.a(new_n277), .b(new_n278), .o1(\s[26] ));
  and002aa1n06x5               g184(.a(new_n275), .b(new_n273), .o(new_n280));
  nand23aa1d12x5               g185(.a(new_n217), .b(new_n258), .c(new_n280), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[26] ), .b(\b[25] ), .c(new_n272), .carry(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  tech160nm_fiaoi012aa1n05x5   g188(.a(new_n283), .b(new_n267), .c(new_n280), .o1(new_n284));
  aoai13aa1n04x5               g189(.a(new_n284), .b(new_n281), .c(new_n196), .d(new_n183), .o1(new_n285));
  xorb03aa1n02x5               g190(.a(new_n285), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  inv040aa1n03x5               g192(.a(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[28] ), .b(\b[27] ), .out0(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  nanp02aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n281), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n280), .o1(new_n293));
  aoai13aa1n06x5               g198(.a(new_n282), .b(new_n293), .c(new_n266), .d(new_n264), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n291), .b(new_n294), .c(new_n186), .d(new_n292), .o1(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n290), .b(new_n295), .c(new_n288), .o1(new_n296));
  aoi112aa1n03x4               g201(.a(new_n289), .b(new_n287), .c(new_n285), .d(new_n291), .o1(new_n297));
  nor002aa1n02x5               g202(.a(new_n296), .b(new_n297), .o1(\s[28] ));
  nano22aa1n02x4               g203(.a(new_n290), .b(new_n288), .c(new_n291), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n294), .c(new_n186), .d(new_n292), .o1(new_n300));
  oao003aa1n09x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n288), .carry(new_n301));
  xorc02aa1n06x5               g206(.a(\a[29] ), .b(\b[28] ), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n300), .c(new_n301), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n301), .o1(new_n305));
  aoi112aa1n03x4               g210(.a(new_n302), .b(new_n305), .c(new_n285), .d(new_n299), .o1(new_n306));
  nor002aa1n02x5               g211(.a(new_n304), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n113), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g213(.a(new_n303), .b(new_n289), .c(new_n291), .d(new_n288), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n294), .c(new_n186), .d(new_n292), .o1(new_n310));
  oao003aa1n12x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .carry(new_n311));
  xorc02aa1n12x5               g216(.a(\a[30] ), .b(\b[29] ), .out0(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n313), .b(new_n310), .c(new_n311), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n311), .o1(new_n315));
  aoi112aa1n03x4               g220(.a(new_n312), .b(new_n315), .c(new_n285), .d(new_n309), .o1(new_n316));
  nor002aa1n02x5               g221(.a(new_n314), .b(new_n316), .o1(\s[30] ));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  and003aa1n02x5               g223(.a(new_n299), .b(new_n312), .c(new_n302), .o(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n294), .c(new_n186), .d(new_n292), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n321));
  aoi012aa1n03x5               g226(.a(new_n318), .b(new_n320), .c(new_n321), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n318), .o1(new_n323));
  inv000aa1n02x5               g228(.a(new_n321), .o1(new_n324));
  aoi112aa1n02x5               g229(.a(new_n323), .b(new_n324), .c(new_n285), .d(new_n319), .o1(new_n325));
  norp02aa1n03x5               g230(.a(new_n322), .b(new_n325), .o1(\s[31] ));
  xnrb03aa1n02x5               g231(.a(new_n115), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g232(.a(\a[3] ), .b(\b[2] ), .c(new_n115), .o1(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g234(.a(new_n118), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g235(.a(new_n120), .b(new_n118), .c(new_n103), .o1(new_n331));
  xnrb03aa1n02x5               g236(.a(new_n331), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oab012aa1n06x5               g237(.a(new_n102), .b(new_n331), .c(new_n119), .out0(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n105), .c(new_n99), .out0(\s[7] ));
  oaoi03aa1n02x5               g239(.a(\a[7] ), .b(\b[6] ), .c(new_n333), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrc02aa1n02x5               g241(.a(new_n123), .b(new_n133), .out0(\s[9] ));
endmodule


