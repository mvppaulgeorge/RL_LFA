// Benchmark "adder" written by ABC on Wed Jul 17 18:54:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n336, new_n339, new_n340,
    new_n341, new_n343, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n06x4               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1n12x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1n04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  aoi012aa1n12x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  inv040aa1d32x5               g009(.a(\a[4] ), .o1(new_n105));
  inv040aa1d28x5               g010(.a(\b[3] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(new_n106), .b(new_n105), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand02aa1d04x5               g013(.a(new_n107), .b(new_n108), .o1(new_n109));
  inv040aa1d32x5               g014(.a(\a[3] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[2] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(new_n112), .b(new_n113), .o1(new_n114));
  nor003aa1n03x5               g019(.a(new_n104), .b(new_n109), .c(new_n114), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  oaoi03aa1n12x5               g021(.a(new_n105), .b(new_n106), .c(new_n116), .o1(new_n117));
  inv000aa1d42x5               g022(.a(new_n117), .o1(new_n118));
  xnrc02aa1n02x5               g023(.a(\b[5] ), .b(\a[6] ), .out0(new_n119));
  xnrc02aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .out0(new_n120));
  nor022aa1n08x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nand42aa1n08x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  norp02aa1n12x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nand42aa1n06x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nona23aa1n09x5               g029(.a(new_n124), .b(new_n122), .c(new_n121), .d(new_n123), .out0(new_n125));
  nor043aa1n03x5               g030(.a(new_n125), .b(new_n120), .c(new_n119), .o1(new_n126));
  oai012aa1n09x5               g031(.a(new_n126), .b(new_n115), .c(new_n118), .o1(new_n127));
  norb02aa1n06x4               g032(.a(new_n122), .b(new_n121), .out0(new_n128));
  nand42aa1n03x5               g033(.a(\b[5] ), .b(\a[6] ), .o1(new_n129));
  nano22aa1n03x7               g034(.a(new_n123), .b(new_n129), .c(new_n124), .out0(new_n130));
  oai022aa1n02x5               g035(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n131));
  tech160nm_fiao0012aa1n02p5x5 g036(.a(new_n121), .b(new_n123), .c(new_n122), .o(new_n132));
  aoi013aa1n06x4               g037(.a(new_n132), .b(new_n130), .c(new_n128), .d(new_n131), .o1(new_n133));
  nanp02aa1n06x5               g038(.a(new_n127), .b(new_n133), .o1(new_n134));
  nand02aa1n03x5               g039(.a(\b[8] ), .b(\a[9] ), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n100), .b(new_n134), .c(new_n135), .o1(new_n136));
  xnrc02aa1n02x5               g041(.a(new_n136), .b(new_n99), .out0(\s[10] ));
  norb02aa1n03x5               g042(.a(new_n135), .b(new_n100), .out0(new_n138));
  aoi012aa1d24x5               g043(.a(new_n97), .b(new_n100), .c(new_n98), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  aoi013aa1n06x4               g045(.a(new_n140), .b(new_n134), .c(new_n138), .d(new_n99), .o1(new_n141));
  nor002aa1d32x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  nand02aa1d06x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n141), .b(new_n144), .c(new_n143), .out0(\s[11] ));
  norb02aa1n15x5               g050(.a(new_n144), .b(new_n142), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  nor042aa1n03x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nand02aa1d08x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nanb02aa1n02x5               g054(.a(new_n148), .b(new_n149), .out0(new_n150));
  oaoi13aa1n06x5               g055(.a(new_n150), .b(new_n143), .c(new_n141), .d(new_n147), .o1(new_n151));
  oai112aa1n02x7               g056(.a(new_n150), .b(new_n143), .c(new_n141), .d(new_n147), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(\s[12] ));
  nano23aa1n03x7               g058(.a(new_n100), .b(new_n148), .c(new_n149), .d(new_n135), .out0(new_n154));
  nand23aa1n03x5               g059(.a(new_n154), .b(new_n99), .c(new_n146), .o1(new_n155));
  nanb03aa1n12x5               g060(.a(new_n142), .b(new_n149), .c(new_n144), .out0(new_n156));
  aoi012aa1n09x5               g061(.a(new_n148), .b(new_n142), .c(new_n149), .o1(new_n157));
  oai012aa1d24x5               g062(.a(new_n157), .b(new_n156), .c(new_n139), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n159), .b(new_n155), .c(new_n127), .d(new_n133), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n16x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand22aa1n04x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n162), .b(new_n160), .c(new_n163), .o1(new_n164));
  xnrb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  oai013aa1n06x5               g070(.a(new_n117), .b(new_n104), .c(new_n109), .d(new_n114), .o1(new_n166));
  nanp03aa1n03x5               g071(.a(new_n130), .b(new_n128), .c(new_n131), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n132), .b(new_n167), .out0(new_n168));
  nano32aa1n03x7               g073(.a(new_n150), .b(new_n146), .c(new_n138), .d(new_n99), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n168), .c(new_n166), .d(new_n126), .o1(new_n170));
  nor002aa1d32x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand22aa1n12x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nona23aa1n03x5               g077(.a(new_n172), .b(new_n163), .c(new_n162), .d(new_n171), .out0(new_n173));
  aoi012aa1d18x5               g078(.a(new_n171), .b(new_n162), .c(new_n172), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n173), .c(new_n170), .d(new_n159), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  nano23aa1n03x7               g083(.a(new_n162), .b(new_n171), .c(new_n172), .d(new_n163), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n174), .o1(new_n180));
  nanp02aa1n04x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  nanb02aa1n12x5               g086(.a(new_n177), .b(new_n181), .out0(new_n182));
  inv030aa1n02x5               g087(.a(new_n182), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n183), .b(new_n180), .c(new_n160), .d(new_n179), .o1(new_n184));
  nor042aa1n06x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nand02aa1n04x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nanb02aa1n09x5               g091(.a(new_n185), .b(new_n186), .out0(new_n187));
  aoi012aa1n02x5               g092(.a(new_n187), .b(new_n184), .c(new_n178), .o1(new_n188));
  inv000aa1n02x5               g093(.a(new_n187), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(new_n177), .b(new_n189), .c(new_n175), .d(new_n183), .o1(new_n190));
  norp02aa1n02x5               g095(.a(new_n188), .b(new_n190), .o1(\s[16] ));
  nor043aa1n06x5               g096(.a(new_n173), .b(new_n182), .c(new_n187), .o1(new_n192));
  nand22aa1n03x5               g097(.a(new_n169), .b(new_n192), .o1(new_n193));
  nanb03aa1n02x5               g098(.a(new_n177), .b(new_n186), .c(new_n181), .out0(new_n194));
  aoi012aa1n02x5               g099(.a(new_n185), .b(new_n177), .c(new_n186), .o1(new_n195));
  oai012aa1n06x5               g100(.a(new_n195), .b(new_n194), .c(new_n174), .o1(new_n196));
  aoi012aa1d24x5               g101(.a(new_n196), .b(new_n192), .c(new_n158), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n193), .c(new_n127), .d(new_n133), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g104(.a(\a[18] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\a[17] ), .o1(new_n201));
  inv000aa1d42x5               g106(.a(\b[16] ), .o1(new_n202));
  oaoi03aa1n03x5               g107(.a(new_n201), .b(new_n202), .c(new_n198), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[17] ), .c(new_n200), .out0(\s[18] ));
  nano32aa1n03x7               g109(.a(new_n155), .b(new_n189), .c(new_n179), .d(new_n183), .out0(new_n205));
  aoai13aa1n12x5               g110(.a(new_n205), .b(new_n168), .c(new_n166), .d(new_n126), .o1(new_n206));
  xroi22aa1d06x4               g111(.a(new_n201), .b(\b[16] ), .c(new_n200), .d(\b[17] ), .out0(new_n207));
  inv000aa1n02x5               g112(.a(new_n207), .o1(new_n208));
  nor042aa1n02x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  aoi112aa1n09x5               g114(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n210));
  nor002aa1n02x5               g115(.a(new_n210), .b(new_n209), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n208), .c(new_n206), .d(new_n197), .o1(new_n212));
  xorb03aa1n03x5               g117(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  inv040aa1n02x5               g120(.a(new_n215), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n211), .o1(new_n217));
  nand02aa1d24x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  norb02aa1n15x5               g123(.a(new_n218), .b(new_n215), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n198), .d(new_n207), .o1(new_n220));
  xnrc02aa1n06x5               g125(.a(\b[19] ), .b(\a[20] ), .out0(new_n221));
  aoi012aa1n03x5               g126(.a(new_n221), .b(new_n220), .c(new_n216), .o1(new_n222));
  inv040aa1n02x5               g127(.a(new_n221), .o1(new_n223));
  aoi112aa1n03x5               g128(.a(new_n215), .b(new_n223), .c(new_n212), .d(new_n219), .o1(new_n224));
  nor002aa1n02x5               g129(.a(new_n222), .b(new_n224), .o1(\s[20] ));
  nand23aa1d12x5               g130(.a(new_n207), .b(new_n219), .c(new_n223), .o1(new_n226));
  nanp02aa1n02x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  oai112aa1n06x5               g132(.a(new_n219), .b(new_n227), .c(new_n210), .d(new_n209), .o1(new_n228));
  oao003aa1n09x5               g133(.a(\a[20] ), .b(\b[19] ), .c(new_n216), .carry(new_n229));
  nand02aa1d06x5               g134(.a(new_n228), .b(new_n229), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n226), .c(new_n206), .d(new_n197), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n226), .o1(new_n236));
  nand42aa1n20x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n234), .out0(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n230), .c(new_n198), .d(new_n236), .o1(new_n239));
  nor002aa1n16x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nand02aa1d28x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  norb02aa1n12x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n03x5               g148(.a(new_n243), .b(new_n239), .c(new_n235), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(new_n234), .b(new_n242), .c(new_n232), .d(new_n238), .o1(new_n245));
  nor002aa1n02x5               g150(.a(new_n244), .b(new_n245), .o1(\s[22] ));
  nano23aa1d15x5               g151(.a(new_n234), .b(new_n240), .c(new_n241), .d(new_n237), .out0(new_n247));
  nano32aa1n03x7               g152(.a(new_n208), .b(new_n247), .c(new_n219), .d(new_n223), .out0(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoi012aa1n06x5               g154(.a(new_n240), .b(new_n234), .c(new_n241), .o1(new_n250));
  inv000aa1n06x5               g155(.a(new_n250), .o1(new_n251));
  aoi012aa1d18x5               g156(.a(new_n251), .b(new_n230), .c(new_n247), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n249), .c(new_n206), .d(new_n197), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1d18x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  inv040aa1n03x5               g160(.a(new_n255), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n252), .o1(new_n257));
  nand42aa1n04x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  norb02aa1n03x5               g163(.a(new_n258), .b(new_n255), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n257), .c(new_n198), .d(new_n248), .o1(new_n260));
  xnrc02aa1n02x5               g165(.a(\b[23] ), .b(\a[24] ), .out0(new_n261));
  aoi012aa1n03x5               g166(.a(new_n261), .b(new_n260), .c(new_n256), .o1(new_n262));
  tech160nm_fixorc02aa1n04x5   g167(.a(\a[24] ), .b(\b[23] ), .out0(new_n263));
  aoi112aa1n02x5               g168(.a(new_n255), .b(new_n263), .c(new_n253), .d(new_n259), .o1(new_n264));
  nor002aa1n02x5               g169(.a(new_n262), .b(new_n264), .o1(\s[24] ));
  nand23aa1n06x5               g170(.a(new_n247), .b(new_n259), .c(new_n263), .o1(new_n266));
  nano32aa1n02x4               g171(.a(new_n266), .b(new_n207), .c(new_n219), .d(new_n223), .out0(new_n267));
  inv020aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  tech160nm_finand02aa1n03p5x5 g173(.a(\b[23] ), .b(\a[24] ), .o1(new_n269));
  nano22aa1n03x5               g174(.a(new_n255), .b(new_n258), .c(new_n269), .out0(new_n270));
  oaoi03aa1n12x5               g175(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .o1(new_n271));
  aoi012aa1n12x5               g176(.a(new_n271), .b(new_n251), .c(new_n270), .o1(new_n272));
  aoai13aa1n12x5               g177(.a(new_n272), .b(new_n266), .c(new_n228), .d(new_n229), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n02x5               g179(.a(new_n274), .b(new_n268), .c(new_n206), .d(new_n197), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  inv000aa1n02x5               g182(.a(new_n277), .o1(new_n278));
  tech160nm_fixorc02aa1n03p5x5 g183(.a(\a[25] ), .b(\b[24] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n273), .c(new_n198), .d(new_n267), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[26] ), .b(\b[25] ), .out0(new_n281));
  inv000aa1d42x5               g186(.a(new_n281), .o1(new_n282));
  aoi012aa1n03x5               g187(.a(new_n282), .b(new_n280), .c(new_n278), .o1(new_n283));
  aoi112aa1n03x4               g188(.a(new_n277), .b(new_n281), .c(new_n275), .d(new_n279), .o1(new_n284));
  nor002aa1n02x5               g189(.a(new_n283), .b(new_n284), .o1(\s[26] ));
  nano32aa1n03x7               g190(.a(new_n261), .b(new_n259), .c(new_n242), .d(new_n238), .out0(new_n286));
  and002aa1n02x5               g191(.a(new_n281), .b(new_n279), .o(new_n287));
  nano22aa1n06x5               g192(.a(new_n226), .b(new_n286), .c(new_n287), .out0(new_n288));
  inv020aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[26] ), .b(\b[25] ), .c(new_n278), .carry(new_n290));
  aobi12aa1n06x5               g195(.a(new_n290), .b(new_n273), .c(new_n287), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n289), .c(new_n206), .d(new_n197), .o1(new_n292));
  xorb03aa1n03x5               g197(.a(new_n292), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv000aa1n03x5               g199(.a(new_n294), .o1(new_n295));
  nand02aa1d04x5               g200(.a(new_n230), .b(new_n286), .o1(new_n296));
  nanp02aa1n02x5               g201(.a(new_n281), .b(new_n279), .o1(new_n297));
  aoai13aa1n04x5               g202(.a(new_n290), .b(new_n297), .c(new_n296), .d(new_n272), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[27] ), .b(\b[26] ), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n198), .d(new_n288), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[28] ), .b(\b[27] ), .out0(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  aoi012aa1n02x7               g207(.a(new_n302), .b(new_n300), .c(new_n295), .o1(new_n303));
  aoi112aa1n03x4               g208(.a(new_n294), .b(new_n301), .c(new_n292), .d(new_n299), .o1(new_n304));
  norp02aa1n03x5               g209(.a(new_n303), .b(new_n304), .o1(\s[28] ));
  and002aa1n02x5               g210(.a(new_n301), .b(new_n299), .o(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n298), .c(new_n198), .d(new_n288), .o1(new_n307));
  oao003aa1n09x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n308));
  tech160nm_fixorc02aa1n03p5x5 g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  aoi012aa1n03x5               g215(.a(new_n310), .b(new_n307), .c(new_n308), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n308), .o1(new_n312));
  aoi112aa1n03x4               g217(.a(new_n309), .b(new_n312), .c(new_n292), .d(new_n306), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g220(.a(new_n310), .b(new_n299), .c(new_n301), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n298), .c(new_n198), .d(new_n288), .o1(new_n317));
  tech160nm_fioaoi03aa1n03p5x5 g222(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .o1(new_n318));
  inv000aa1n03x5               g223(.a(new_n318), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .out0(new_n320));
  inv000aa1n02x5               g225(.a(new_n320), .o1(new_n321));
  aoi012aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n319), .o1(new_n322));
  aoi112aa1n03x4               g227(.a(new_n320), .b(new_n318), .c(new_n292), .d(new_n316), .o1(new_n323));
  norp02aa1n03x5               g228(.a(new_n322), .b(new_n323), .o1(\s[30] ));
  nano32aa1n02x4               g229(.a(new_n321), .b(new_n309), .c(new_n301), .d(new_n299), .out0(new_n325));
  oao003aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .c(new_n319), .carry(new_n326));
  inv000aa1n02x5               g231(.a(new_n326), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[31] ), .b(\b[30] ), .out0(new_n328));
  aoi112aa1n03x4               g233(.a(new_n328), .b(new_n327), .c(new_n292), .d(new_n325), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n325), .b(new_n298), .c(new_n198), .d(new_n288), .o1(new_n330));
  inv000aa1d42x5               g235(.a(new_n328), .o1(new_n331));
  tech160nm_fiaoi012aa1n02p5x5 g236(.a(new_n331), .b(new_n330), .c(new_n326), .o1(new_n332));
  norp02aa1n03x5               g237(.a(new_n332), .b(new_n329), .o1(\s[31] ));
  xnbna2aa1n03x5               g238(.a(new_n104), .b(new_n113), .c(new_n112), .out0(\s[3] ));
  orn002aa1n02x5               g239(.a(new_n104), .b(new_n114), .o(new_n335));
  aoi022aa1n02x5               g240(.a(new_n107), .b(new_n108), .c(new_n111), .d(new_n110), .o1(new_n336));
  aoi022aa1n02x5               g241(.a(new_n166), .b(new_n107), .c(new_n336), .d(new_n335), .o1(\s[4] ));
  xorb03aa1n02x5               g242(.a(new_n166), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g243(.a(\a[6] ), .o1(new_n339));
  norp02aa1n02x5               g244(.a(\b[4] ), .b(\a[5] ), .o1(new_n340));
  aoib12aa1n02x5               g245(.a(new_n340), .b(new_n166), .c(new_n120), .out0(new_n341));
  xorb03aa1n02x5               g246(.a(new_n341), .b(\b[5] ), .c(new_n339), .out0(\s[6] ));
  norb02aa1n02x5               g247(.a(new_n124), .b(new_n123), .out0(new_n343));
  oaib12aa1n03x5               g248(.a(new_n341), .b(\b[5] ), .c(new_n339), .out0(new_n344));
  xobna2aa1n03x5               g249(.a(new_n343), .b(new_n344), .c(new_n129), .out0(\s[7] ));
  tech160nm_fiaoi012aa1n05x5   g250(.a(new_n123), .b(new_n344), .c(new_n130), .o1(new_n346));
  xnrc02aa1n02x5               g251(.a(new_n346), .b(new_n128), .out0(\s[8] ));
  xnbna2aa1n03x5               g252(.a(new_n138), .b(new_n127), .c(new_n133), .out0(\s[9] ));
endmodule


