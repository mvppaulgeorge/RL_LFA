// Benchmark "adder" written by ABC on Wed Jul 17 20:16:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n332, new_n335, new_n337, new_n338, new_n339, new_n340, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1n09x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  and002aa1n06x5               g004(.a(\b[3] ), .b(\a[4] ), .o(new_n100));
  inv040aa1d32x5               g005(.a(\a[3] ), .o1(new_n101));
  inv030aa1d32x5               g006(.a(\b[2] ), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(new_n103), .b(new_n104), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nand22aa1n04x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nand22aa1n09x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  aoi012aa1n12x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  oa0022aa1n09x5               g014(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n110));
  oaoi13aa1n12x5               g015(.a(new_n100), .b(new_n110), .c(new_n109), .d(new_n105), .o1(new_n111));
  xnrc02aa1n02x5               g016(.a(\b[5] ), .b(\a[6] ), .out0(new_n112));
  nor002aa1n12x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nor002aa1d32x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  xnrc02aa1n06x5               g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  nor043aa1n02x5               g023(.a(new_n117), .b(new_n118), .c(new_n112), .o1(new_n119));
  and002aa1n02x5               g024(.a(\b[5] ), .b(\a[6] ), .o(new_n120));
  oai012aa1n02x5               g025(.a(new_n114), .b(new_n116), .c(new_n113), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\a[5] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\a[6] ), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\b[4] ), .o1(new_n124));
  aboi22aa1n12x5               g029(.a(\b[5] ), .b(new_n123), .c(new_n122), .d(new_n124), .out0(new_n125));
  oai013aa1n03x5               g030(.a(new_n121), .b(new_n117), .c(new_n120), .d(new_n125), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n126), .c(new_n111), .d(new_n119), .o1(new_n128));
  nor002aa1d32x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1n03x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  inv030aa1n02x5               g036(.a(new_n131), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n128), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g038(.a(new_n129), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n130), .o1(new_n135));
  nor042aa1n06x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanp02aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanb02aa1n09x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  aoi113aa1n03x7               g043(.a(new_n138), .b(new_n135), .c(new_n128), .d(new_n134), .e(new_n99), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n111), .b(new_n119), .o1(new_n140));
  nano23aa1n03x7               g045(.a(new_n116), .b(new_n113), .c(new_n114), .d(new_n115), .out0(new_n141));
  norp02aa1n02x5               g046(.a(new_n125), .b(new_n120), .o1(new_n142));
  aobi12aa1n06x5               g047(.a(new_n121), .b(new_n141), .c(new_n142), .out0(new_n143));
  inv000aa1d42x5               g048(.a(new_n127), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n99), .b(new_n144), .c(new_n140), .d(new_n143), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n138), .o1(new_n146));
  aoai13aa1n12x5               g051(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  aoi112aa1n02x5               g053(.a(new_n148), .b(new_n146), .c(new_n145), .d(new_n132), .o1(new_n149));
  norp02aa1n02x5               g054(.a(new_n149), .b(new_n139), .o1(\s[11] ));
  nor002aa1n16x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nand02aa1n03x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  aoi112aa1n03x5               g058(.a(new_n139), .b(new_n136), .c(new_n152), .d(new_n153), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n146), .b(new_n148), .c(new_n145), .d(new_n132), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n151), .b(new_n153), .out0(new_n156));
  oaoi13aa1n02x5               g061(.a(new_n156), .b(new_n155), .c(\a[11] ), .d(\b[10] ), .o1(new_n157));
  norp02aa1n03x5               g062(.a(new_n157), .b(new_n154), .o1(\s[12] ));
  nona23aa1n03x5               g063(.a(new_n153), .b(new_n137), .c(new_n136), .d(new_n151), .out0(new_n159));
  norb03aa1n02x7               g064(.a(new_n127), .b(new_n159), .c(new_n131), .out0(new_n160));
  aoai13aa1n03x5               g065(.a(new_n160), .b(new_n126), .c(new_n111), .d(new_n119), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(new_n136), .b(new_n153), .o1(new_n162));
  nor043aa1n03x5               g067(.a(new_n147), .b(new_n138), .c(new_n156), .o1(new_n163));
  nano22aa1n03x7               g068(.a(new_n163), .b(new_n152), .c(new_n162), .out0(new_n164));
  nor002aa1d32x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand42aa1d28x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n161), .c(new_n164), .out0(\s[13] ));
  inv040aa1n08x5               g073(.a(new_n165), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n100), .o1(new_n170));
  tech160nm_fioai012aa1n04x5   g075(.a(new_n110), .b(new_n109), .c(new_n105), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n170), .o1(new_n172));
  nona22aa1n02x4               g077(.a(new_n141), .b(new_n118), .c(new_n112), .out0(new_n173));
  tech160nm_fioai012aa1n05x5   g078(.a(new_n143), .b(new_n172), .c(new_n173), .o1(new_n174));
  oai112aa1n06x5               g079(.a(new_n162), .b(new_n152), .c(new_n159), .d(new_n147), .o1(new_n175));
  aoai13aa1n02x5               g080(.a(new_n167), .b(new_n175), .c(new_n174), .d(new_n160), .o1(new_n176));
  nor042aa1n04x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nand42aa1n16x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n176), .c(new_n169), .out0(\s[14] ));
  oaoi03aa1n12x5               g085(.a(\a[14] ), .b(\b[13] ), .c(new_n169), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  nano23aa1d15x5               g087(.a(new_n165), .b(new_n177), .c(new_n178), .d(new_n166), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  aoai13aa1n04x5               g089(.a(new_n182), .b(new_n184), .c(new_n161), .d(new_n164), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  nand42aa1n02x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  norb02aa1n06x4               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  nor042aa1n02x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nand42aa1n02x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  norb02aa1n09x5               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  aoi112aa1n02x5               g097(.a(new_n192), .b(new_n187), .c(new_n185), .d(new_n189), .o1(new_n193));
  aoai13aa1n03x5               g098(.a(new_n192), .b(new_n187), .c(new_n185), .d(new_n188), .o1(new_n194));
  norb02aa1n02x7               g099(.a(new_n194), .b(new_n193), .out0(\s[16] ));
  nano23aa1n06x5               g100(.a(new_n136), .b(new_n151), .c(new_n153), .d(new_n137), .out0(new_n196));
  nand23aa1n09x5               g101(.a(new_n183), .b(new_n189), .c(new_n192), .o1(new_n197));
  nano32aa1n03x7               g102(.a(new_n197), .b(new_n196), .c(new_n132), .d(new_n127), .out0(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n126), .c(new_n111), .d(new_n119), .o1(new_n199));
  inv000aa1n02x5               g104(.a(new_n197), .o1(new_n200));
  aoi112aa1n02x5               g105(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n201));
  nanp03aa1n02x5               g106(.a(new_n181), .b(new_n189), .c(new_n192), .o1(new_n202));
  nona22aa1n03x5               g107(.a(new_n202), .b(new_n201), .c(new_n190), .out0(new_n203));
  aoi012aa1n12x5               g108(.a(new_n203), .b(new_n175), .c(new_n200), .o1(new_n204));
  xorc02aa1n12x5               g109(.a(\a[17] ), .b(\b[16] ), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n199), .c(new_n204), .out0(\s[17] ));
  inv000aa1d42x5               g111(.a(\a[17] ), .o1(new_n207));
  inv000aa1d42x5               g112(.a(\b[16] ), .o1(new_n208));
  nanp02aa1n06x5               g113(.a(new_n199), .b(new_n204), .o1(new_n209));
  tech160nm_fioaoi03aa1n03p5x5 g114(.a(new_n207), .b(new_n208), .c(new_n209), .o1(new_n210));
  nor022aa1n04x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nand42aa1n03x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nanb02aa1n12x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  xorc02aa1n02x5               g118(.a(new_n210), .b(new_n213), .out0(\s[18] ));
  norb02aa1n03x5               g119(.a(new_n205), .b(new_n213), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n04x5               g121(.a(new_n212), .b(new_n211), .c(new_n207), .d(new_n208), .o1(new_n217));
  aoai13aa1n04x5               g122(.a(new_n217), .b(new_n216), .c(new_n199), .d(new_n204), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  nand42aa1n06x5               g126(.a(\b[18] ), .b(\a[19] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\b[19] ), .o1(new_n223));
  nanb02aa1n02x5               g128(.a(\a[20] ), .b(new_n223), .out0(new_n224));
  nand42aa1n04x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  aoi122aa1n03x5               g130(.a(new_n221), .b(new_n225), .c(new_n224), .d(new_n218), .e(new_n222), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n221), .o1(new_n227));
  nanb02aa1n12x5               g132(.a(new_n221), .b(new_n222), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  nanp02aa1n03x5               g134(.a(new_n218), .b(new_n229), .o1(new_n230));
  nanp02aa1n02x5               g135(.a(new_n224), .b(new_n225), .o1(new_n231));
  tech160nm_fiaoi012aa1n02p5x5 g136(.a(new_n231), .b(new_n230), .c(new_n227), .o1(new_n232));
  norp02aa1n03x5               g137(.a(new_n232), .b(new_n226), .o1(\s[20] ));
  nona23aa1n02x4               g138(.a(new_n229), .b(new_n205), .c(new_n213), .d(new_n231), .out0(new_n234));
  nand42aa1n03x5               g139(.a(new_n221), .b(new_n225), .o1(new_n235));
  nor043aa1n03x5               g140(.a(new_n217), .b(new_n228), .c(new_n231), .o1(new_n236));
  nano22aa1n03x7               g141(.a(new_n236), .b(new_n224), .c(new_n235), .out0(new_n237));
  aoai13aa1n04x5               g142(.a(new_n237), .b(new_n234), .c(new_n199), .d(new_n204), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  xnrc02aa1n12x5               g145(.a(\b[20] ), .b(\a[21] ), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoi112aa1n02x7               g149(.a(new_n240), .b(new_n244), .c(new_n238), .d(new_n242), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n244), .b(new_n240), .c(new_n238), .d(new_n242), .o1(new_n246));
  norb02aa1n02x7               g151(.a(new_n246), .b(new_n245), .out0(\s[22] ));
  norp02aa1n02x5               g152(.a(\b[19] ), .b(\a[20] ), .o1(new_n248));
  nona23aa1n12x5               g153(.a(new_n225), .b(new_n222), .c(new_n221), .d(new_n248), .out0(new_n249));
  nor042aa1n06x5               g154(.a(new_n243), .b(new_n241), .o1(new_n250));
  nona23aa1n12x5               g155(.a(new_n250), .b(new_n205), .c(new_n249), .d(new_n213), .out0(new_n251));
  oai112aa1n03x5               g156(.a(new_n235), .b(new_n224), .c(new_n249), .d(new_n217), .o1(new_n252));
  inv020aa1n02x5               g157(.a(new_n240), .o1(new_n253));
  tech160nm_fioaoi03aa1n03p5x5 g158(.a(\a[22] ), .b(\b[21] ), .c(new_n253), .o1(new_n254));
  aoi012aa1n02x5               g159(.a(new_n254), .b(new_n252), .c(new_n250), .o1(new_n255));
  aoai13aa1n04x5               g160(.a(new_n255), .b(new_n251), .c(new_n199), .d(new_n204), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  xorc02aa1n12x5               g164(.a(\a[24] ), .b(\b[23] ), .out0(new_n260));
  aoi112aa1n02x7               g165(.a(new_n258), .b(new_n260), .c(new_n256), .d(new_n259), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n260), .b(new_n258), .c(new_n256), .d(new_n259), .o1(new_n262));
  norb02aa1n02x7               g167(.a(new_n262), .b(new_n261), .out0(\s[24] ));
  nanp02aa1n02x5               g168(.a(new_n260), .b(new_n259), .o1(new_n264));
  nona23aa1n06x5               g169(.a(new_n250), .b(new_n215), .c(new_n264), .d(new_n249), .out0(new_n265));
  xnrc02aa1n02x5               g170(.a(\b[22] ), .b(\a[23] ), .out0(new_n266));
  norb02aa1n02x5               g171(.a(new_n260), .b(new_n266), .out0(new_n267));
  norp02aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .o1(new_n268));
  aoi112aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n269));
  nanp03aa1n02x5               g174(.a(new_n254), .b(new_n259), .c(new_n260), .o1(new_n270));
  nona22aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n268), .out0(new_n271));
  aoi013aa1n02x4               g176(.a(new_n271), .b(new_n252), .c(new_n250), .d(new_n267), .o1(new_n272));
  aoai13aa1n04x5               g177(.a(new_n272), .b(new_n265), .c(new_n199), .d(new_n204), .o1(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor002aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  aoi112aa1n03x5               g182(.a(new_n275), .b(new_n277), .c(new_n273), .d(new_n276), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n277), .b(new_n275), .c(new_n273), .d(new_n276), .o1(new_n279));
  norb02aa1n03x4               g184(.a(new_n279), .b(new_n278), .out0(\s[26] ));
  aoi113aa1n02x5               g185(.a(new_n201), .b(new_n190), .c(new_n181), .d(new_n189), .e(new_n191), .o1(new_n281));
  tech160nm_fioai012aa1n05x5   g186(.a(new_n281), .b(new_n164), .c(new_n197), .o1(new_n282));
  and002aa1n09x5               g187(.a(new_n277), .b(new_n276), .o(new_n283));
  nano22aa1n03x7               g188(.a(new_n251), .b(new_n267), .c(new_n283), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n282), .c(new_n174), .d(new_n198), .o1(new_n285));
  nano22aa1n03x7               g190(.a(new_n237), .b(new_n250), .c(new_n267), .out0(new_n286));
  inv000aa1d42x5               g191(.a(\a[26] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[25] ), .o1(new_n288));
  oaoi03aa1n03x5               g193(.a(new_n287), .b(new_n288), .c(new_n275), .o1(new_n289));
  inv000aa1n02x5               g194(.a(new_n289), .o1(new_n290));
  oaoi13aa1n12x5               g195(.a(new_n290), .b(new_n283), .c(new_n286), .d(new_n271), .o1(new_n291));
  xorc02aa1n12x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  xnbna2aa1n06x5               g197(.a(new_n292), .b(new_n291), .c(new_n285), .out0(\s[27] ));
  nor042aa1n03x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  aobi12aa1n02x7               g200(.a(new_n292), .b(new_n291), .c(new_n285), .out0(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[27] ), .b(\a[28] ), .out0(new_n297));
  nano22aa1n02x4               g202(.a(new_n296), .b(new_n295), .c(new_n297), .out0(new_n298));
  nona32aa1n02x5               g203(.a(new_n252), .b(new_n264), .c(new_n243), .d(new_n241), .out0(new_n299));
  inv040aa1n03x5               g204(.a(new_n271), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n283), .o1(new_n301));
  aoai13aa1n06x5               g206(.a(new_n289), .b(new_n301), .c(new_n299), .d(new_n300), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n292), .b(new_n302), .c(new_n209), .d(new_n284), .o1(new_n303));
  aoi012aa1n03x5               g208(.a(new_n297), .b(new_n303), .c(new_n295), .o1(new_n304));
  nor002aa1n02x5               g209(.a(new_n304), .b(new_n298), .o1(\s[28] ));
  xnrc02aa1n02x5               g210(.a(\b[28] ), .b(\a[29] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n292), .b(new_n297), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n302), .c(new_n209), .d(new_n284), .o1(new_n308));
  oao003aa1n03x5               g213(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n309));
  aoi012aa1n02x7               g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  aobi12aa1n02x7               g215(.a(new_n307), .b(new_n291), .c(new_n285), .out0(new_n311));
  nano22aa1n03x5               g216(.a(new_n311), .b(new_n306), .c(new_n309), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n310), .b(new_n312), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g219(.a(new_n292), .b(new_n306), .c(new_n297), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n302), .c(new_n209), .d(new_n284), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .out0(new_n318));
  aoi012aa1n03x5               g223(.a(new_n318), .b(new_n316), .c(new_n317), .o1(new_n319));
  aobi12aa1n06x5               g224(.a(new_n315), .b(new_n291), .c(new_n285), .out0(new_n320));
  nano22aa1n02x4               g225(.a(new_n320), .b(new_n317), .c(new_n318), .out0(new_n321));
  nor002aa1n02x5               g226(.a(new_n319), .b(new_n321), .o1(\s[30] ));
  xnrc02aa1n02x5               g227(.a(\b[30] ), .b(\a[31] ), .out0(new_n323));
  norb02aa1n02x5               g228(.a(new_n315), .b(new_n318), .out0(new_n324));
  aobi12aa1n02x7               g229(.a(new_n324), .b(new_n291), .c(new_n285), .out0(new_n325));
  oao003aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n326));
  nano22aa1n03x5               g231(.a(new_n325), .b(new_n323), .c(new_n326), .out0(new_n327));
  aoai13aa1n03x5               g232(.a(new_n324), .b(new_n302), .c(new_n209), .d(new_n284), .o1(new_n328));
  aoi012aa1n03x5               g233(.a(new_n323), .b(new_n328), .c(new_n326), .o1(new_n329));
  nor002aa1n02x5               g234(.a(new_n329), .b(new_n327), .o1(\s[31] ));
  xnbna2aa1n03x5               g235(.a(new_n109), .b(new_n103), .c(new_n104), .out0(\s[3] ));
  oaoi03aa1n02x5               g236(.a(\a[3] ), .b(\b[2] ), .c(new_n109), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnbna2aa1n03x5               g238(.a(new_n118), .b(new_n171), .c(new_n170), .out0(\s[5] ));
  oaoi03aa1n02x5               g239(.a(new_n122), .b(new_n124), .c(new_n111), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[5] ), .c(new_n123), .out0(\s[6] ));
  oai012aa1n02x5               g241(.a(new_n125), .b(new_n172), .c(new_n118), .o1(new_n337));
  nona23aa1n02x4               g242(.a(new_n337), .b(new_n115), .c(new_n120), .d(new_n116), .out0(new_n338));
  inv000aa1d42x5               g243(.a(new_n116), .o1(new_n339));
  aboi22aa1n03x5               g244(.a(new_n120), .b(new_n337), .c(new_n115), .d(new_n339), .out0(new_n340));
  norb02aa1n02x5               g245(.a(new_n338), .b(new_n340), .out0(\s[7] ));
  norb02aa1n02x5               g246(.a(new_n114), .b(new_n113), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n342), .b(new_n338), .c(new_n339), .out0(\s[8] ));
  xnbna2aa1n03x5               g248(.a(new_n127), .b(new_n140), .c(new_n143), .out0(\s[9] ));
endmodule


