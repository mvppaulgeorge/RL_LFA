// Benchmark "adder" written by ABC on Wed Jul 17 23:01:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n336, new_n338,
    new_n340, new_n342, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n09x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  norp02aa1n04x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nanp02aa1n06x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norb02aa1n09x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  nand22aa1n06x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nor042aa1n03x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nona22aa1n09x5               g010(.a(new_n104), .b(new_n105), .c(new_n103), .out0(new_n106));
  nor042aa1n06x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1n06x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nano22aa1n12x5               g013(.a(new_n107), .b(new_n104), .c(new_n108), .out0(new_n109));
  tech160nm_fiaoi012aa1n04x5   g014(.a(new_n100), .b(new_n107), .c(new_n101), .o1(new_n110));
  inv000aa1n02x5               g015(.a(new_n110), .o1(new_n111));
  aoi013aa1n06x4               g016(.a(new_n111), .b(new_n109), .c(new_n106), .d(new_n102), .o1(new_n112));
  nor042aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1n10x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n16x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n06x5               g021(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n117));
  nor002aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nand42aa1n08x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  norb02aa1n03x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  xorc02aa1n12x5               g025(.a(\a[5] ), .b(\b[4] ), .out0(new_n121));
  nand43aa1n06x5               g026(.a(new_n117), .b(new_n120), .c(new_n121), .o1(new_n122));
  orn002aa1n24x5               g027(.a(\a[5] ), .b(\b[4] ), .o(new_n123));
  nanb03aa1n06x5               g028(.a(new_n118), .b(new_n123), .c(new_n119), .out0(new_n124));
  inv000aa1d42x5               g029(.a(\b[7] ), .o1(new_n125));
  nanb02aa1n06x5               g030(.a(\a[8] ), .b(new_n125), .out0(new_n126));
  nanb02aa1n12x5               g031(.a(new_n115), .b(new_n116), .out0(new_n127));
  nano32aa1n02x4               g032(.a(new_n127), .b(new_n126), .c(new_n119), .d(new_n114), .out0(new_n128));
  aoi012aa1n02x5               g033(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n129));
  aobi12aa1n02x7               g034(.a(new_n129), .b(new_n128), .c(new_n124), .out0(new_n130));
  oai012aa1n03x5               g035(.a(new_n130), .b(new_n112), .c(new_n122), .o1(new_n131));
  aob012aa1n06x5               g036(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(new_n132));
  oai012aa1n02x5               g037(.a(new_n132), .b(\b[8] ), .c(\a[9] ), .o1(new_n133));
  norp02aa1n02x5               g038(.a(\b[8] ), .b(\a[9] ), .o1(new_n134));
  nona22aa1n06x5               g039(.a(new_n132), .b(new_n134), .c(new_n99), .out0(new_n135));
  aob012aa1n02x5               g040(.a(new_n135), .b(new_n133), .c(new_n99), .out0(\s[10] ));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  inv040aa1n08x5               g042(.a(new_n137), .o1(new_n138));
  aoi022aa1n02x5               g043(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n139));
  nand02aa1d28x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  aoi022aa1n02x5               g045(.a(new_n135), .b(new_n98), .c(new_n140), .d(new_n138), .o1(new_n141));
  aoi013aa1n02x4               g046(.a(new_n141), .b(new_n139), .c(new_n138), .d(new_n135), .o1(\s[11] ));
  nor042aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand22aa1n12x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n06x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  aoi112aa1n02x5               g050(.a(new_n137), .b(new_n145), .c(new_n135), .d(new_n139), .o1(new_n146));
  aoai13aa1n03x5               g051(.a(new_n145), .b(new_n137), .c(new_n135), .d(new_n139), .o1(new_n147));
  norb02aa1n03x4               g052(.a(new_n147), .b(new_n146), .out0(\s[12] ));
  nanp03aa1n06x5               g053(.a(new_n109), .b(new_n106), .c(new_n102), .o1(new_n149));
  aoi012aa1n06x5               g054(.a(new_n122), .b(new_n149), .c(new_n110), .o1(new_n150));
  aob012aa1n06x5               g055(.a(new_n129), .b(new_n128), .c(new_n124), .out0(new_n151));
  nano23aa1n03x7               g056(.a(new_n137), .b(new_n143), .c(new_n144), .d(new_n140), .out0(new_n152));
  xnrc02aa1n02x5               g057(.a(\b[8] ), .b(\a[9] ), .out0(new_n153));
  nona22aa1n02x4               g058(.a(new_n152), .b(new_n153), .c(new_n99), .out0(new_n154));
  oabi12aa1n02x5               g059(.a(new_n154), .b(new_n150), .c(new_n151), .out0(new_n155));
  tech160nm_fiao0012aa1n03p5x5 g060(.a(new_n97), .b(new_n134), .c(new_n98), .o(new_n156));
  oaoi03aa1n12x5               g061(.a(\a[12] ), .b(\b[11] ), .c(new_n138), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n157), .b(new_n152), .c(new_n156), .o1(new_n158));
  nor002aa1d32x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand02aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  aob012aa1n02x5               g066(.a(new_n161), .b(new_n155), .c(new_n158), .out0(new_n162));
  aoi112aa1n02x5               g067(.a(new_n161), .b(new_n157), .c(new_n152), .d(new_n156), .o1(new_n163));
  aobi12aa1n02x5               g068(.a(new_n162), .b(new_n163), .c(new_n155), .out0(\s[13] ));
  nor002aa1d32x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand02aa1n06x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  aoib12aa1n02x5               g071(.a(new_n159), .b(new_n166), .c(new_n165), .out0(new_n167));
  nona23aa1d24x5               g072(.a(new_n166), .b(new_n160), .c(new_n159), .d(new_n165), .out0(new_n168));
  nona22aa1n02x4               g073(.a(new_n131), .b(new_n154), .c(new_n168), .out0(new_n169));
  norb02aa1n12x5               g074(.a(new_n140), .b(new_n137), .out0(new_n170));
  aoi112aa1n09x5               g075(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n171));
  oai112aa1n06x5               g076(.a(new_n145), .b(new_n170), .c(new_n171), .d(new_n97), .o1(new_n172));
  inv030aa1n08x5               g077(.a(new_n157), .o1(new_n173));
  tech160nm_fioai012aa1n03p5x5 g078(.a(new_n166), .b(new_n165), .c(new_n159), .o1(new_n174));
  aoai13aa1n12x5               g079(.a(new_n174), .b(new_n168), .c(new_n172), .d(new_n173), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(new_n169), .b(new_n176), .o1(new_n177));
  aboi22aa1n03x5               g082(.a(new_n165), .b(new_n177), .c(new_n162), .d(new_n167), .out0(\s[14] ));
  nor042aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nand22aa1n02x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n169), .c(new_n176), .out0(\s[15] ));
  nanp02aa1n02x5               g087(.a(new_n177), .b(new_n181), .o1(new_n183));
  nor042aa1n02x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand22aa1n02x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  aoib12aa1n02x5               g090(.a(new_n179), .b(new_n185), .c(new_n184), .out0(new_n186));
  nona23aa1n02x4               g091(.a(new_n144), .b(new_n140), .c(new_n137), .d(new_n143), .out0(new_n187));
  nor042aa1n02x5               g092(.a(new_n153), .b(new_n99), .o1(new_n188));
  nano23aa1d15x5               g093(.a(new_n179), .b(new_n184), .c(new_n185), .d(new_n180), .out0(new_n189));
  nona23aa1n09x5               g094(.a(new_n189), .b(new_n188), .c(new_n187), .d(new_n168), .out0(new_n190));
  oabi12aa1n18x5               g095(.a(new_n190), .b(new_n150), .c(new_n151), .out0(new_n191));
  oai012aa1n03x5               g096(.a(new_n185), .b(new_n184), .c(new_n179), .o1(new_n192));
  aobi12aa1n12x5               g097(.a(new_n192), .b(new_n175), .c(new_n189), .out0(new_n193));
  nand02aa1d12x5               g098(.a(new_n193), .b(new_n191), .o1(new_n194));
  aboi22aa1n03x5               g099(.a(new_n184), .b(new_n194), .c(new_n183), .d(new_n186), .out0(\s[16] ));
  xorc02aa1n12x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  nanb02aa1n02x5               g101(.a(new_n196), .b(new_n192), .out0(new_n197));
  aoi012aa1n02x5               g102(.a(new_n197), .b(new_n175), .c(new_n189), .o1(new_n198));
  aoi022aa1n02x5               g103(.a(new_n194), .b(new_n196), .c(new_n191), .d(new_n198), .o1(\s[17] ));
  oaoi13aa1n09x5               g104(.a(new_n190), .b(new_n130), .c(new_n112), .d(new_n122), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n168), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n201), .b(new_n157), .c(new_n152), .d(new_n156), .o1(new_n202));
  inv040aa1n03x5               g107(.a(new_n189), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n192), .b(new_n203), .c(new_n202), .d(new_n174), .o1(new_n204));
  inv040aa1d32x5               g109(.a(\a[17] ), .o1(new_n205));
  inv040aa1d28x5               g110(.a(\b[16] ), .o1(new_n206));
  nanp02aa1n02x5               g111(.a(new_n206), .b(new_n205), .o1(new_n207));
  nor042aa1n02x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand42aa1n02x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  oaib12aa1n02x5               g114(.a(new_n207), .b(new_n208), .c(new_n209), .out0(new_n210));
  oaoi13aa1n02x5               g115(.a(new_n210), .b(new_n196), .c(new_n204), .d(new_n200), .o1(new_n211));
  nano22aa1n03x7               g116(.a(new_n208), .b(new_n196), .c(new_n209), .out0(new_n212));
  oaih12aa1n02x5               g117(.a(new_n212), .b(new_n204), .c(new_n200), .o1(new_n213));
  aoai13aa1n06x5               g118(.a(new_n209), .b(new_n208), .c(new_n205), .d(new_n206), .o1(new_n214));
  aoi012aa1n02x5               g119(.a(new_n208), .b(new_n213), .c(new_n214), .o1(new_n215));
  norp02aa1n02x5               g120(.a(new_n215), .b(new_n211), .o1(\s[18] ));
  nor042aa1n06x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nanp02aa1n03x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n213), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g125(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n02x5               g126(.a(new_n217), .o1(new_n222));
  tech160nm_fioaoi03aa1n04x5   g127(.a(\a[18] ), .b(\b[17] ), .c(new_n207), .o1(new_n223));
  aoai13aa1n06x5               g128(.a(new_n219), .b(new_n223), .c(new_n194), .d(new_n212), .o1(new_n224));
  norp02aa1n06x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand02aa1n03x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  norb03aa1n02x5               g132(.a(new_n226), .b(new_n217), .c(new_n225), .out0(new_n228));
  tech160nm_finand02aa1n03p5x5 g133(.a(new_n224), .b(new_n228), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n227), .c(new_n222), .d(new_n224), .o1(\s[20] ));
  nona23aa1n03x5               g135(.a(new_n226), .b(new_n218), .c(new_n217), .d(new_n225), .out0(new_n231));
  nano23aa1n02x4               g136(.a(new_n231), .b(new_n208), .c(new_n196), .d(new_n209), .out0(new_n232));
  oaoi03aa1n02x5               g137(.a(\a[20] ), .b(\b[19] ), .c(new_n222), .o1(new_n233));
  oabi12aa1n03x5               g138(.a(new_n233), .b(new_n231), .c(new_n214), .out0(new_n234));
  nor042aa1n06x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nanp02aa1n02x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n234), .c(new_n194), .d(new_n232), .o1(new_n238));
  nano23aa1n06x5               g143(.a(new_n217), .b(new_n225), .c(new_n226), .d(new_n218), .out0(new_n239));
  aoi112aa1n02x5               g144(.a(new_n233), .b(new_n237), .c(new_n239), .d(new_n223), .o1(new_n240));
  aobi12aa1n02x5               g145(.a(new_n240), .b(new_n194), .c(new_n232), .out0(new_n241));
  norb02aa1n03x4               g146(.a(new_n238), .b(new_n241), .out0(\s[21] ));
  inv000aa1n06x5               g147(.a(new_n235), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[21] ), .b(\a[22] ), .out0(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  and002aa1n02x5               g150(.a(\b[21] ), .b(\a[22] ), .o(new_n246));
  oai022aa1n02x5               g151(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n247));
  nona22aa1n02x5               g152(.a(new_n238), .b(new_n246), .c(new_n247), .out0(new_n248));
  aoai13aa1n03x5               g153(.a(new_n248), .b(new_n245), .c(new_n243), .d(new_n238), .o1(\s[22] ));
  nano22aa1n12x5               g154(.a(new_n244), .b(new_n243), .c(new_n236), .out0(new_n250));
  nand23aa1n04x5               g155(.a(new_n212), .b(new_n250), .c(new_n239), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n250), .b(new_n233), .c(new_n239), .d(new_n223), .o1(new_n253));
  oaoi03aa1n02x5               g158(.a(\a[22] ), .b(\b[21] ), .c(new_n243), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  nanp02aa1n02x5               g160(.a(new_n253), .b(new_n255), .o1(new_n256));
  xnrc02aa1n12x5               g161(.a(\b[22] ), .b(\a[23] ), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n256), .c(new_n194), .d(new_n252), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(new_n258), .b(new_n256), .c(new_n194), .d(new_n252), .o1(new_n260));
  norb02aa1n03x4               g165(.a(new_n259), .b(new_n260), .out0(\s[23] ));
  norp02aa1n02x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .out0(new_n264));
  and002aa1n02x5               g169(.a(\b[23] ), .b(\a[24] ), .o(new_n265));
  oai022aa1n02x5               g170(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n266));
  nona22aa1n03x5               g171(.a(new_n259), .b(new_n265), .c(new_n266), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n264), .c(new_n263), .d(new_n259), .o1(\s[24] ));
  norb02aa1n02x5               g173(.a(new_n264), .b(new_n257), .out0(new_n269));
  inv020aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  nano32aa1n02x4               g175(.a(new_n270), .b(new_n212), .c(new_n250), .d(new_n239), .out0(new_n271));
  aob012aa1n02x5               g176(.a(new_n266), .b(\b[23] ), .c(\a[24] ), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n270), .c(new_n253), .d(new_n255), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n194), .d(new_n271), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(new_n274), .b(new_n273), .c(new_n194), .d(new_n271), .o1(new_n276));
  norb02aa1n03x4               g181(.a(new_n275), .b(new_n276), .out0(\s[25] ));
  norp02aa1n02x5               g182(.a(\b[24] ), .b(\a[25] ), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  tech160nm_fixorc02aa1n03p5x5 g184(.a(\a[26] ), .b(\b[25] ), .out0(new_n280));
  and002aa1n02x5               g185(.a(\b[25] ), .b(\a[26] ), .o(new_n281));
  oai022aa1n02x5               g186(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n282));
  nona22aa1n02x5               g187(.a(new_n275), .b(new_n281), .c(new_n282), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n280), .c(new_n279), .d(new_n275), .o1(\s[26] ));
  and002aa1n06x5               g189(.a(new_n280), .b(new_n274), .o(new_n285));
  nano22aa1n09x5               g190(.a(new_n251), .b(new_n285), .c(new_n269), .out0(new_n286));
  tech160nm_fioai012aa1n04x5   g191(.a(new_n286), .b(new_n204), .c(new_n200), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n281), .o1(new_n288));
  aoi022aa1n02x7               g193(.a(new_n273), .b(new_n285), .c(new_n288), .d(new_n282), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[27] ), .b(\b[26] ), .out0(new_n290));
  xnbna2aa1n03x5               g195(.a(new_n290), .b(new_n287), .c(new_n289), .out0(\s[27] ));
  nor042aa1n03x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  inv040aa1n03x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n269), .b(new_n254), .c(new_n234), .d(new_n250), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n285), .o1(new_n295));
  aob012aa1n02x5               g200(.a(new_n282), .b(\b[25] ), .c(\a[26] ), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n295), .c(new_n294), .d(new_n272), .o1(new_n297));
  aoai13aa1n06x5               g202(.a(new_n290), .b(new_n297), .c(new_n194), .d(new_n286), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  oai022aa1n02x5               g204(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n300));
  aoi012aa1n02x5               g205(.a(new_n300), .b(\a[28] ), .c(\b[27] ), .o1(new_n301));
  tech160nm_finand02aa1n03p5x5 g206(.a(new_n298), .b(new_n301), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n299), .c(new_n293), .d(new_n298), .o1(\s[28] ));
  xorc02aa1n12x5               g208(.a(\a[29] ), .b(\b[28] ), .out0(new_n304));
  and002aa1n02x5               g209(.a(new_n299), .b(new_n290), .o(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n297), .c(new_n194), .d(new_n286), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n304), .o1(new_n307));
  oaoi03aa1n09x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n293), .o1(new_n308));
  nona22aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n308), .out0(new_n309));
  inv000aa1n06x5               g214(.a(new_n286), .o1(new_n310));
  aoi012aa1n06x5               g215(.a(new_n310), .b(new_n193), .c(new_n191), .o1(new_n311));
  oaoi13aa1n02x7               g216(.a(new_n308), .b(new_n305), .c(new_n311), .d(new_n297), .o1(new_n312));
  oai012aa1n03x5               g217(.a(new_n309), .b(new_n312), .c(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g219(.a(new_n307), .b(new_n290), .c(new_n299), .out0(new_n315));
  inv000aa1n03x5               g220(.a(new_n308), .o1(new_n316));
  oaoi03aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .o1(new_n317));
  oaoi13aa1n03x5               g222(.a(new_n317), .b(new_n315), .c(new_n311), .d(new_n297), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  inv000aa1d42x5               g224(.a(new_n315), .o1(new_n320));
  norb02aa1n02x5               g225(.a(new_n319), .b(new_n317), .out0(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n320), .c(new_n287), .d(new_n289), .o1(new_n322));
  oai012aa1n03x5               g227(.a(new_n322), .b(new_n318), .c(new_n319), .o1(\s[30] ));
  nano32aa1n06x5               g228(.a(new_n307), .b(new_n319), .c(new_n290), .d(new_n299), .out0(new_n324));
  inv000aa1d42x5               g229(.a(new_n324), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\a[30] ), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\b[29] ), .o1(new_n327));
  oaoi03aa1n12x5               g232(.a(new_n326), .b(new_n327), .c(new_n317), .o1(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n325), .c(new_n287), .d(new_n289), .o1(new_n329));
  xnrc02aa1n02x5               g234(.a(\b[30] ), .b(\a[31] ), .out0(new_n330));
  nand02aa1n02x5               g235(.a(new_n329), .b(new_n330), .o1(new_n331));
  aoai13aa1n03x5               g236(.a(new_n324), .b(new_n297), .c(new_n194), .d(new_n286), .o1(new_n332));
  inv000aa1d42x5               g237(.a(new_n328), .o1(new_n333));
  nona22aa1n03x5               g238(.a(new_n332), .b(new_n333), .c(new_n330), .out0(new_n334));
  nanp02aa1n03x5               g239(.a(new_n331), .b(new_n334), .o1(\s[31] ));
  norb02aa1n02x5               g240(.a(new_n108), .b(new_n107), .out0(new_n336));
  xobna2aa1n03x5               g241(.a(new_n336), .b(new_n106), .c(new_n104), .out0(\s[3] ));
  aoi012aa1n02x5               g242(.a(new_n107), .b(new_n109), .c(new_n106), .o1(new_n338));
  xnrc02aa1n02x5               g243(.a(new_n338), .b(new_n102), .out0(\s[4] ));
  aoi112aa1n02x5               g244(.a(new_n121), .b(new_n100), .c(new_n101), .d(new_n107), .o1(new_n340));
  aboi22aa1n03x5               g245(.a(new_n112), .b(new_n121), .c(new_n340), .d(new_n149), .out0(\s[5] ));
  aob012aa1n02x5               g246(.a(new_n121), .b(new_n149), .c(new_n110), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n120), .b(new_n342), .c(new_n123), .out0(\s[6] ));
  nanb02aa1n02x5               g248(.a(new_n124), .b(new_n342), .out0(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n127), .b(new_n344), .c(new_n119), .out0(\s[7] ));
  aoi013aa1n02x4               g250(.a(new_n115), .b(new_n344), .c(new_n119), .d(new_n116), .o1(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n126), .c(new_n114), .out0(\s[8] ));
  xorb03aa1n02x5               g252(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


