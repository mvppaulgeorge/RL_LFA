// Benchmark "adder" written by ABC on Wed Jul 17 20:42:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n325, new_n327, new_n328, new_n329, new_n330, new_n333,
    new_n335, new_n337, new_n338, new_n339, new_n340;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[5] ), .b(\a[6] ), .o1(new_n99));
  norp02aa1n02x5               g004(.a(\b[5] ), .b(\a[6] ), .o1(new_n100));
  norp02aa1n02x5               g005(.a(\b[4] ), .b(\a[5] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[4] ), .b(\a[5] ), .o1(new_n102));
  nano23aa1n02x4               g007(.a(new_n101), .b(new_n100), .c(new_n102), .d(new_n99), .out0(new_n103));
  norp02aa1n02x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  nand42aa1n03x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nano23aa1n02x4               g012(.a(new_n104), .b(new_n106), .c(new_n107), .d(new_n105), .out0(new_n108));
  nand42aa1n02x5               g013(.a(new_n108), .b(new_n103), .o1(new_n109));
  nand42aa1n04x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  norp02aa1n02x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nano22aa1n02x4               g018(.a(new_n112), .b(new_n111), .c(new_n113), .out0(new_n114));
  nanp02aa1n02x5               g019(.a(\b[0] ), .b(\a[1] ), .o1(new_n115));
  norp02aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nona22aa1n02x4               g021(.a(new_n111), .b(new_n116), .c(new_n115), .out0(new_n117));
  orn002aa1n12x5               g022(.a(\a[4] ), .b(\b[3] ), .o(new_n118));
  oai112aa1n06x5               g023(.a(new_n118), .b(new_n110), .c(\b[2] ), .d(\a[3] ), .o1(new_n119));
  aoai13aa1n04x5               g024(.a(new_n110), .b(new_n119), .c(new_n114), .d(new_n117), .o1(new_n120));
  oai012aa1n02x5               g025(.a(new_n105), .b(new_n106), .c(new_n104), .o1(new_n121));
  oa0012aa1n02x5               g026(.a(new_n99), .b(new_n100), .c(new_n101), .o(new_n122));
  aobi12aa1n06x5               g027(.a(new_n121), .b(new_n108), .c(new_n122), .out0(new_n123));
  tech160nm_fioai012aa1n05x5   g028(.a(new_n123), .b(new_n120), .c(new_n109), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nanp03aa1n02x5               g030(.a(new_n124), .b(new_n98), .c(new_n125), .o1(new_n126));
  norp02aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nona23aa1n02x4               g034(.a(new_n126), .b(new_n128), .c(new_n127), .d(new_n97), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .d(new_n126), .o1(\s[10] ));
  nano23aa1n09x5               g036(.a(new_n97), .b(new_n127), .c(new_n128), .d(new_n125), .out0(new_n132));
  tech160nm_fioaoi03aa1n03p5x5 g037(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n133));
  tech160nm_fiaoi012aa1n04x5   g038(.a(new_n133), .b(new_n124), .c(new_n132), .o1(new_n134));
  nor002aa1n06x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv000aa1n02x5               g040(.a(new_n135), .o1(new_n136));
  nand42aa1n02x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n134), .b(new_n137), .c(new_n136), .out0(\s[11] ));
  nanb02aa1n02x5               g043(.a(new_n135), .b(new_n137), .out0(new_n139));
  oab012aa1n02x4               g044(.a(new_n135), .b(new_n134), .c(new_n139), .out0(new_n140));
  orn002aa1n02x5               g045(.a(\a[12] ), .b(\b[11] ), .o(new_n141));
  nanp02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nor002aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nona22aa1n02x4               g048(.a(new_n142), .b(new_n143), .c(new_n135), .out0(new_n144));
  oabi12aa1n02x5               g049(.a(new_n144), .b(new_n134), .c(new_n139), .out0(new_n145));
  aoai13aa1n02x5               g050(.a(new_n145), .b(new_n140), .c(new_n142), .d(new_n141), .o1(\s[12] ));
  nano23aa1n06x5               g051(.a(new_n135), .b(new_n143), .c(new_n142), .d(new_n137), .out0(new_n147));
  nanp02aa1n02x5               g052(.a(new_n147), .b(new_n132), .o1(new_n148));
  oaoi03aa1n02x5               g053(.a(\a[12] ), .b(\b[11] ), .c(new_n136), .o1(new_n149));
  aoi012aa1n02x5               g054(.a(new_n149), .b(new_n147), .c(new_n133), .o1(new_n150));
  oaib12aa1n03x5               g055(.a(new_n150), .b(new_n148), .c(new_n124), .out0(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  tech160nm_fixnrc02aa1n04x5   g057(.a(\b[12] ), .b(\a[13] ), .out0(new_n153));
  norb02aa1n02x5               g058(.a(new_n151), .b(new_n153), .out0(new_n154));
  norp02aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  aoib12aa1n02x5               g060(.a(new_n155), .b(new_n151), .c(new_n153), .out0(new_n156));
  tech160nm_fixnrc02aa1n04x5   g061(.a(\b[13] ), .b(\a[14] ), .out0(new_n157));
  nanp02aa1n02x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  oai022aa1n02x5               g063(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n159));
  nanb02aa1n02x5               g064(.a(new_n159), .b(new_n158), .out0(new_n160));
  obai22aa1n02x7               g065(.a(new_n157), .b(new_n156), .c(new_n154), .d(new_n160), .out0(\s[14] ));
  nor042aa1n02x5               g066(.a(new_n157), .b(new_n153), .o1(new_n162));
  aboi22aa1n03x5               g067(.a(new_n150), .b(new_n162), .c(new_n158), .d(new_n159), .out0(new_n163));
  nona32aa1n02x4               g068(.a(new_n124), .b(new_n157), .c(new_n153), .d(new_n148), .out0(new_n164));
  nor002aa1d32x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanp02aa1n04x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n164), .c(new_n163), .out0(\s[15] ));
  inv000aa1d42x5               g073(.a(new_n165), .o1(new_n169));
  aob012aa1n02x5               g074(.a(new_n167), .b(new_n164), .c(new_n163), .out0(new_n170));
  nor022aa1n12x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nand42aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  nona23aa1n02x4               g078(.a(new_n170), .b(new_n172), .c(new_n171), .d(new_n165), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n173), .c(new_n169), .d(new_n170), .o1(\s[16] ));
  nona23aa1n06x5               g080(.a(new_n142), .b(new_n137), .c(new_n135), .d(new_n143), .out0(new_n176));
  nona23aa1d16x5               g081(.a(new_n172), .b(new_n166), .c(new_n165), .d(new_n171), .out0(new_n177));
  nona23aa1d18x5               g082(.a(new_n162), .b(new_n132), .c(new_n177), .d(new_n176), .out0(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  nand02aa1d04x5               g084(.a(new_n124), .b(new_n179), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n172), .b(new_n171), .c(new_n165), .o1(new_n181));
  aoai13aa1n04x5               g086(.a(new_n162), .b(new_n149), .c(new_n147), .d(new_n133), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(new_n159), .b(new_n158), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n177), .o1(new_n184));
  aob012aa1n02x5               g089(.a(new_n184), .b(new_n182), .c(new_n183), .out0(new_n185));
  nand23aa1n06x5               g090(.a(new_n180), .b(new_n185), .c(new_n181), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  inv040aa1n08x5               g093(.a(new_n188), .o1(new_n189));
  oaoi13aa1n12x5               g094(.a(new_n178), .b(new_n123), .c(new_n120), .d(new_n109), .o1(new_n190));
  aoai13aa1n06x5               g095(.a(new_n181), .b(new_n177), .c(new_n182), .d(new_n183), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  oai012aa1n02x5               g097(.a(new_n192), .b(new_n191), .c(new_n190), .o1(new_n193));
  xorc02aa1n02x5               g098(.a(\a[18] ), .b(\b[17] ), .out0(new_n194));
  inv000aa1d42x5               g099(.a(\a[18] ), .o1(new_n195));
  inv000aa1d42x5               g100(.a(\b[17] ), .o1(new_n196));
  aoi012aa1n02x5               g101(.a(new_n188), .b(new_n195), .c(new_n196), .o1(new_n197));
  oai112aa1n02x5               g102(.a(new_n193), .b(new_n197), .c(new_n196), .d(new_n195), .o1(new_n198));
  aoai13aa1n02x5               g103(.a(new_n198), .b(new_n194), .c(new_n189), .d(new_n193), .o1(\s[18] ));
  and002aa1n02x5               g104(.a(new_n194), .b(new_n192), .o(new_n200));
  oaih12aa1n02x5               g105(.a(new_n200), .b(new_n191), .c(new_n190), .o1(new_n201));
  oaoi03aa1n12x5               g106(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  nor042aa1n09x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanp02aa1n02x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n201), .c(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g114(.a(new_n204), .o1(new_n210));
  aoai13aa1n03x5               g115(.a(new_n207), .b(new_n202), .c(new_n186), .d(new_n200), .o1(new_n211));
  nor042aa1n02x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand02aa1n16x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n213), .o1(new_n215));
  oai022aa1n02x5               g120(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n216));
  norp02aa1n02x5               g121(.a(new_n216), .b(new_n215), .o1(new_n217));
  aoai13aa1n02x5               g122(.a(new_n217), .b(new_n206), .c(new_n201), .d(new_n203), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n214), .c(new_n211), .d(new_n210), .o1(\s[20] ));
  nano23aa1n03x7               g124(.a(new_n204), .b(new_n212), .c(new_n213), .d(new_n205), .out0(new_n220));
  nand23aa1n03x5               g125(.a(new_n220), .b(new_n192), .c(new_n194), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oaih12aa1n02x5               g127(.a(new_n222), .b(new_n191), .c(new_n190), .o1(new_n223));
  aoi022aa1n02x7               g128(.a(new_n220), .b(new_n202), .c(new_n213), .d(new_n216), .o1(new_n224));
  xnrc02aa1n12x5               g129(.a(\b[20] ), .b(\a[21] ), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n224), .out0(\s[21] ));
  norp02aa1n02x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n224), .o1(new_n230));
  aoai13aa1n03x5               g135(.a(new_n226), .b(new_n230), .c(new_n186), .d(new_n222), .o1(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  nanp02aa1n02x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  oai022aa1n02x5               g139(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n234), .b(new_n235), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n225), .c(new_n223), .d(new_n224), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n233), .c(new_n231), .d(new_n229), .o1(\s[22] ));
  nor002aa1n04x5               g143(.a(new_n232), .b(new_n225), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n221), .out0(new_n240));
  oaih12aa1n02x5               g145(.a(new_n240), .b(new_n191), .c(new_n190), .o1(new_n241));
  oab012aa1n02x4               g146(.a(new_n215), .b(new_n204), .c(new_n212), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n239), .b(new_n242), .c(new_n220), .d(new_n202), .o1(new_n243));
  nanp02aa1n02x5               g148(.a(new_n235), .b(new_n234), .o1(new_n244));
  nanp02aa1n02x5               g149(.a(new_n243), .b(new_n244), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[22] ), .b(\a[23] ), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  xnbna2aa1n03x5               g153(.a(new_n248), .b(new_n241), .c(new_n246), .out0(\s[23] ));
  norp02aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n248), .b(new_n245), .c(new_n186), .d(new_n240), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .out0(new_n253));
  nanp02aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .o1(new_n254));
  oai022aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n254), .b(new_n255), .out0(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n247), .c(new_n241), .d(new_n246), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n253), .c(new_n252), .d(new_n251), .o1(\s[24] ));
  nano32aa1n02x5               g163(.a(new_n221), .b(new_n253), .c(new_n239), .d(new_n248), .out0(new_n259));
  oaih12aa1n02x5               g164(.a(new_n259), .b(new_n191), .c(new_n190), .o1(new_n260));
  norb02aa1n02x5               g165(.a(new_n253), .b(new_n247), .out0(new_n261));
  inv000aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(new_n255), .b(new_n254), .o1(new_n263));
  aoai13aa1n12x5               g168(.a(new_n263), .b(new_n262), .c(new_n243), .d(new_n244), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n260), .c(new_n265), .out0(\s[25] ));
  norp02aa1n02x5               g172(.a(\b[24] ), .b(\a[25] ), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  aoai13aa1n03x5               g174(.a(new_n266), .b(new_n264), .c(new_n186), .d(new_n259), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[26] ), .b(\b[25] ), .out0(new_n271));
  inv000aa1d42x5               g176(.a(new_n266), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .o1(new_n273));
  oai022aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n274));
  norb02aa1n02x5               g179(.a(new_n273), .b(new_n274), .out0(new_n275));
  aoai13aa1n02x5               g180(.a(new_n275), .b(new_n272), .c(new_n260), .d(new_n265), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n271), .c(new_n270), .d(new_n269), .o1(\s[26] ));
  and002aa1n02x5               g182(.a(new_n271), .b(new_n266), .o(new_n278));
  nano32aa1n06x5               g183(.a(new_n221), .b(new_n278), .c(new_n239), .d(new_n261), .out0(new_n279));
  oai012aa1n12x5               g184(.a(new_n279), .b(new_n191), .c(new_n190), .o1(new_n280));
  aoi022aa1d18x5               g185(.a(new_n264), .b(new_n278), .c(new_n273), .d(new_n274), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n06x5               g187(.a(new_n282), .b(new_n280), .c(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  nanp02aa1n03x5               g190(.a(new_n264), .b(new_n278), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(new_n274), .b(new_n273), .o1(new_n287));
  nanp02aa1n03x5               g192(.a(new_n286), .b(new_n287), .o1(new_n288));
  aoai13aa1n02x5               g193(.a(new_n282), .b(new_n288), .c(new_n186), .d(new_n279), .o1(new_n289));
  xorc02aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n282), .o1(new_n291));
  oai022aa1n02x5               g196(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n292));
  aoi012aa1n02x5               g197(.a(new_n292), .b(\a[28] ), .c(\b[27] ), .o1(new_n293));
  aoai13aa1n02x7               g198(.a(new_n293), .b(new_n291), .c(new_n280), .d(new_n281), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n290), .c(new_n289), .d(new_n285), .o1(\s[28] ));
  and002aa1n02x5               g200(.a(new_n290), .b(new_n282), .o(new_n296));
  inv000aa1d42x5               g201(.a(new_n296), .o1(new_n297));
  aob012aa1n02x5               g202(.a(new_n292), .b(\b[27] ), .c(\a[28] ), .out0(new_n298));
  xorc02aa1n12x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  and002aa1n02x5               g204(.a(new_n299), .b(new_n298), .o(new_n300));
  aoai13aa1n02x5               g205(.a(new_n300), .b(new_n297), .c(new_n280), .d(new_n281), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n299), .o1(new_n302));
  aoai13aa1n06x5               g207(.a(new_n298), .b(new_n297), .c(new_n280), .d(new_n281), .o1(new_n303));
  nanp02aa1n03x5               g208(.a(new_n303), .b(new_n302), .o1(new_n304));
  nanp02aa1n03x5               g209(.a(new_n304), .b(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n115), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g211(.a(new_n290), .b(new_n282), .c(new_n299), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n308));
  aoai13aa1n06x5               g213(.a(new_n308), .b(new_n307), .c(new_n280), .d(new_n281), .o1(new_n309));
  xorc02aa1n12x5               g214(.a(\a[30] ), .b(\b[29] ), .out0(new_n310));
  inv000aa1d42x5               g215(.a(new_n310), .o1(new_n311));
  nanp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(new_n312));
  norb02aa1n02x5               g217(.a(new_n308), .b(new_n311), .out0(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n307), .c(new_n280), .d(new_n281), .o1(new_n314));
  nanp02aa1n03x5               g219(.a(new_n312), .b(new_n314), .o1(\s[30] ));
  nano32aa1n03x7               g220(.a(new_n291), .b(new_n310), .c(new_n290), .d(new_n299), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n288), .c(new_n186), .d(new_n279), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[31] ), .b(\b[30] ), .out0(new_n318));
  inv000aa1d42x5               g223(.a(new_n316), .o1(new_n319));
  oai012aa1n02x5               g224(.a(new_n318), .b(\b[29] ), .c(\a[30] ), .o1(new_n320));
  oab012aa1n02x4               g225(.a(new_n320), .b(new_n308), .c(new_n311), .out0(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n319), .c(new_n280), .d(new_n281), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n323));
  aoai13aa1n03x5               g228(.a(new_n322), .b(new_n318), .c(new_n317), .d(new_n323), .o1(\s[31] ));
  norb02aa1n02x5               g229(.a(new_n113), .b(new_n112), .out0(new_n325));
  xobna2aa1n03x5               g230(.a(new_n325), .b(new_n117), .c(new_n111), .out0(\s[3] ));
  oai112aa1n02x5               g231(.a(new_n325), .b(new_n111), .c(new_n115), .d(new_n116), .o1(new_n327));
  inv000aa1d42x5               g232(.a(new_n119), .o1(new_n328));
  nanp02aa1n02x5               g233(.a(new_n327), .b(new_n328), .o1(new_n329));
  aoi012aa1n02x5               g234(.a(new_n112), .b(new_n114), .c(new_n117), .o1(new_n330));
  aoai13aa1n02x5               g235(.a(new_n329), .b(new_n330), .c(new_n118), .d(new_n110), .o1(\s[4] ));
  xnrb03aa1n02x5               g236(.a(new_n120), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi013aa1n02x4               g237(.a(new_n101), .b(new_n329), .c(new_n110), .d(new_n102), .o1(new_n333));
  xnrb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g239(.a(\a[6] ), .b(\b[5] ), .c(new_n333), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  norb02aa1n02x5               g241(.a(new_n107), .b(new_n106), .out0(new_n337));
  nona22aa1n02x4               g242(.a(new_n105), .b(new_n106), .c(new_n104), .out0(new_n338));
  nanb02aa1n02x5               g243(.a(new_n104), .b(new_n105), .out0(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n106), .c(new_n335), .d(new_n107), .o1(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n338), .c(new_n337), .d(new_n335), .o1(\s[8] ));
  xorb03aa1n02x5               g246(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


