// Benchmark "adder" written by ABC on Thu Jul 18 12:00:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n306,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n324, new_n326, new_n327, new_n328, new_n330, new_n331, new_n332,
    new_n334, new_n335, new_n336, new_n338, new_n339, new_n340, new_n342,
    new_n343, new_n344, new_n345, new_n347, new_n348, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  oa0022aa1n06x5               g002(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n98));
  oai112aa1n06x5               g003(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n99));
  inv040aa1d32x5               g004(.a(\a[3] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[2] ), .o1(new_n101));
  nand02aa1n06x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nand42aa1n04x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand23aa1n06x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  oaib12aa1n18x5               g010(.a(new_n98), .b(new_n105), .c(new_n99), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\a[8] ), .o1(new_n107));
  inv040aa1d32x5               g012(.a(\b[7] ), .o1(new_n108));
  nand42aa1d28x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  inv040aa1d32x5               g014(.a(\a[5] ), .o1(new_n110));
  inv000aa1d48x5               g015(.a(\b[4] ), .o1(new_n111));
  nand02aa1n10x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  oai112aa1n04x5               g017(.a(new_n112), .b(new_n109), .c(new_n108), .d(new_n107), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  inv040aa1d32x5               g019(.a(\a[7] ), .o1(new_n115));
  inv040aa1d32x5               g020(.a(\b[6] ), .o1(new_n116));
  nand02aa1d16x5               g021(.a(new_n116), .b(new_n115), .o1(new_n117));
  nand22aa1n12x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand03aa1n02x5               g023(.a(new_n117), .b(new_n114), .c(new_n118), .o1(new_n119));
  nand42aa1n16x5               g024(.a(\b[3] ), .b(\a[4] ), .o1(new_n120));
  oai122aa1n06x5               g025(.a(new_n120), .b(\a[8] ), .c(\b[7] ), .d(\a[6] ), .e(\b[5] ), .o1(new_n121));
  nor043aa1n06x5               g026(.a(new_n113), .b(new_n119), .c(new_n121), .o1(new_n122));
  and002aa1n06x5               g027(.a(\b[7] ), .b(\a[8] ), .o(new_n123));
  nanp02aa1n02x5               g028(.a(new_n108), .b(new_n107), .o1(new_n124));
  oai022aa1d18x5               g029(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n125));
  nanp03aa1n03x5               g030(.a(new_n125), .b(new_n114), .c(new_n118), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n124), .b(new_n123), .c(new_n126), .d(new_n117), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n127), .c(new_n106), .d(new_n122), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n97), .out0(\s[10] ));
  nanp02aa1n02x5               g036(.a(new_n129), .b(new_n97), .o1(new_n132));
  oaoi03aa1n09x5               g037(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n133));
  nor022aa1n16x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  aoai13aa1n06x5               g041(.a(new_n136), .b(new_n133), .c(new_n132), .d(new_n130), .o1(new_n137));
  aoi112aa1n02x5               g042(.a(new_n136), .b(new_n133), .c(new_n132), .d(new_n130), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(\s[11] ));
  orn002aa1n24x5               g044(.a(\a[11] ), .b(\b[10] ), .o(new_n140));
  nor022aa1n16x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanp02aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  nona23aa1n02x4               g048(.a(new_n137), .b(new_n142), .c(new_n141), .d(new_n134), .out0(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n143), .c(new_n140), .d(new_n137), .o1(\s[12] ));
  nona23aa1n09x5               g050(.a(new_n142), .b(new_n135), .c(new_n134), .d(new_n141), .out0(new_n146));
  nano22aa1n03x7               g051(.a(new_n146), .b(new_n128), .c(new_n130), .out0(new_n147));
  aoai13aa1n03x5               g052(.a(new_n147), .b(new_n127), .c(new_n106), .d(new_n122), .o1(new_n148));
  oai022aa1n02x7               g053(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n149));
  aob012aa1n03x5               g054(.a(new_n149), .b(\b[9] ), .c(\a[10] ), .out0(new_n150));
  oaoi03aa1n09x5               g055(.a(\a[12] ), .b(\b[11] ), .c(new_n140), .o1(new_n151));
  oabi12aa1n06x5               g056(.a(new_n151), .b(new_n146), .c(new_n150), .out0(new_n152));
  nanb02aa1n06x5               g057(.a(new_n152), .b(new_n148), .out0(new_n153));
  nor002aa1d32x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nanp02aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  norb02aa1n06x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  nano23aa1n03x5               g061(.a(new_n134), .b(new_n141), .c(new_n142), .d(new_n135), .out0(new_n157));
  aoi112aa1n02x5               g062(.a(new_n151), .b(new_n156), .c(new_n157), .d(new_n133), .o1(new_n158));
  aoi022aa1n02x5               g063(.a(new_n153), .b(new_n156), .c(new_n148), .d(new_n158), .o1(\s[13] ));
  xnrc02aa1n02x5               g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n154), .c(new_n153), .d(new_n156), .o1(new_n161));
  inv000aa1d42x5               g066(.a(\b[13] ), .o1(new_n162));
  inv000aa1d42x5               g067(.a(\a[14] ), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n154), .b(new_n163), .c(new_n162), .o1(new_n164));
  oaib12aa1n02x5               g069(.a(new_n164), .b(new_n162), .c(\a[14] ), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n161), .b(new_n165), .c(new_n156), .d(new_n153), .o1(\s[14] ));
  inv030aa1n06x5               g071(.a(new_n154), .o1(new_n167));
  nano22aa1n03x7               g072(.a(new_n160), .b(new_n167), .c(new_n155), .out0(new_n168));
  oaoi03aa1n09x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n169));
  xorc02aa1n12x5               g074(.a(\a[15] ), .b(\b[14] ), .out0(new_n170));
  aoai13aa1n04x5               g075(.a(new_n170), .b(new_n169), .c(new_n153), .d(new_n168), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n170), .b(new_n169), .c(new_n153), .d(new_n168), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[15] ));
  nor002aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  nor042aa1n06x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nand02aa1n16x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  norb02aa1n03x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  nona23aa1n03x5               g083(.a(new_n171), .b(new_n177), .c(new_n176), .d(new_n174), .out0(new_n179));
  aoai13aa1n02x5               g084(.a(new_n179), .b(new_n178), .c(new_n175), .d(new_n171), .o1(\s[16] ));
  tech160nm_fiaoi012aa1n05x5   g085(.a(new_n127), .b(new_n106), .c(new_n122), .o1(new_n181));
  tech160nm_fixorc02aa1n02p5x5 g086(.a(\a[14] ), .b(\b[13] ), .out0(new_n182));
  nand22aa1n03x5               g087(.a(new_n170), .b(new_n178), .o1(new_n183));
  nano22aa1n02x4               g088(.a(new_n183), .b(new_n156), .c(new_n182), .out0(new_n184));
  nand02aa1n02x5               g089(.a(new_n184), .b(new_n147), .o1(new_n185));
  inv000aa1n02x5               g090(.a(new_n183), .o1(new_n186));
  aoai13aa1n04x5               g091(.a(new_n186), .b(new_n169), .c(new_n152), .d(new_n168), .o1(new_n187));
  tech160nm_fiaoi012aa1n05x5   g092(.a(new_n176), .b(new_n174), .c(new_n177), .o1(new_n188));
  oai112aa1n06x5               g093(.a(new_n187), .b(new_n188), .c(new_n181), .d(new_n185), .o1(new_n189));
  nor042aa1n06x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nand42aa1n08x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  norb02aa1n02x7               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  norp02aa1n02x5               g097(.a(new_n181), .b(new_n185), .o1(new_n193));
  nano23aa1n02x4               g098(.a(new_n192), .b(new_n193), .c(new_n187), .d(new_n188), .out0(new_n194));
  aoi012aa1n02x5               g099(.a(new_n194), .b(new_n189), .c(new_n192), .o1(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[17] ), .o1(new_n197));
  nand42aa1n08x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  nand02aa1n04x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  aoi122aa1n02x7               g104(.a(new_n190), .b(new_n198), .c(new_n199), .d(new_n189), .e(new_n192), .o1(new_n200));
  tech160nm_fiao0012aa1n02p5x5 g105(.a(new_n190), .b(new_n189), .c(new_n191), .o(new_n201));
  aoi013aa1n02x5               g106(.a(new_n200), .b(new_n201), .c(new_n198), .d(new_n199), .o1(\s[18] ));
  nano32aa1n02x4               g107(.a(new_n190), .b(new_n199), .c(new_n191), .d(new_n198), .out0(new_n203));
  aob012aa1d15x5               g108(.a(new_n198), .b(new_n190), .c(new_n199), .out0(new_n204));
  nor042aa1n06x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanp02aa1n02x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  aoai13aa1n04x5               g112(.a(new_n207), .b(new_n204), .c(new_n189), .d(new_n203), .o1(new_n208));
  aoi112aa1n02x7               g113(.a(new_n207), .b(new_n204), .c(new_n189), .d(new_n203), .o1(new_n209));
  norb02aa1n03x4               g114(.a(new_n208), .b(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g116(.a(new_n205), .o1(new_n212));
  norp02aa1n04x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1n03x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  norb03aa1n02x5               g120(.a(new_n214), .b(new_n205), .c(new_n213), .out0(new_n216));
  nanp02aa1n03x5               g121(.a(new_n208), .b(new_n216), .o1(new_n217));
  aoai13aa1n03x5               g122(.a(new_n217), .b(new_n215), .c(new_n212), .d(new_n208), .o1(\s[20] ));
  nona23aa1n09x5               g123(.a(new_n214), .b(new_n206), .c(new_n205), .d(new_n213), .out0(new_n219));
  nano32aa1n03x7               g124(.a(new_n219), .b(new_n192), .c(new_n198), .d(new_n199), .out0(new_n220));
  oaoi03aa1n02x5               g125(.a(new_n196), .b(new_n197), .c(new_n190), .o1(new_n221));
  oaoi03aa1n06x5               g126(.a(\a[20] ), .b(\b[19] ), .c(new_n212), .o1(new_n222));
  oabi12aa1n06x5               g127(.a(new_n222), .b(new_n219), .c(new_n221), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[21] ), .b(\b[20] ), .out0(new_n224));
  aoai13aa1n04x5               g129(.a(new_n224), .b(new_n223), .c(new_n189), .d(new_n220), .o1(new_n225));
  nano23aa1n06x5               g130(.a(new_n205), .b(new_n213), .c(new_n214), .d(new_n206), .out0(new_n226));
  orn002aa1n02x5               g131(.a(new_n222), .b(new_n224), .o(new_n227));
  aoi122aa1n06x5               g132(.a(new_n227), .b(new_n204), .c(new_n226), .d(new_n189), .e(new_n220), .o1(new_n228));
  norb02aa1n03x4               g133(.a(new_n225), .b(new_n228), .out0(\s[21] ));
  nor042aa1n03x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  inv040aa1n03x5               g135(.a(new_n230), .o1(new_n231));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  and002aa1n02x5               g137(.a(\b[21] ), .b(\a[22] ), .o(new_n233));
  oai022aa1n02x5               g138(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n234));
  nona22aa1n03x5               g139(.a(new_n225), .b(new_n233), .c(new_n234), .out0(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n232), .c(new_n231), .d(new_n225), .o1(\s[22] ));
  nanp02aa1n02x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  xnrc02aa1n02x5               g142(.a(\b[21] ), .b(\a[22] ), .out0(new_n238));
  nano22aa1n03x7               g143(.a(new_n238), .b(new_n231), .c(new_n237), .out0(new_n239));
  and003aa1n02x5               g144(.a(new_n203), .b(new_n239), .c(new_n226), .o(new_n240));
  aoai13aa1n06x5               g145(.a(new_n239), .b(new_n222), .c(new_n226), .d(new_n204), .o1(new_n241));
  oao003aa1n06x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n231), .carry(new_n242));
  nanp02aa1n02x5               g147(.a(new_n241), .b(new_n242), .o1(new_n243));
  tech160nm_fixorc02aa1n03p5x5 g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  aoai13aa1n04x5               g149(.a(new_n244), .b(new_n243), .c(new_n189), .d(new_n240), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n169), .o1(new_n246));
  aoai13aa1n02x5               g151(.a(new_n168), .b(new_n151), .c(new_n157), .d(new_n133), .o1(new_n247));
  aoai13aa1n03x5               g152(.a(new_n188), .b(new_n183), .c(new_n247), .d(new_n246), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n242), .o1(new_n249));
  nona22aa1n02x4               g154(.a(new_n241), .b(new_n249), .c(new_n244), .out0(new_n250));
  oaoi13aa1n02x5               g155(.a(new_n250), .b(new_n240), .c(new_n248), .d(new_n193), .o1(new_n251));
  norb02aa1n03x4               g156(.a(new_n245), .b(new_n251), .out0(\s[23] ));
  nor042aa1n03x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[24] ), .b(\b[23] ), .out0(new_n255));
  and002aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o(new_n256));
  oai022aa1n02x5               g161(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n257));
  nona22aa1n03x5               g162(.a(new_n245), .b(new_n256), .c(new_n257), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n255), .c(new_n254), .d(new_n245), .o1(\s[24] ));
  and002aa1n06x5               g164(.a(new_n255), .b(new_n244), .o(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  nano32aa1n02x5               g166(.a(new_n261), .b(new_n239), .c(new_n203), .d(new_n226), .out0(new_n262));
  oao003aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n254), .carry(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n261), .c(new_n241), .d(new_n242), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[25] ), .b(\b[24] ), .out0(new_n265));
  aoai13aa1n04x5               g170(.a(new_n265), .b(new_n264), .c(new_n189), .d(new_n262), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n260), .b(new_n249), .c(new_n223), .d(new_n239), .o1(new_n267));
  nanb03aa1n02x5               g172(.a(new_n265), .b(new_n267), .c(new_n263), .out0(new_n268));
  aoi012aa1n02x5               g173(.a(new_n268), .b(new_n189), .c(new_n262), .o1(new_n269));
  norb02aa1n03x4               g174(.a(new_n266), .b(new_n269), .out0(\s[25] ));
  nor042aa1n03x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  tech160nm_fixorc02aa1n05x5   g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  and002aa1n02x5               g178(.a(\b[25] ), .b(\a[26] ), .o(new_n274));
  oai022aa1n02x5               g179(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n275));
  nona22aa1n03x5               g180(.a(new_n266), .b(new_n274), .c(new_n275), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n273), .c(new_n272), .d(new_n266), .o1(\s[26] ));
  and002aa1n02x5               g182(.a(new_n273), .b(new_n265), .o(new_n278));
  inv000aa1n02x5               g183(.a(new_n278), .o1(new_n279));
  nano32aa1n03x7               g184(.a(new_n279), .b(new_n220), .c(new_n260), .d(new_n239), .out0(new_n280));
  oai012aa1n06x5               g185(.a(new_n280), .b(new_n248), .c(new_n193), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[26] ), .b(\b[25] ), .c(new_n272), .carry(new_n282));
  aoai13aa1n04x5               g187(.a(new_n282), .b(new_n279), .c(new_n267), .d(new_n263), .o1(new_n283));
  xorc02aa1n12x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n283), .c(new_n189), .d(new_n280), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n282), .o1(new_n286));
  aoi112aa1n02x5               g191(.a(new_n284), .b(new_n286), .c(new_n264), .d(new_n278), .o1(new_n287));
  aobi12aa1n02x7               g192(.a(new_n285), .b(new_n287), .c(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .out0(new_n291));
  aoi012aa1n06x5               g196(.a(new_n286), .b(new_n264), .c(new_n278), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n284), .o1(new_n293));
  oai022aa1n02x5               g198(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n294));
  aoi012aa1n02x5               g199(.a(new_n294), .b(\a[28] ), .c(\b[27] ), .o1(new_n295));
  aoai13aa1n02x7               g200(.a(new_n295), .b(new_n293), .c(new_n292), .d(new_n281), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n291), .c(new_n285), .d(new_n290), .o1(\s[28] ));
  and002aa1n02x5               g202(.a(new_n291), .b(new_n284), .o(new_n298));
  aoai13aa1n02x7               g203(.a(new_n298), .b(new_n283), .c(new_n189), .d(new_n280), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n298), .o1(new_n300));
  aob012aa1n02x5               g205(.a(new_n294), .b(\b[27] ), .c(\a[28] ), .out0(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n300), .c(new_n292), .d(new_n281), .o1(new_n302));
  tech160nm_fixorc02aa1n03p5x5 g207(.a(\a[29] ), .b(\b[28] ), .out0(new_n303));
  norb02aa1n02x5               g208(.a(new_n301), .b(new_n303), .out0(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n299), .d(new_n304), .o1(\s[29] ));
  nanp02aa1n02x5               g210(.a(\b[0] ), .b(\a[1] ), .o1(new_n306));
  xorb03aa1n02x5               g211(.a(new_n306), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g212(.a(new_n293), .b(new_n291), .c(new_n303), .out0(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n283), .c(new_n189), .d(new_n280), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n308), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .carry(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n310), .c(new_n292), .d(new_n281), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n311), .b(new_n313), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[30] ));
  nano32aa1n03x7               g220(.a(new_n293), .b(new_n313), .c(new_n291), .d(new_n303), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n283), .c(new_n189), .d(new_n280), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n316), .o1(new_n318));
  oao003aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n318), .c(new_n292), .d(new_n281), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[31] ), .b(\b[30] ), .out0(new_n321));
  norb02aa1n02x5               g226(.a(new_n319), .b(new_n321), .out0(new_n322));
  aoi022aa1n03x5               g227(.a(new_n320), .b(new_n321), .c(new_n317), .d(new_n322), .o1(\s[31] ));
  nanp02aa1n02x5               g228(.a(new_n102), .b(new_n104), .o1(new_n324));
  xnbna2aa1n03x5               g229(.a(new_n324), .b(new_n99), .c(new_n103), .out0(\s[3] ));
  nano22aa1n02x4               g230(.a(new_n324), .b(new_n99), .c(new_n103), .out0(new_n326));
  xorc02aa1n02x5               g231(.a(\a[4] ), .b(\b[3] ), .out0(new_n327));
  norb02aa1n02x5               g232(.a(new_n102), .b(new_n327), .out0(new_n328));
  aboi22aa1n03x5               g233(.a(new_n326), .b(new_n328), .c(new_n106), .d(new_n327), .out0(\s[4] ));
  aoi022aa1n02x5               g234(.a(new_n106), .b(new_n120), .c(new_n109), .d(new_n112), .o1(new_n330));
  nanp03aa1n02x5               g235(.a(new_n112), .b(new_n109), .c(new_n120), .o1(new_n331));
  aoib12aa1n06x5               g236(.a(new_n331), .b(new_n98), .c(new_n326), .out0(new_n332));
  norp02aa1n02x5               g237(.a(new_n330), .b(new_n332), .o1(\s[5] ));
  xorc02aa1n02x5               g238(.a(\a[6] ), .b(\b[5] ), .out0(new_n334));
  aoai13aa1n02x5               g239(.a(new_n334), .b(new_n332), .c(new_n110), .d(new_n111), .o1(new_n335));
  aoi112aa1n02x5               g240(.a(new_n332), .b(new_n334), .c(new_n110), .d(new_n111), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n335), .b(new_n336), .out0(\s[6] ));
  xorc02aa1n02x5               g242(.a(\a[7] ), .b(\b[6] ), .out0(new_n338));
  oaoi03aa1n02x5               g243(.a(\a[6] ), .b(\b[5] ), .c(new_n112), .o1(new_n339));
  inv000aa1d42x5               g244(.a(new_n339), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n338), .b(new_n335), .c(new_n340), .out0(\s[7] ));
  aob012aa1n03x5               g246(.a(new_n338), .b(new_n335), .c(new_n340), .out0(new_n342));
  nanp02aa1n02x5               g247(.a(new_n342), .b(new_n117), .o1(new_n343));
  xorc02aa1n02x5               g248(.a(\a[8] ), .b(\b[7] ), .out0(new_n344));
  aboi22aa1n03x5               g249(.a(new_n123), .b(new_n124), .c(new_n115), .d(new_n116), .out0(new_n345));
  aoi022aa1n02x5               g250(.a(new_n343), .b(new_n344), .c(new_n342), .d(new_n345), .o1(\s[8] ));
  norb02aa1n02x5               g251(.a(new_n124), .b(new_n128), .out0(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n123), .c(new_n126), .d(new_n117), .o1(new_n348));
  aoi012aa1n02x5               g253(.a(new_n348), .b(new_n106), .c(new_n122), .o1(new_n349));
  norb02aa1n02x5               g254(.a(new_n129), .b(new_n349), .out0(\s[9] ));
endmodule


