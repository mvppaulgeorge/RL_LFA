// Benchmark "adder" written by ABC on Thu Jul 18 02:21:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n330, new_n333,
    new_n335, new_n336, new_n337, new_n339;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n03x5               g001(.a(\b[3] ), .b(\a[4] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  nor022aa1n16x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nona23aa1n06x5               g005(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n101));
  nanp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand02aa1d04x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor002aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  tech160nm_fioai012aa1n04x5   g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  aoi012aa1n02x7               g010(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n101), .c(new_n105), .o1(new_n107));
  nor022aa1n04x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nanp02aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor022aa1n16x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n09x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  nor043aa1n06x5               g019(.a(new_n112), .b(new_n113), .c(new_n114), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\a[6] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[5] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[5] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[4] ), .o1(new_n120));
  oai112aa1n04x5               g025(.a(new_n119), .b(new_n120), .c(new_n117), .d(new_n116), .o1(new_n121));
  tech160nm_fioai012aa1n03p5x5 g026(.a(new_n109), .b(new_n110), .c(new_n108), .o1(new_n122));
  aoai13aa1n06x5               g027(.a(new_n122), .b(new_n112), .c(new_n121), .d(new_n118), .o1(new_n123));
  aoi012aa1d18x5               g028(.a(new_n123), .b(new_n107), .c(new_n115), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  xorb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n09x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand22aa1n09x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nor042aa1n06x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nona23aa1n02x4               g035(.a(new_n130), .b(new_n128), .c(new_n127), .d(new_n129), .out0(new_n131));
  aoi012aa1d24x5               g036(.a(new_n127), .b(new_n129), .c(new_n128), .o1(new_n132));
  tech160nm_fioai012aa1n05x5   g037(.a(new_n132), .b(new_n124), .c(new_n131), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv040aa1n08x5               g040(.a(new_n135), .o1(new_n136));
  nand02aa1d28x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n06x5               g042(.a(new_n137), .b(new_n135), .out0(new_n138));
  nanp02aa1n02x5               g043(.a(new_n133), .b(new_n138), .o1(new_n139));
  nor002aa1n20x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand02aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n12x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n139), .c(new_n136), .out0(\s[12] ));
  nona23aa1d18x5               g048(.a(new_n141), .b(new_n137), .c(new_n135), .d(new_n140), .out0(new_n144));
  oaoi03aa1n09x5               g049(.a(\a[12] ), .b(\b[11] ), .c(new_n136), .o1(new_n145));
  inv030aa1n06x5               g050(.a(new_n145), .o1(new_n146));
  oaih12aa1n12x5               g051(.a(new_n146), .b(new_n144), .c(new_n132), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  oai013aa1n03x5               g053(.a(new_n148), .b(new_n124), .c(new_n131), .d(new_n144), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n09x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1n08x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  aoi012aa1n03x5               g057(.a(new_n151), .b(new_n149), .c(new_n152), .o1(new_n153));
  xnrb03aa1n03x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  aoi112aa1n09x5               g059(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n155));
  oai112aa1n06x5               g060(.a(new_n138), .b(new_n142), .c(new_n155), .d(new_n127), .o1(new_n156));
  nor042aa1n06x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand42aa1d28x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nano23aa1n09x5               g063(.a(new_n151), .b(new_n157), .c(new_n158), .d(new_n152), .out0(new_n159));
  inv020aa1n04x5               g064(.a(new_n159), .o1(new_n160));
  aoi012aa1d24x5               g065(.a(new_n157), .b(new_n151), .c(new_n158), .o1(new_n161));
  aoai13aa1n12x5               g066(.a(new_n161), .b(new_n160), .c(new_n156), .d(new_n146), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  inv000aa1n02x5               g068(.a(new_n124), .o1(new_n164));
  nona32aa1n02x4               g069(.a(new_n164), .b(new_n160), .c(new_n144), .d(new_n131), .out0(new_n165));
  nanp02aa1n02x5               g070(.a(new_n165), .b(new_n163), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1d28x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nanp02aa1n24x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  aoi112aa1n02x5               g077(.a(new_n168), .b(new_n172), .c(new_n166), .d(new_n169), .o1(new_n173));
  aoai13aa1n02x5               g078(.a(new_n172), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(\s[16] ));
  norb02aa1n02x5               g080(.a(new_n128), .b(new_n127), .out0(new_n176));
  norb02aa1n03x5               g081(.a(new_n130), .b(new_n129), .out0(new_n177));
  nano23aa1d15x5               g082(.a(new_n135), .b(new_n140), .c(new_n141), .d(new_n137), .out0(new_n178));
  nano23aa1d15x5               g083(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n179));
  nand02aa1d04x5               g084(.a(new_n179), .b(new_n159), .o1(new_n180));
  nano32aa1n03x7               g085(.a(new_n180), .b(new_n178), .c(new_n177), .d(new_n176), .out0(new_n181));
  aoai13aa1n12x5               g086(.a(new_n181), .b(new_n123), .c(new_n107), .d(new_n115), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n161), .o1(new_n183));
  aoai13aa1n04x5               g088(.a(new_n179), .b(new_n183), .c(new_n147), .d(new_n159), .o1(new_n184));
  oai012aa1n02x5               g089(.a(new_n171), .b(new_n170), .c(new_n168), .o1(new_n185));
  nand23aa1n06x5               g090(.a(new_n182), .b(new_n184), .c(new_n185), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nand42aa1n16x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  nor042aa1n06x5               g093(.a(\b[17] ), .b(\a[18] ), .o1(new_n189));
  nand42aa1n10x5               g094(.a(\b[17] ), .b(\a[18] ), .o1(new_n190));
  nanb02aa1n02x5               g095(.a(new_n189), .b(new_n190), .out0(new_n191));
  aobi12aa1n12x5               g096(.a(new_n185), .b(new_n162), .c(new_n179), .out0(new_n192));
  oai112aa1n02x5               g097(.a(new_n192), .b(new_n182), .c(\b[16] ), .d(\a[17] ), .o1(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n191), .b(new_n193), .c(new_n188), .out0(\s[18] ));
  nor002aa1n04x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  nano23aa1d15x5               g100(.a(new_n195), .b(new_n189), .c(new_n190), .d(new_n188), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  aoi012aa1n06x5               g102(.a(new_n189), .b(new_n195), .c(new_n190), .o1(new_n198));
  aoai13aa1n02x7               g103(.a(new_n198), .b(new_n197), .c(new_n192), .d(new_n182), .o1(new_n199));
  xorb03aa1n03x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n24x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand42aa1n06x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nor002aa1n16x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand42aa1d28x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  norb02aa1d27x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  aoi112aa1n03x4               g111(.a(new_n202), .b(new_n206), .c(new_n199), .d(new_n203), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n202), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n198), .o1(new_n209));
  norb02aa1n06x4               g114(.a(new_n203), .b(new_n202), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n209), .c(new_n186), .d(new_n196), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n206), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n212), .b(new_n211), .c(new_n208), .o1(new_n213));
  nor002aa1n02x5               g118(.a(new_n213), .b(new_n207), .o1(\s[20] ));
  nano23aa1n03x7               g119(.a(new_n202), .b(new_n204), .c(new_n205), .d(new_n203), .out0(new_n215));
  nand22aa1n09x5               g120(.a(new_n215), .b(new_n196), .o1(new_n216));
  aoi112aa1n09x5               g121(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n217));
  oai112aa1n06x5               g122(.a(new_n210), .b(new_n206), .c(new_n217), .d(new_n189), .o1(new_n218));
  oai012aa1d24x5               g123(.a(new_n205), .b(new_n204), .c(new_n202), .o1(new_n219));
  nand22aa1n12x5               g124(.a(new_n218), .b(new_n219), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n216), .c(new_n192), .d(new_n182), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  xorc02aa1n12x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoi112aa1n02x7               g132(.a(new_n224), .b(new_n227), .c(new_n222), .d(new_n225), .o1(new_n228));
  inv040aa1n08x5               g133(.a(new_n224), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n216), .o1(new_n230));
  aoai13aa1n03x5               g135(.a(new_n225), .b(new_n220), .c(new_n186), .d(new_n230), .o1(new_n231));
  aoi012aa1n03x5               g136(.a(new_n226), .b(new_n231), .c(new_n229), .o1(new_n232));
  norp02aa1n03x5               g137(.a(new_n232), .b(new_n228), .o1(\s[22] ));
  nanb02aa1n12x5               g138(.a(new_n226), .b(new_n225), .out0(new_n234));
  nano22aa1n12x5               g139(.a(new_n234), .b(new_n196), .c(new_n215), .out0(new_n235));
  oaoi03aa1n12x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n229), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n218), .d(new_n219), .o1(new_n238));
  xorc02aa1n12x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n238), .c(new_n186), .d(new_n235), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n132), .o1(new_n242));
  aoai13aa1n02x5               g147(.a(new_n159), .b(new_n145), .c(new_n178), .d(new_n242), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n179), .o1(new_n244));
  aoai13aa1n02x5               g149(.a(new_n185), .b(new_n244), .c(new_n243), .d(new_n161), .o1(new_n245));
  aoai13aa1n02x5               g150(.a(new_n235), .b(new_n245), .c(new_n164), .d(new_n181), .o1(new_n246));
  nona22aa1n02x4               g151(.a(new_n246), .b(new_n238), .c(new_n240), .out0(new_n247));
  nanp02aa1n02x5               g152(.a(new_n241), .b(new_n247), .o1(\s[23] ));
  nanp02aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  aoi112aa1n03x5               g154(.a(new_n240), .b(new_n238), .c(new_n186), .d(new_n235), .o1(new_n250));
  tech160nm_fixorc02aa1n05x5   g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  nano22aa1n03x5               g156(.a(new_n250), .b(new_n249), .c(new_n251), .out0(new_n252));
  aoi012aa1n02x5               g157(.a(new_n251), .b(new_n247), .c(new_n249), .o1(new_n253));
  norp02aa1n02x5               g158(.a(new_n253), .b(new_n252), .o1(\s[24] ));
  nand02aa1n04x5               g159(.a(new_n251), .b(new_n239), .o1(new_n255));
  nor043aa1n02x5               g160(.a(new_n216), .b(new_n234), .c(new_n255), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  norb02aa1d21x5               g162(.a(new_n225), .b(new_n226), .out0(new_n258));
  inv030aa1n06x5               g163(.a(new_n255), .o1(new_n259));
  norp02aa1n02x5               g164(.a(\b[23] ), .b(\a[24] ), .o1(new_n260));
  aoi112aa1n02x5               g165(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n261));
  nanp03aa1d12x5               g166(.a(new_n236), .b(new_n239), .c(new_n251), .o1(new_n262));
  nona22aa1d18x5               g167(.a(new_n262), .b(new_n261), .c(new_n260), .out0(new_n263));
  aoi013aa1n09x5               g168(.a(new_n263), .b(new_n220), .c(new_n259), .d(new_n258), .o1(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n257), .c(new_n192), .d(new_n182), .o1(new_n265));
  xorb03aa1n02x5               g170(.a(new_n265), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1d18x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  tech160nm_fixorc02aa1n04x5   g172(.a(\a[25] ), .b(\b[24] ), .out0(new_n268));
  xorc02aa1n12x5               g173(.a(\a[26] ), .b(\b[25] ), .out0(new_n269));
  aoi112aa1n03x5               g174(.a(new_n267), .b(new_n269), .c(new_n265), .d(new_n268), .o1(new_n270));
  inv020aa1n03x5               g175(.a(new_n267), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n264), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n268), .b(new_n272), .c(new_n186), .d(new_n256), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n269), .o1(new_n274));
  aoi012aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n271), .o1(new_n275));
  nor002aa1n02x5               g180(.a(new_n275), .b(new_n270), .o1(\s[26] ));
  and002aa1n12x5               g181(.a(new_n269), .b(new_n268), .o(new_n277));
  nano23aa1n06x5               g182(.a(new_n216), .b(new_n255), .c(new_n277), .d(new_n258), .out0(new_n278));
  inv020aa1n03x5               g183(.a(new_n278), .o1(new_n279));
  aoi112aa1n06x5               g184(.a(new_n234), .b(new_n255), .c(new_n218), .d(new_n219), .o1(new_n280));
  tech160nm_fioaoi03aa1n02p5x5 g185(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .o1(new_n281));
  oaoi13aa1n09x5               g186(.a(new_n281), .b(new_n277), .c(new_n280), .d(new_n263), .o1(new_n282));
  aoai13aa1n04x5               g187(.a(new_n282), .b(new_n279), .c(new_n192), .d(new_n182), .o1(new_n283));
  xorb03aa1n03x5               g188(.a(new_n283), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nanp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .out0(new_n286));
  inv000aa1d42x5               g191(.a(new_n263), .o1(new_n287));
  nanp03aa1n03x5               g192(.a(new_n220), .b(new_n258), .c(new_n259), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n277), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n281), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n289), .c(new_n287), .d(new_n288), .o1(new_n291));
  nor042aa1d18x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  aoi112aa1n03x4               g197(.a(new_n292), .b(new_n291), .c(new_n186), .d(new_n278), .o1(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n285), .c(new_n286), .out0(new_n294));
  aoai13aa1n02x5               g199(.a(new_n278), .b(new_n245), .c(new_n164), .d(new_n181), .o1(new_n295));
  nona22aa1n03x5               g200(.a(new_n295), .b(new_n291), .c(new_n292), .out0(new_n296));
  aoi012aa1n03x5               g201(.a(new_n286), .b(new_n296), .c(new_n285), .o1(new_n297));
  norp02aa1n03x5               g202(.a(new_n297), .b(new_n294), .o1(\s[28] ));
  nano22aa1n02x4               g203(.a(new_n292), .b(new_n286), .c(new_n285), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n291), .c(new_n186), .d(new_n278), .o1(new_n300));
  inv000aa1d42x5               g205(.a(\a[28] ), .o1(new_n301));
  inv000aa1d42x5               g206(.a(\b[27] ), .o1(new_n302));
  oaoi03aa1n12x5               g207(.a(new_n301), .b(new_n302), .c(new_n292), .o1(new_n303));
  tech160nm_fixorc02aa1n02p5x5 g208(.a(\a[29] ), .b(\b[28] ), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  tech160nm_fiaoi012aa1n02p5x5 g210(.a(new_n305), .b(new_n300), .c(new_n303), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n303), .o1(new_n307));
  aoi112aa1n02x7               g212(.a(new_n304), .b(new_n307), .c(new_n283), .d(new_n299), .o1(new_n308));
  nor002aa1n02x5               g213(.a(new_n306), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g215(.a(new_n305), .b(new_n292), .c(new_n286), .d(new_n285), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n291), .c(new_n186), .d(new_n278), .o1(new_n312));
  tech160nm_fioaoi03aa1n03p5x5 g217(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .o1(new_n313));
  inv030aa1n02x5               g218(.a(new_n313), .o1(new_n314));
  tech160nm_fixorc02aa1n02p5x5 g219(.a(\a[30] ), .b(\b[29] ), .out0(new_n315));
  inv000aa1d42x5               g220(.a(new_n315), .o1(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n312), .c(new_n314), .o1(new_n317));
  aoi112aa1n03x4               g222(.a(new_n315), .b(new_n313), .c(new_n283), .d(new_n311), .o1(new_n318));
  norp02aa1n03x5               g223(.a(new_n317), .b(new_n318), .o1(\s[30] ));
  and003aa1n03x7               g224(.a(new_n299), .b(new_n315), .c(new_n304), .o(new_n320));
  oaoi03aa1n03x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n314), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  aoi112aa1n03x4               g227(.a(new_n322), .b(new_n321), .c(new_n283), .d(new_n320), .o1(new_n323));
  aoai13aa1n03x5               g228(.a(new_n320), .b(new_n291), .c(new_n186), .d(new_n278), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n321), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n322), .o1(new_n326));
  tech160nm_fiaoi012aa1n02p5x5 g231(.a(new_n326), .b(new_n324), .c(new_n325), .o1(new_n327));
  norp02aa1n03x5               g232(.a(new_n327), .b(new_n323), .o1(\s[31] ));
  xnrb03aa1n02x5               g233(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g234(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g236(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g237(.a(new_n119), .b(new_n120), .c(new_n107), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(new_n116), .out0(\s[6] ));
  nanb02aa1n02x5               g239(.a(new_n110), .b(new_n111), .out0(new_n335));
  oaoi13aa1n02x5               g240(.a(new_n335), .b(new_n118), .c(new_n333), .d(new_n113), .o1(new_n336));
  oai112aa1n02x5               g241(.a(new_n118), .b(new_n335), .c(new_n333), .d(new_n113), .o1(new_n337));
  norb02aa1n02x5               g242(.a(new_n337), .b(new_n336), .out0(\s[7] ));
  norp02aa1n02x5               g243(.a(new_n336), .b(new_n110), .o1(new_n339));
  xnrb03aa1n02x5               g244(.a(new_n339), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrc02aa1n02x5               g245(.a(new_n124), .b(new_n177), .out0(\s[9] ));
endmodule


