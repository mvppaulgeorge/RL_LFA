// Benchmark "adder" written by ABC on Wed Jul 17 20:14:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n338,
    new_n341, new_n343, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d30x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nand02aa1d04x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nona23aa1n09x5               g008(.a(new_n102), .b(new_n101), .c(new_n103), .d(new_n100), .out0(new_n104));
  norp02aa1n03x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nand22aa1n03x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nor022aa1n03x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nona23aa1n03x5               g013(.a(new_n107), .b(new_n106), .c(new_n108), .d(new_n105), .out0(new_n109));
  nor042aa1n02x5               g014(.a(new_n109), .b(new_n104), .o1(new_n110));
  and002aa1n06x5               g015(.a(\b[3] ), .b(\a[4] ), .o(new_n111));
  inv000aa1d42x5               g016(.a(\a[3] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[2] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(new_n113), .b(new_n112), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(new_n114), .b(new_n115), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  nor042aa1n02x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  nand22aa1n03x5               g023(.a(\b[0] ), .b(\a[1] ), .o1(new_n119));
  tech160nm_fioai012aa1n05x5   g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  oa0022aa1n02x5               g025(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n121));
  oaoi13aa1n12x5               g026(.a(new_n111), .b(new_n121), .c(new_n120), .d(new_n116), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n100), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n103), .b(new_n101), .o1(new_n124));
  oai012aa1n02x5               g029(.a(new_n106), .b(new_n108), .c(new_n105), .o1(new_n125));
  oai112aa1n03x5               g030(.a(new_n123), .b(new_n124), .c(new_n104), .d(new_n125), .o1(new_n126));
  xorc02aa1n02x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n128));
  nor002aa1d32x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n128), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g037(.a(new_n129), .o1(new_n133));
  inv000aa1n04x5               g038(.a(new_n130), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand22aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  aoi113aa1n02x5               g043(.a(new_n138), .b(new_n134), .c(new_n128), .d(new_n133), .e(new_n99), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n111), .o1(new_n140));
  oai012aa1n04x7               g045(.a(new_n121), .b(new_n120), .c(new_n116), .o1(new_n141));
  nona23aa1n09x5               g046(.a(new_n141), .b(new_n140), .c(new_n104), .d(new_n109), .out0(new_n142));
  norp02aa1n02x5               g047(.a(new_n104), .b(new_n125), .o1(new_n143));
  nano22aa1n03x7               g048(.a(new_n143), .b(new_n123), .c(new_n124), .out0(new_n144));
  and002aa1n02x5               g049(.a(\b[8] ), .b(\a[9] ), .o(new_n145));
  aoai13aa1n02x5               g050(.a(new_n99), .b(new_n145), .c(new_n142), .d(new_n144), .o1(new_n146));
  aoai13aa1n12x5               g051(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  aoi112aa1n02x5               g053(.a(new_n148), .b(new_n137), .c(new_n146), .d(new_n131), .o1(new_n149));
  norp02aa1n02x5               g054(.a(new_n149), .b(new_n139), .o1(\s[11] ));
  nor022aa1n12x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nanp02aa1n12x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  norp03aa1n02x5               g058(.a(new_n139), .b(new_n153), .c(new_n135), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n135), .o1(new_n155));
  aoai13aa1n03x5               g060(.a(new_n137), .b(new_n148), .c(new_n146), .d(new_n131), .o1(new_n156));
  aobi12aa1n02x5               g061(.a(new_n153), .b(new_n156), .c(new_n155), .out0(new_n157));
  norp02aa1n03x5               g062(.a(new_n157), .b(new_n154), .o1(\s[12] ));
  inv000aa1n02x5               g063(.a(new_n136), .o1(new_n159));
  aoi112aa1n06x5               g064(.a(new_n134), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n160));
  norb03aa1n12x5               g065(.a(new_n152), .b(new_n135), .c(new_n151), .out0(new_n161));
  nona23aa1d18x5               g066(.a(new_n160), .b(new_n161), .c(new_n159), .d(new_n145), .out0(new_n162));
  nona23aa1n09x5               g067(.a(new_n152), .b(new_n136), .c(new_n135), .d(new_n151), .out0(new_n163));
  tech160nm_fioai012aa1n03p5x5 g068(.a(new_n152), .b(new_n151), .c(new_n135), .o1(new_n164));
  oai012aa1d24x5               g069(.a(new_n164), .b(new_n163), .c(new_n147), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n162), .c(new_n142), .d(new_n144), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n12x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nand42aa1n02x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n169), .b(new_n167), .c(new_n170), .o1(new_n171));
  xnrb03aa1n02x5               g076(.a(new_n171), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g077(.a(new_n162), .o1(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n174));
  nor022aa1n06x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nand42aa1n03x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  oai012aa1n12x5               g081(.a(new_n176), .b(new_n175), .c(new_n169), .o1(new_n177));
  nona23aa1n03x5               g082(.a(new_n176), .b(new_n170), .c(new_n169), .d(new_n175), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n177), .b(new_n178), .c(new_n174), .d(new_n166), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n02x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  nand02aa1n02x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nanb02aa1n02x5               g087(.a(new_n181), .b(new_n182), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  norp02aa1n02x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nanp02aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nanb02aa1n02x5               g091(.a(new_n185), .b(new_n186), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(new_n188), .b(new_n181), .c(new_n179), .d(new_n184), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n177), .o1(new_n190));
  nano23aa1n02x4               g095(.a(new_n169), .b(new_n175), .c(new_n176), .d(new_n170), .out0(new_n191));
  aoai13aa1n02x7               g096(.a(new_n184), .b(new_n190), .c(new_n167), .d(new_n191), .o1(new_n192));
  oaoi13aa1n03x5               g097(.a(new_n187), .b(new_n192), .c(\a[15] ), .d(\b[14] ), .o1(new_n193));
  nor002aa1n02x5               g098(.a(new_n193), .b(new_n189), .o1(\s[16] ));
  nano23aa1n02x4               g099(.a(new_n181), .b(new_n185), .c(new_n186), .d(new_n182), .out0(new_n195));
  nano22aa1n03x7               g100(.a(new_n162), .b(new_n191), .c(new_n195), .out0(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n126), .c(new_n122), .d(new_n110), .o1(new_n197));
  nona23aa1n03x5               g102(.a(new_n186), .b(new_n182), .c(new_n181), .d(new_n185), .out0(new_n198));
  nor002aa1n02x5               g103(.a(new_n198), .b(new_n178), .o1(new_n199));
  aoi112aa1n02x5               g104(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n200));
  oai022aa1n03x5               g105(.a(new_n198), .b(new_n177), .c(\b[15] ), .d(\a[16] ), .o1(new_n201));
  aoi112aa1n09x5               g106(.a(new_n201), .b(new_n200), .c(new_n165), .d(new_n199), .o1(new_n202));
  nanp02aa1n06x5               g107(.a(new_n197), .b(new_n202), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g109(.a(\a[17] ), .o1(new_n205));
  inv000aa1d42x5               g110(.a(\b[16] ), .o1(new_n206));
  oaoi03aa1n03x5               g111(.a(new_n205), .b(new_n206), .c(new_n203), .o1(new_n207));
  xnrb03aa1n03x5               g112(.a(new_n207), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n02x5               g113(.a(new_n206), .b(new_n205), .o1(new_n209));
  nanp02aa1n02x5               g114(.a(\b[16] ), .b(\a[17] ), .o1(new_n210));
  nor022aa1n06x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nand42aa1n03x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nanb02aa1n02x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  nano22aa1n03x7               g118(.a(new_n213), .b(new_n209), .c(new_n210), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n09x5               g120(.a(new_n212), .b(new_n211), .c(new_n205), .d(new_n206), .o1(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n215), .c(new_n197), .d(new_n202), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  nor042aa1n02x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nanb02aa1n02x5               g128(.a(new_n222), .b(new_n223), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  aoi112aa1n02x7               g130(.a(new_n225), .b(new_n220), .c(new_n217), .d(new_n221), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n220), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n221), .b(new_n220), .out0(new_n228));
  nanp02aa1n03x5               g133(.a(new_n217), .b(new_n228), .o1(new_n229));
  aoi012aa1n03x5               g134(.a(new_n224), .b(new_n229), .c(new_n227), .o1(new_n230));
  norp02aa1n03x5               g135(.a(new_n230), .b(new_n226), .o1(\s[20] ));
  nano23aa1n06x5               g136(.a(new_n220), .b(new_n222), .c(new_n223), .d(new_n221), .out0(new_n232));
  nanp02aa1n02x5               g137(.a(new_n214), .b(new_n232), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n216), .o1(new_n234));
  oaih12aa1n02x5               g139(.a(new_n223), .b(new_n222), .c(new_n220), .o1(new_n235));
  aobi12aa1n06x5               g140(.a(new_n235), .b(new_n232), .c(new_n234), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n233), .c(new_n197), .d(new_n202), .o1(new_n237));
  xorb03aa1n02x5               g142(.a(new_n237), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  xorc02aa1n02x5               g144(.a(\a[21] ), .b(\b[20] ), .out0(new_n240));
  xorc02aa1n02x5               g145(.a(\a[22] ), .b(\b[21] ), .out0(new_n241));
  aoi112aa1n03x5               g146(.a(new_n239), .b(new_n241), .c(new_n237), .d(new_n240), .o1(new_n242));
  inv000aa1n02x5               g147(.a(new_n239), .o1(new_n243));
  nanp02aa1n03x5               g148(.a(new_n237), .b(new_n240), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n241), .o1(new_n245));
  tech160nm_fiaoi012aa1n05x5   g150(.a(new_n245), .b(new_n244), .c(new_n243), .o1(new_n246));
  nor042aa1n03x5               g151(.a(new_n246), .b(new_n242), .o1(\s[22] ));
  inv000aa1d42x5               g152(.a(\a[21] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(\a[22] ), .o1(new_n249));
  xroi22aa1d04x5               g154(.a(new_n248), .b(\b[20] ), .c(new_n249), .d(\b[21] ), .out0(new_n250));
  nand23aa1n03x5               g155(.a(new_n250), .b(new_n214), .c(new_n232), .o1(new_n251));
  nona23aa1n09x5               g156(.a(new_n223), .b(new_n221), .c(new_n220), .d(new_n222), .out0(new_n252));
  tech160nm_fioai012aa1n03p5x5 g157(.a(new_n235), .b(new_n252), .c(new_n216), .o1(new_n253));
  oao003aa1n02x5               g158(.a(\a[22] ), .b(\b[21] ), .c(new_n243), .carry(new_n254));
  aobi12aa1n02x5               g159(.a(new_n254), .b(new_n253), .c(new_n250), .out0(new_n255));
  aoai13aa1n04x5               g160(.a(new_n255), .b(new_n251), .c(new_n197), .d(new_n202), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n04x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  nor002aa1n02x5               g164(.a(\b[23] ), .b(\a[24] ), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(\b[23] ), .b(\a[24] ), .o1(new_n261));
  norb02aa1n02x5               g166(.a(new_n261), .b(new_n260), .out0(new_n262));
  aoi112aa1n02x7               g167(.a(new_n258), .b(new_n262), .c(new_n256), .d(new_n259), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n258), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n259), .b(new_n258), .out0(new_n265));
  nand42aa1n02x5               g170(.a(new_n256), .b(new_n265), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n262), .o1(new_n267));
  aoi012aa1n03x5               g172(.a(new_n267), .b(new_n266), .c(new_n264), .o1(new_n268));
  nor042aa1n03x5               g173(.a(new_n268), .b(new_n263), .o1(\s[24] ));
  nona23aa1d18x5               g174(.a(new_n261), .b(new_n259), .c(new_n258), .d(new_n260), .out0(new_n270));
  nona23aa1n02x4               g175(.a(new_n250), .b(new_n214), .c(new_n270), .d(new_n252), .out0(new_n271));
  inv000aa1d42x5               g176(.a(new_n270), .o1(new_n272));
  oai012aa1n02x5               g177(.a(new_n261), .b(new_n260), .c(new_n258), .o1(new_n273));
  oai012aa1n12x5               g178(.a(new_n273), .b(new_n254), .c(new_n270), .o1(new_n274));
  aoi013aa1n02x4               g179(.a(new_n274), .b(new_n253), .c(new_n250), .d(new_n272), .o1(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n271), .c(new_n197), .d(new_n202), .o1(new_n276));
  xorb03aa1n02x5               g181(.a(new_n276), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g182(.a(\b[24] ), .b(\a[25] ), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[25] ), .b(\b[24] ), .out0(new_n279));
  xorc02aa1n12x5               g184(.a(\a[26] ), .b(\b[25] ), .out0(new_n280));
  aoi112aa1n02x5               g185(.a(new_n278), .b(new_n280), .c(new_n276), .d(new_n279), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n278), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(new_n276), .b(new_n279), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n280), .o1(new_n284));
  aoi012aa1n03x5               g189(.a(new_n284), .b(new_n283), .c(new_n282), .o1(new_n285));
  norp02aa1n02x5               g190(.a(new_n285), .b(new_n281), .o1(\s[26] ));
  nand42aa1n02x5               g191(.a(new_n142), .b(new_n144), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(new_n165), .b(new_n199), .o1(new_n288));
  nona22aa1n03x5               g193(.a(new_n288), .b(new_n201), .c(new_n200), .out0(new_n289));
  and002aa1n06x5               g194(.a(new_n280), .b(new_n279), .o(new_n290));
  nano22aa1n03x7               g195(.a(new_n251), .b(new_n290), .c(new_n272), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n289), .c(new_n287), .d(new_n196), .o1(new_n292));
  nano22aa1n03x7               g197(.a(new_n236), .b(new_n250), .c(new_n272), .out0(new_n293));
  oao003aa1n02x5               g198(.a(\a[26] ), .b(\b[25] ), .c(new_n282), .carry(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  oaoi13aa1n09x5               g200(.a(new_n295), .b(new_n290), .c(new_n293), .d(new_n274), .o1(new_n296));
  nor042aa1n03x5               g201(.a(\b[26] ), .b(\a[27] ), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  norb02aa1n02x5               g203(.a(new_n298), .b(new_n297), .out0(new_n299));
  xnbna2aa1n03x5               g204(.a(new_n299), .b(new_n292), .c(new_n296), .out0(\s[27] ));
  inv000aa1d42x5               g205(.a(new_n297), .o1(new_n301));
  aobi12aa1n02x5               g206(.a(new_n299), .b(new_n292), .c(new_n296), .out0(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .out0(new_n303));
  nano22aa1n02x4               g208(.a(new_n302), .b(new_n301), .c(new_n303), .out0(new_n304));
  inv000aa1n02x5               g209(.a(new_n274), .o1(new_n305));
  nanp03aa1n02x5               g210(.a(new_n253), .b(new_n250), .c(new_n272), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n290), .o1(new_n307));
  aoai13aa1n06x5               g212(.a(new_n294), .b(new_n307), .c(new_n306), .d(new_n305), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n299), .b(new_n308), .c(new_n203), .d(new_n291), .o1(new_n309));
  aoi012aa1n03x5               g214(.a(new_n303), .b(new_n309), .c(new_n301), .o1(new_n310));
  nor002aa1n02x5               g215(.a(new_n310), .b(new_n304), .o1(\s[28] ));
  xnrc02aa1n02x5               g216(.a(\b[28] ), .b(\a[29] ), .out0(new_n312));
  nano22aa1n02x4               g217(.a(new_n303), .b(new_n301), .c(new_n298), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n308), .c(new_n203), .d(new_n291), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[28] ), .b(\b[27] ), .c(new_n301), .carry(new_n315));
  aoi012aa1n03x5               g220(.a(new_n312), .b(new_n314), .c(new_n315), .o1(new_n316));
  aobi12aa1n02x5               g221(.a(new_n313), .b(new_n292), .c(new_n296), .out0(new_n317));
  nano22aa1n02x4               g222(.a(new_n317), .b(new_n312), .c(new_n315), .out0(new_n318));
  nor002aa1n02x5               g223(.a(new_n316), .b(new_n318), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n119), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g225(.a(new_n312), .b(new_n303), .c(new_n298), .d(new_n301), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n308), .c(new_n203), .d(new_n291), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(new_n315), .carry(new_n323));
  xnrc02aa1n02x5               g228(.a(\b[29] ), .b(\a[30] ), .out0(new_n324));
  aoi012aa1n03x5               g229(.a(new_n324), .b(new_n322), .c(new_n323), .o1(new_n325));
  aobi12aa1n02x5               g230(.a(new_n321), .b(new_n292), .c(new_n296), .out0(new_n326));
  nano22aa1n02x4               g231(.a(new_n326), .b(new_n323), .c(new_n324), .out0(new_n327));
  nor002aa1n02x5               g232(.a(new_n325), .b(new_n327), .o1(\s[30] ));
  norb03aa1n02x5               g233(.a(new_n313), .b(new_n312), .c(new_n324), .out0(new_n329));
  aobi12aa1n02x5               g234(.a(new_n329), .b(new_n292), .c(new_n296), .out0(new_n330));
  oao003aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .c(new_n323), .carry(new_n331));
  xnrc02aa1n02x5               g236(.a(\b[30] ), .b(\a[31] ), .out0(new_n332));
  nano22aa1n02x4               g237(.a(new_n330), .b(new_n331), .c(new_n332), .out0(new_n333));
  aoai13aa1n03x5               g238(.a(new_n329), .b(new_n308), .c(new_n203), .d(new_n291), .o1(new_n334));
  aoi012aa1n03x5               g239(.a(new_n332), .b(new_n334), .c(new_n331), .o1(new_n335));
  nor002aa1n02x5               g240(.a(new_n335), .b(new_n333), .o1(\s[31] ));
  xnbna2aa1n03x5               g241(.a(new_n120), .b(new_n114), .c(new_n115), .out0(\s[3] ));
  oaoi03aa1n02x5               g242(.a(\a[3] ), .b(\b[2] ), .c(new_n120), .o1(new_n338));
  xorb03aa1n02x5               g243(.a(new_n338), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g244(.a(new_n122), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi013aa1n02x4               g245(.a(new_n108), .b(new_n141), .c(new_n140), .d(new_n107), .o1(new_n341));
  xnrb03aa1n02x5               g246(.a(new_n341), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi113aa1n02x5               g247(.a(new_n108), .b(new_n105), .c(new_n141), .d(new_n140), .e(new_n107), .o1(new_n343));
  norb02aa1n02x5               g248(.a(new_n106), .b(new_n343), .out0(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g250(.a(new_n103), .b(new_n344), .c(new_n102), .o1(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n123), .c(new_n101), .out0(\s[8] ));
  xnbna2aa1n03x5               g252(.a(new_n127), .b(new_n142), .c(new_n144), .out0(\s[9] ));
endmodule


