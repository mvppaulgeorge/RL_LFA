// Benchmark "adder" written by ABC on Thu Jul 18 02:23:27 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n331,
    new_n334, new_n335, new_n336, new_n338, new_n339, new_n341, new_n342,
    new_n343;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv030aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[4] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[3] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand02aa1d10x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nor042aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n03x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb02aa1n02x5               g010(.a(new_n104), .b(new_n105), .out0(new_n106));
  nano32aa1n03x7               g011(.a(new_n106), .b(new_n101), .c(new_n102), .d(new_n103), .out0(new_n107));
  nand02aa1n04x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  norb03aa1n03x5               g014(.a(new_n103), .b(new_n109), .c(new_n108), .out0(new_n110));
  inv000aa1n06x5               g015(.a(new_n110), .o1(new_n111));
  oaoi03aa1n09x5               g016(.a(new_n99), .b(new_n100), .c(new_n104), .o1(new_n112));
  inv000aa1d42x5               g017(.a(new_n112), .o1(new_n113));
  nor002aa1d24x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor022aa1n06x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nand42aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nona23aa1n03x5               g022(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n118));
  nor022aa1n04x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nand22aa1n09x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nor002aa1d32x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nand02aa1n03x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  nona23aa1n09x5               g027(.a(new_n122), .b(new_n120), .c(new_n119), .d(new_n121), .out0(new_n123));
  nor042aa1n03x5               g028(.a(new_n123), .b(new_n118), .o1(new_n124));
  aoai13aa1n12x5               g029(.a(new_n124), .b(new_n113), .c(new_n107), .d(new_n111), .o1(new_n125));
  inv000aa1d42x5               g030(.a(new_n114), .o1(new_n126));
  aob012aa1n02x5               g031(.a(new_n126), .b(new_n116), .c(new_n115), .out0(new_n127));
  oai022aa1n02x5               g032(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n128));
  aboi22aa1n09x5               g033(.a(new_n123), .b(new_n127), .c(new_n128), .d(new_n120), .out0(new_n129));
  nand02aa1d08x5               g034(.a(new_n125), .b(new_n129), .o1(new_n130));
  nand02aa1n04x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n97), .b(new_n131), .out0(new_n132));
  nanb02aa1n02x5               g037(.a(new_n132), .b(new_n130), .out0(new_n133));
  nor002aa1n04x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nanp02aa1n04x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n136), .b(new_n133), .c(new_n98), .out0(\s[10] ));
  nona23aa1d18x5               g042(.a(new_n135), .b(new_n131), .c(new_n97), .d(new_n134), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  oaoi03aa1n09x5               g044(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n140));
  nor002aa1n10x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nand42aa1n06x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  norb02aa1n02x7               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  aoai13aa1n06x5               g048(.a(new_n143), .b(new_n140), .c(new_n130), .d(new_n139), .o1(new_n144));
  aoi112aa1n02x5               g049(.a(new_n143), .b(new_n140), .c(new_n130), .d(new_n139), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n144), .b(new_n145), .out0(\s[11] ));
  inv000aa1n02x5               g051(.a(new_n141), .o1(new_n147));
  nor042aa1n02x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nanp02aa1n03x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  norb02aa1n06x4               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n144), .c(new_n147), .out0(\s[12] ));
  nano22aa1n12x5               g056(.a(new_n138), .b(new_n143), .c(new_n150), .out0(new_n152));
  nano23aa1n09x5               g057(.a(new_n141), .b(new_n148), .c(new_n149), .d(new_n142), .out0(new_n153));
  oaoi03aa1n02x5               g058(.a(\a[12] ), .b(\b[11] ), .c(new_n147), .o1(new_n154));
  tech160nm_fiao0012aa1n02p5x5 g059(.a(new_n154), .b(new_n153), .c(new_n140), .o(new_n155));
  xnrc02aa1n12x5               g060(.a(\b[12] ), .b(\a[13] ), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n155), .c(new_n130), .d(new_n152), .o1(new_n158));
  aoi112aa1n02x5               g063(.a(new_n157), .b(new_n155), .c(new_n130), .d(new_n152), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(\s[13] ));
  orn002aa1n02x5               g065(.a(\a[13] ), .b(\b[12] ), .o(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[13] ), .b(\a[14] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n158), .c(new_n161), .out0(\s[14] ));
  nor042aa1n06x5               g069(.a(new_n162), .b(new_n156), .o1(new_n165));
  nano22aa1n02x4               g070(.a(new_n138), .b(new_n165), .c(new_n153), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n165), .b(new_n154), .c(new_n153), .d(new_n140), .o1(new_n167));
  oao003aa1n02x5               g072(.a(\a[14] ), .b(\b[13] ), .c(new_n161), .carry(new_n168));
  nand22aa1n03x5               g073(.a(new_n167), .b(new_n168), .o1(new_n169));
  xorc02aa1n02x5               g074(.a(\a[15] ), .b(\b[14] ), .out0(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n169), .c(new_n130), .d(new_n166), .o1(new_n171));
  nanb03aa1n02x5               g076(.a(new_n170), .b(new_n167), .c(new_n168), .out0(new_n172));
  aoi012aa1n02x5               g077(.a(new_n172), .b(new_n130), .c(new_n166), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n171), .b(new_n173), .out0(\s[15] ));
  inv000aa1d42x5               g079(.a(\a[15] ), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(\b[14] ), .b(new_n175), .out0(new_n176));
  xorc02aa1n02x5               g081(.a(\a[16] ), .b(\b[15] ), .out0(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n171), .c(new_n176), .out0(\s[16] ));
  inv000aa1d42x5               g083(.a(\a[17] ), .o1(new_n179));
  inv020aa1n04x5               g084(.a(\a[16] ), .o1(new_n180));
  xroi22aa1d06x4               g085(.a(new_n175), .b(\b[14] ), .c(new_n180), .d(\b[15] ), .out0(new_n181));
  nand23aa1n06x5               g086(.a(new_n152), .b(new_n165), .c(new_n181), .o1(new_n182));
  aoi012aa1d18x5               g087(.a(new_n182), .b(new_n125), .c(new_n129), .o1(new_n183));
  inv000aa1n02x5               g088(.a(new_n181), .o1(new_n184));
  oao003aa1n02x5               g089(.a(\a[16] ), .b(\b[15] ), .c(new_n176), .carry(new_n185));
  aoai13aa1n12x5               g090(.a(new_n185), .b(new_n184), .c(new_n167), .d(new_n168), .o1(new_n186));
  nor042aa1n03x5               g091(.a(new_n186), .b(new_n183), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(new_n179), .out0(\s[17] ));
  obai22aa1n02x7               g093(.a(\b[16] ), .b(new_n179), .c(\b[17] ), .d(\a[18] ), .out0(new_n189));
  aoi012aa1n02x5               g094(.a(new_n189), .b(\a[18] ), .c(\b[17] ), .o1(new_n190));
  oaib12aa1n06x5               g095(.a(new_n187), .b(\b[16] ), .c(new_n179), .out0(new_n191));
  xnrc02aa1n02x5               g096(.a(\b[17] ), .b(\a[18] ), .out0(new_n192));
  oaib12aa1n02x5               g097(.a(new_n191), .b(new_n179), .c(\b[16] ), .out0(new_n193));
  aoi022aa1n02x5               g098(.a(new_n193), .b(new_n192), .c(new_n190), .d(new_n191), .o1(\s[18] ));
  inv040aa1n16x5               g099(.a(\a[18] ), .o1(new_n195));
  xroi22aa1d06x4               g100(.a(new_n179), .b(\b[16] ), .c(new_n195), .d(\b[17] ), .out0(new_n196));
  oai012aa1n06x5               g101(.a(new_n196), .b(new_n186), .c(new_n183), .o1(new_n197));
  inv040aa1d32x5               g102(.a(\b[17] ), .o1(new_n198));
  nor042aa1n06x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  oao003aa1n12x5               g104(.a(new_n195), .b(new_n198), .c(new_n199), .carry(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  nor042aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand42aa1n04x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n197), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g111(.a(new_n101), .b(new_n102), .o1(new_n207));
  nanb03aa1n06x5               g112(.a(new_n104), .b(new_n105), .c(new_n103), .out0(new_n208));
  oai013aa1n06x5               g113(.a(new_n112), .b(new_n110), .c(new_n208), .d(new_n207), .o1(new_n209));
  oai012aa1n02x5               g114(.a(new_n120), .b(new_n121), .c(new_n119), .o1(new_n210));
  oaib12aa1n02x5               g115(.a(new_n210), .b(new_n123), .c(new_n127), .out0(new_n211));
  tech160nm_fiaoi012aa1n05x5   g116(.a(new_n211), .b(new_n209), .c(new_n124), .o1(new_n212));
  nanp02aa1n03x5               g117(.a(new_n169), .b(new_n181), .o1(new_n213));
  oai112aa1n06x5               g118(.a(new_n213), .b(new_n185), .c(new_n212), .d(new_n182), .o1(new_n214));
  aoai13aa1n02x5               g119(.a(new_n204), .b(new_n200), .c(new_n214), .d(new_n196), .o1(new_n215));
  nor002aa1n03x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand02aa1n06x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  aoib12aa1n02x5               g123(.a(new_n202), .b(new_n217), .c(new_n216), .out0(new_n219));
  inv000aa1n02x5               g124(.a(new_n202), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n204), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n220), .b(new_n221), .c(new_n197), .d(new_n201), .o1(new_n222));
  aoi022aa1n02x7               g127(.a(new_n222), .b(new_n218), .c(new_n215), .d(new_n219), .o1(\s[20] ));
  nano23aa1d15x5               g128(.a(new_n202), .b(new_n216), .c(new_n217), .d(new_n203), .out0(new_n224));
  nand02aa1n04x5               g129(.a(new_n196), .b(new_n224), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  oai012aa1n06x5               g131(.a(new_n226), .b(new_n186), .c(new_n183), .o1(new_n227));
  oaoi03aa1n12x5               g132(.a(\a[20] ), .b(\b[19] ), .c(new_n220), .o1(new_n228));
  aoi012aa1d24x5               g133(.a(new_n228), .b(new_n224), .c(new_n200), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  xnbna2aa1n03x5               g136(.a(new_n231), .b(new_n227), .c(new_n229), .out0(\s[21] ));
  inv000aa1d42x5               g137(.a(new_n229), .o1(new_n233));
  aoai13aa1n03x5               g138(.a(new_n231), .b(new_n233), .c(new_n214), .d(new_n226), .o1(new_n234));
  nor002aa1n06x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  nand02aa1d06x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  nanb02aa1d24x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  nor042aa1n09x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  aoib12aa1n02x5               g144(.a(new_n239), .b(new_n236), .c(new_n235), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n239), .o1(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n230), .c(new_n227), .d(new_n229), .o1(new_n242));
  aoi022aa1n02x5               g147(.a(new_n242), .b(new_n238), .c(new_n234), .d(new_n240), .o1(\s[22] ));
  nor042aa1n06x5               g148(.a(new_n230), .b(new_n237), .o1(new_n244));
  and003aa1n02x5               g149(.a(new_n196), .b(new_n244), .c(new_n224), .o(new_n245));
  aoi012aa1n02x5               g150(.a(new_n235), .b(new_n239), .c(new_n236), .o1(new_n246));
  oaib12aa1n03x5               g151(.a(new_n246), .b(new_n229), .c(new_n244), .out0(new_n247));
  xnrc02aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .out0(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n247), .c(new_n214), .d(new_n245), .o1(new_n249));
  oaih12aa1n02x5               g154(.a(new_n245), .b(new_n186), .c(new_n183), .o1(new_n250));
  norp02aa1n02x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  and002aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o(new_n252));
  nona32aa1n03x5               g157(.a(new_n250), .b(new_n252), .c(new_n251), .d(new_n247), .out0(new_n253));
  nanp02aa1n02x5               g158(.a(new_n249), .b(new_n253), .o1(\s[23] ));
  and002aa1n02x5               g159(.a(\b[23] ), .b(\a[24] ), .o(new_n255));
  norp02aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n255), .b(new_n256), .c(\a[23] ), .d(\b[22] ), .o1(new_n257));
  xnrc02aa1n02x5               g162(.a(\b[23] ), .b(\a[24] ), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n252), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(new_n253), .b(new_n259), .o1(new_n260));
  aoi022aa1n02x7               g165(.a(new_n260), .b(new_n258), .c(new_n253), .d(new_n257), .o1(\s[24] ));
  norp02aa1n04x5               g166(.a(new_n258), .b(new_n248), .o1(new_n262));
  nand02aa1d04x5               g167(.a(new_n262), .b(new_n244), .o1(new_n263));
  nano22aa1n02x4               g168(.a(new_n263), .b(new_n196), .c(new_n224), .out0(new_n264));
  tech160nm_fioai012aa1n04x5   g169(.a(new_n264), .b(new_n186), .c(new_n183), .o1(new_n265));
  aob012aa1n02x5               g170(.a(new_n251), .b(\b[23] ), .c(\a[24] ), .out0(new_n266));
  oai012aa1n02x5               g171(.a(new_n266), .b(\b[23] ), .c(\a[24] ), .o1(new_n267));
  aoib12aa1n06x5               g172(.a(new_n267), .b(new_n262), .c(new_n246), .out0(new_n268));
  oai012aa1d24x5               g173(.a(new_n268), .b(new_n229), .c(new_n263), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  nanp02aa1n02x5               g175(.a(new_n265), .b(new_n270), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  oai112aa1n02x5               g178(.a(new_n268), .b(new_n273), .c(new_n229), .d(new_n263), .o1(new_n274));
  aboi22aa1n03x5               g179(.a(new_n274), .b(new_n265), .c(new_n271), .d(new_n272), .out0(\s[25] ));
  aoai13aa1n02x5               g180(.a(new_n272), .b(new_n269), .c(new_n214), .d(new_n264), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  orn002aa1n02x5               g182(.a(\a[25] ), .b(\b[24] ), .o(new_n278));
  norb02aa1n02x5               g183(.a(new_n278), .b(new_n277), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n278), .b(new_n273), .c(new_n265), .d(new_n270), .o1(new_n280));
  aoi022aa1n02x5               g185(.a(new_n280), .b(new_n277), .c(new_n276), .d(new_n279), .o1(\s[26] ));
  and002aa1n02x5               g186(.a(new_n277), .b(new_n272), .o(new_n282));
  inv000aa1n02x5               g187(.a(new_n282), .o1(new_n283));
  nor043aa1n06x5               g188(.a(new_n283), .b(new_n225), .c(new_n263), .o1(new_n284));
  oai012aa1n06x5               g189(.a(new_n284), .b(new_n186), .c(new_n183), .o1(new_n285));
  oaoi03aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .c(new_n278), .o1(new_n286));
  aoi012aa1n12x5               g191(.a(new_n286), .b(new_n269), .c(new_n282), .o1(new_n287));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  nanb02aa1n02x5               g194(.a(new_n288), .b(new_n289), .out0(new_n290));
  xobna2aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n287), .out0(\s[27] ));
  oai012aa1n02x5               g196(.a(new_n289), .b(\b[27] ), .c(\a[28] ), .o1(new_n292));
  aoi012aa1n02x5               g197(.a(new_n292), .b(\a[28] ), .c(\b[27] ), .o1(new_n293));
  oaoi13aa1n02x5               g198(.a(new_n283), .b(new_n268), .c(new_n229), .d(new_n263), .o1(new_n294));
  nona32aa1n03x5               g199(.a(new_n285), .b(new_n288), .c(new_n286), .d(new_n294), .out0(new_n295));
  tech160nm_fixnrc02aa1n04x5   g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  nanp02aa1n03x5               g201(.a(new_n295), .b(new_n289), .o1(new_n297));
  aoi022aa1n03x5               g202(.a(new_n297), .b(new_n296), .c(new_n293), .d(new_n295), .o1(\s[28] ));
  inv000aa1n06x5               g203(.a(new_n287), .o1(new_n299));
  nor042aa1n03x5               g204(.a(new_n296), .b(new_n290), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n299), .c(new_n214), .d(new_n284), .o1(new_n301));
  inv000aa1n02x5               g206(.a(new_n300), .o1(new_n302));
  orn002aa1n02x5               g207(.a(\a[27] ), .b(\b[26] ), .o(new_n303));
  oao003aa1n03x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n303), .carry(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n302), .c(new_n285), .d(new_n287), .o1(new_n305));
  xorc02aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n304), .b(new_n306), .out0(new_n307));
  aoi022aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n301), .d(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1d15x5               g214(.a(new_n306), .b(new_n290), .c(new_n296), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n299), .c(new_n214), .d(new_n284), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n310), .o1(new_n312));
  oaoi03aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .o1(new_n313));
  inv000aa1n03x5               g218(.a(new_n313), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n312), .c(new_n285), .d(new_n287), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n304), .b(\a[29] ), .c(\b[28] ), .o1(new_n317));
  oabi12aa1n02x5               g222(.a(new_n316), .b(\a[29] ), .c(\b[28] ), .out0(new_n318));
  norp02aa1n02x5               g223(.a(new_n317), .b(new_n318), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n315), .b(new_n316), .c(new_n311), .d(new_n319), .o1(\s[30] ));
  nano22aa1n06x5               g225(.a(new_n302), .b(new_n306), .c(new_n316), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n299), .c(new_n214), .d(new_n284), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[31] ), .b(\b[30] ), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n314), .carry(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(new_n325));
  inv000aa1d42x5               g230(.a(new_n321), .o1(new_n326));
  aoai13aa1n03x5               g231(.a(new_n324), .b(new_n326), .c(new_n285), .d(new_n287), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n323), .c(new_n322), .d(new_n325), .o1(\s[31] ));
  oai012aa1n02x5               g233(.a(new_n103), .b(new_n109), .c(new_n108), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(new_n329), .b(new_n106), .out0(\s[3] ));
  oaoi03aa1n02x5               g235(.a(\a[3] ), .b(\b[2] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g237(.a(new_n209), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g238(.a(new_n115), .b(new_n114), .out0(new_n334));
  oaoi13aa1n02x5               g239(.a(new_n334), .b(new_n117), .c(new_n209), .d(new_n116), .o1(new_n335));
  oai112aa1n02x5               g240(.a(new_n117), .b(new_n334), .c(new_n209), .d(new_n116), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n336), .b(new_n335), .out0(\s[6] ));
  nanb02aa1n02x5               g242(.a(new_n121), .b(new_n122), .out0(new_n338));
  inv000aa1d42x5               g243(.a(new_n338), .o1(new_n339));
  xnbna2aa1n03x5               g244(.a(new_n339), .b(new_n336), .c(new_n126), .out0(\s[7] ));
  nanb02aa1n02x5               g245(.a(new_n119), .b(new_n120), .out0(new_n341));
  inv000aa1d42x5               g246(.a(new_n121), .o1(new_n342));
  aob012aa1n03x5               g247(.a(new_n339), .b(new_n336), .c(new_n126), .out0(new_n343));
  xobna2aa1n03x5               g248(.a(new_n341), .b(new_n343), .c(new_n342), .out0(\s[8] ));
  xobna2aa1n03x5               g249(.a(new_n132), .b(new_n125), .c(new_n129), .out0(\s[9] ));
endmodule


