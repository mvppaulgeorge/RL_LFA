// Benchmark "adder" written by ABC on Wed Jul 17 19:46:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n314, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n337, new_n338, new_n339,
    new_n340, new_n342, new_n344, new_n345, new_n346, new_n348;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  nor022aa1n08x5               g002(.a(\b[2] ), .b(\a[3] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nand02aa1n03x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oai112aa1n06x5               g005(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n101));
  nanp02aa1n12x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanb02aa1n02x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  aoi113aa1n06x5               g009(.a(new_n104), .b(new_n98), .c(new_n101), .d(new_n99), .e(new_n100), .o1(new_n105));
  nand02aa1d28x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor042aa1n09x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand42aa1n08x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nano22aa1n09x5               g013(.a(new_n107), .b(new_n106), .c(new_n108), .out0(new_n109));
  xorc02aa1n12x5               g014(.a(\a[8] ), .b(\b[7] ), .out0(new_n110));
  nor042aa1d18x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor002aa1n16x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n04x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nano23aa1n06x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .d(new_n102), .out0(new_n114));
  nand23aa1n03x5               g019(.a(new_n114), .b(new_n109), .c(new_n110), .o1(new_n115));
  inv040aa1n09x5               g020(.a(new_n111), .o1(new_n116));
  oai112aa1n06x5               g021(.a(new_n116), .b(new_n106), .c(\b[4] ), .d(\a[5] ), .o1(new_n117));
  aob012aa1n06x5               g022(.a(new_n107), .b(\b[7] ), .c(\a[8] ), .out0(new_n118));
  oai012aa1n02x5               g023(.a(new_n118), .b(\b[7] ), .c(\a[8] ), .o1(new_n119));
  aoi013aa1n09x5               g024(.a(new_n119), .b(new_n109), .c(new_n117), .d(new_n110), .o1(new_n120));
  oai012aa1d24x5               g025(.a(new_n120), .b(new_n115), .c(new_n105), .o1(new_n121));
  xorc02aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .out0(new_n122));
  nand02aa1d06x5               g027(.a(new_n121), .b(new_n122), .o1(new_n123));
  xorc02aa1n02x5               g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  and002aa1n12x5               g029(.a(\b[9] ), .b(\a[10] ), .o(new_n125));
  oai022aa1d18x5               g030(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n126));
  nor042aa1n09x5               g031(.a(new_n126), .b(new_n125), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(new_n123), .b(new_n127), .o1(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n124), .c(new_n97), .d(new_n123), .o1(\s[10] ));
  and002aa1n03x5               g034(.a(\b[10] ), .b(\a[11] ), .o(new_n130));
  nor002aa1d32x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norp02aa1n02x5               g036(.a(new_n130), .b(new_n131), .o1(new_n132));
  inv000aa1n02x5               g037(.a(new_n132), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n125), .c(new_n123), .d(new_n127), .o1(new_n134));
  aoi112aa1n03x5               g039(.a(new_n125), .b(new_n133), .c(new_n123), .d(new_n127), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(\s[11] ));
  nor002aa1d32x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand42aa1d28x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  norb02aa1n06x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  oabi12aa1n03x5               g044(.a(new_n139), .b(new_n135), .c(new_n131), .out0(new_n140));
  nona22aa1n09x5               g045(.a(new_n139), .b(new_n135), .c(new_n131), .out0(new_n141));
  nanp02aa1n03x5               g046(.a(new_n141), .b(new_n140), .o1(\s[12] ));
  nanb02aa1n06x5               g047(.a(new_n98), .b(new_n99), .out0(new_n143));
  nand02aa1d04x5               g048(.a(new_n101), .b(new_n100), .o1(new_n144));
  norb03aa1n03x5               g049(.a(new_n102), .b(new_n98), .c(new_n103), .out0(new_n145));
  oai012aa1n09x5               g050(.a(new_n145), .b(new_n144), .c(new_n143), .o1(new_n146));
  nanb03aa1n02x5               g051(.a(new_n107), .b(new_n108), .c(new_n106), .out0(new_n147));
  xnrc02aa1n02x5               g052(.a(\b[7] ), .b(\a[8] ), .out0(new_n148));
  nor042aa1n02x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  nanp03aa1n09x5               g054(.a(new_n146), .b(new_n149), .c(new_n114), .o1(new_n150));
  and002aa1n02x5               g055(.a(\b[8] ), .b(\a[9] ), .o(new_n151));
  aoi112aa1n06x5               g056(.a(new_n130), .b(new_n131), .c(\a[10] ), .d(\b[9] ), .o1(new_n152));
  nona23aa1n03x5               g057(.a(new_n152), .b(new_n139), .c(new_n151), .d(new_n126), .out0(new_n153));
  aoi022aa1n12x5               g058(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n154));
  nona23aa1d18x5               g059(.a(new_n154), .b(new_n138), .c(new_n131), .d(new_n137), .out0(new_n155));
  aoi012aa1d18x5               g060(.a(new_n137), .b(new_n131), .c(new_n138), .o1(new_n156));
  oai012aa1d24x5               g061(.a(new_n156), .b(new_n155), .c(new_n127), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n153), .c(new_n150), .d(new_n120), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n03x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand02aa1n06x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n06x4               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  nor042aa1n12x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  tech160nm_fiaoi012aa1n05x5   g070(.a(new_n164), .b(new_n159), .c(new_n165), .o1(new_n166));
  xnrc02aa1n02x5               g071(.a(new_n166), .b(new_n163), .out0(\s[14] ));
  nor043aa1n02x5               g072(.a(new_n155), .b(new_n126), .c(new_n151), .o1(new_n168));
  nano23aa1n09x5               g073(.a(new_n164), .b(new_n161), .c(new_n162), .d(new_n165), .out0(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n157), .c(new_n121), .d(new_n168), .o1(new_n170));
  aoi012aa1n12x5               g075(.a(new_n161), .b(new_n164), .c(new_n162), .o1(new_n171));
  nor042aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand02aa1n04x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n171), .out0(\s[15] ));
  nanp02aa1n02x5               g080(.a(new_n170), .b(new_n171), .o1(new_n176));
  nor002aa1n03x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand02aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  aoai13aa1n03x5               g084(.a(new_n179), .b(new_n172), .c(new_n176), .d(new_n174), .o1(new_n180));
  inv030aa1n03x5               g085(.a(new_n171), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n174), .b(new_n181), .c(new_n159), .d(new_n169), .o1(new_n182));
  nona22aa1n03x5               g087(.a(new_n182), .b(new_n179), .c(new_n172), .out0(new_n183));
  nanp02aa1n03x5               g088(.a(new_n180), .b(new_n183), .o1(\s[16] ));
  inv000aa1d42x5               g089(.a(new_n164), .o1(new_n185));
  nona23aa1n09x5               g090(.a(new_n178), .b(new_n173), .c(new_n172), .d(new_n177), .out0(new_n186));
  nano32aa1n03x7               g091(.a(new_n186), .b(new_n163), .c(new_n165), .d(new_n185), .out0(new_n187));
  nand02aa1n02x5               g092(.a(new_n168), .b(new_n187), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n178), .b(new_n177), .c(new_n172), .o1(new_n189));
  oai012aa1n03x5               g094(.a(new_n189), .b(new_n186), .c(new_n171), .o1(new_n190));
  aoi012aa1n06x5               g095(.a(new_n190), .b(new_n157), .c(new_n187), .o1(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n188), .c(new_n150), .d(new_n120), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g098(.a(\a[18] ), .o1(new_n194));
  norp02aa1n02x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  xorc02aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  tech160nm_fiaoi012aa1n05x5   g101(.a(new_n195), .b(new_n192), .c(new_n196), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[17] ), .c(new_n194), .out0(\s[18] ));
  nano23aa1n06x5               g103(.a(new_n172), .b(new_n177), .c(new_n178), .d(new_n173), .out0(new_n199));
  nand22aa1n02x5               g104(.a(new_n199), .b(new_n169), .o1(new_n200));
  nor042aa1n04x5               g105(.a(new_n153), .b(new_n200), .o1(new_n201));
  oai112aa1n02x5               g106(.a(new_n152), .b(new_n139), .c(new_n126), .d(new_n125), .o1(new_n202));
  aobi12aa1n06x5               g107(.a(new_n189), .b(new_n199), .c(new_n181), .out0(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n200), .c(new_n202), .d(new_n156), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\a[17] ), .o1(new_n205));
  xroi22aa1d06x4               g110(.a(new_n205), .b(\b[16] ), .c(new_n194), .d(\b[17] ), .out0(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n204), .c(new_n121), .d(new_n201), .o1(new_n207));
  nor042aa1n02x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  aoi112aa1n09x5               g113(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n209));
  norp02aa1n02x5               g114(.a(new_n209), .b(new_n208), .o1(new_n210));
  nor042aa1n06x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanp02aa1n09x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n09x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n207), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n03x5               g120(.a(new_n207), .b(new_n210), .o1(new_n216));
  nor002aa1n20x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1d28x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1d27x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n04x5               g125(.a(new_n220), .b(new_n211), .c(new_n216), .d(new_n212), .o1(new_n221));
  inv000aa1n02x5               g126(.a(new_n210), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n213), .b(new_n222), .c(new_n192), .d(new_n206), .o1(new_n223));
  nona22aa1n03x5               g128(.a(new_n223), .b(new_n220), .c(new_n211), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n221), .b(new_n224), .o1(\s[20] ));
  nano23aa1n06x5               g130(.a(new_n211), .b(new_n217), .c(new_n218), .d(new_n212), .out0(new_n226));
  nand22aa1n06x5               g131(.a(new_n206), .b(new_n226), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n204), .c(new_n121), .d(new_n201), .o1(new_n229));
  oai112aa1n06x5               g134(.a(new_n213), .b(new_n219), .c(new_n209), .d(new_n208), .o1(new_n230));
  aoi012aa1n12x5               g135(.a(new_n217), .b(new_n211), .c(new_n218), .o1(new_n231));
  nand22aa1n12x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[20] ), .b(\a[21] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n229), .c(new_n233), .out0(\s[21] ));
  nanp02aa1n02x5               g141(.a(new_n229), .b(new_n233), .o1(new_n237));
  nor022aa1n04x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  aoai13aa1n02x5               g144(.a(new_n239), .b(new_n238), .c(new_n237), .d(new_n235), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n235), .b(new_n232), .c(new_n192), .d(new_n228), .o1(new_n241));
  nona22aa1n03x5               g146(.a(new_n241), .b(new_n239), .c(new_n238), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n240), .b(new_n242), .o1(\s[22] ));
  nor042aa1n06x5               g148(.a(new_n239), .b(new_n234), .o1(new_n244));
  and003aa1n02x5               g149(.a(new_n206), .b(new_n244), .c(new_n226), .o(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n204), .c(new_n121), .d(new_n201), .o1(new_n246));
  norp02aa1n02x5               g151(.a(\b[21] ), .b(\a[22] ), .o1(new_n247));
  nanp02aa1n02x5               g152(.a(\b[21] ), .b(\a[22] ), .o1(new_n248));
  aoi012aa1n02x5               g153(.a(new_n247), .b(new_n238), .c(new_n248), .o1(new_n249));
  aobi12aa1n02x5               g154(.a(new_n249), .b(new_n232), .c(new_n244), .out0(new_n250));
  nor002aa1d32x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  nand02aa1d08x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  nanb02aa1d24x5               g157(.a(new_n251), .b(new_n252), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n246), .c(new_n250), .out0(\s[23] ));
  nand02aa1d04x5               g160(.a(new_n246), .b(new_n250), .o1(new_n256));
  nor002aa1d32x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  nand02aa1n04x5               g162(.a(\b[23] ), .b(\a[24] ), .o1(new_n258));
  nanb02aa1n06x5               g163(.a(new_n257), .b(new_n258), .out0(new_n259));
  aoai13aa1n02x7               g164(.a(new_n259), .b(new_n251), .c(new_n256), .d(new_n254), .o1(new_n260));
  tech160nm_finand02aa1n03p5x5 g165(.a(new_n256), .b(new_n254), .o1(new_n261));
  nona22aa1n03x5               g166(.a(new_n261), .b(new_n259), .c(new_n251), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n262), .b(new_n260), .o1(\s[24] ));
  nona23aa1d18x5               g168(.a(new_n258), .b(new_n252), .c(new_n251), .d(new_n257), .out0(new_n264));
  inv040aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  nano22aa1n03x7               g170(.a(new_n227), .b(new_n244), .c(new_n265), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n204), .c(new_n121), .d(new_n201), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n257), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(new_n251), .b(new_n258), .o1(new_n269));
  oai112aa1n02x5               g174(.a(new_n269), .b(new_n268), .c(new_n264), .d(new_n249), .o1(new_n270));
  aoi013aa1n06x4               g175(.a(new_n270), .b(new_n232), .c(new_n244), .d(new_n265), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n267), .c(new_n271), .out0(\s[25] ));
  nand02aa1d06x5               g178(.a(new_n267), .b(new_n271), .o1(new_n274));
  nor042aa1n03x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xnrc02aa1n12x5               g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .d(new_n272), .o1(new_n277));
  tech160nm_finand02aa1n05x5   g182(.a(new_n274), .b(new_n272), .o1(new_n278));
  nona22aa1n03x5               g183(.a(new_n278), .b(new_n276), .c(new_n275), .out0(new_n279));
  nanp02aa1n03x5               g184(.a(new_n279), .b(new_n277), .o1(\s[26] ));
  norb02aa1d21x5               g185(.a(new_n272), .b(new_n276), .out0(new_n281));
  nano32aa1d15x5               g186(.a(new_n227), .b(new_n281), .c(new_n244), .d(new_n265), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n204), .c(new_n121), .d(new_n201), .o1(new_n283));
  inv040aa1n03x5               g188(.a(new_n244), .o1(new_n284));
  aoi112aa1n02x7               g189(.a(new_n284), .b(new_n264), .c(new_n230), .d(new_n231), .o1(new_n285));
  inv000aa1d42x5               g190(.a(\a[26] ), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\b[25] ), .o1(new_n287));
  oao003aa1n02x5               g192(.a(new_n286), .b(new_n287), .c(new_n275), .carry(new_n288));
  oaoi13aa1n06x5               g193(.a(new_n288), .b(new_n281), .c(new_n285), .d(new_n270), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[27] ), .b(\b[26] ), .out0(new_n290));
  xnbna2aa1n03x5               g195(.a(new_n290), .b(new_n289), .c(new_n283), .out0(\s[27] ));
  nanp02aa1n03x5               g196(.a(new_n289), .b(new_n283), .o1(new_n292));
  nor042aa1n03x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[28] ), .b(\b[27] ), .out0(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n293), .c(new_n292), .d(new_n290), .o1(new_n296));
  norp03aa1n02x5               g201(.a(new_n249), .b(new_n253), .c(new_n259), .o1(new_n297));
  nano22aa1n03x7               g202(.a(new_n297), .b(new_n268), .c(new_n269), .out0(new_n298));
  nona32aa1n03x5               g203(.a(new_n232), .b(new_n264), .c(new_n239), .d(new_n234), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n281), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n288), .o1(new_n301));
  aoai13aa1n12x5               g206(.a(new_n301), .b(new_n300), .c(new_n299), .d(new_n298), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n290), .b(new_n302), .c(new_n192), .d(new_n282), .o1(new_n303));
  nona22aa1n03x5               g208(.a(new_n303), .b(new_n295), .c(new_n293), .out0(new_n304));
  nanp02aa1n03x5               g209(.a(new_n296), .b(new_n304), .o1(\s[28] ));
  and002aa1n02x5               g210(.a(new_n294), .b(new_n290), .o(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n302), .c(new_n192), .d(new_n282), .o1(new_n307));
  inv000aa1n03x5               g212(.a(new_n293), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[28] ), .b(\b[27] ), .c(new_n308), .carry(new_n309));
  nanp02aa1n03x5               g214(.a(new_n307), .b(new_n309), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  norb02aa1n02x5               g216(.a(new_n309), .b(new_n311), .out0(new_n312));
  aoi022aa1n02x7               g217(.a(new_n310), .b(new_n311), .c(new_n307), .d(new_n312), .o1(\s[29] ));
  nanp02aa1n02x5               g218(.a(\b[0] ), .b(\a[1] ), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g220(.a(new_n295), .b(new_n290), .c(new_n311), .out0(new_n316));
  aoai13aa1n06x5               g221(.a(new_n316), .b(new_n302), .c(new_n192), .d(new_n282), .o1(new_n317));
  oaoi03aa1n09x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n318), .o1(new_n319));
  nanp02aa1n03x5               g224(.a(new_n317), .b(new_n319), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .out0(new_n321));
  aoi012aa1n02x5               g226(.a(new_n309), .b(\a[29] ), .c(\b[28] ), .o1(new_n322));
  oabi12aa1n02x5               g227(.a(new_n321), .b(\a[29] ), .c(\b[28] ), .out0(new_n323));
  norp02aa1n02x5               g228(.a(new_n322), .b(new_n323), .o1(new_n324));
  aoi022aa1n02x7               g229(.a(new_n320), .b(new_n321), .c(new_n317), .d(new_n324), .o1(\s[30] ));
  and003aa1n02x5               g230(.a(new_n306), .b(new_n321), .c(new_n311), .o(new_n326));
  aoai13aa1n06x5               g231(.a(new_n326), .b(new_n302), .c(new_n192), .d(new_n282), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n319), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  aoi012aa1n03x5               g234(.a(new_n329), .b(new_n327), .c(new_n328), .o1(new_n330));
  aobi12aa1n06x5               g235(.a(new_n326), .b(new_n289), .c(new_n283), .out0(new_n331));
  nano22aa1n03x7               g236(.a(new_n331), .b(new_n328), .c(new_n329), .out0(new_n332));
  nor002aa1n02x5               g237(.a(new_n330), .b(new_n332), .o1(\s[31] ));
  xnbna2aa1n03x5               g238(.a(new_n143), .b(new_n101), .c(new_n100), .out0(\s[3] ));
  aoi013aa1n02x4               g239(.a(new_n98), .b(new_n101), .c(new_n100), .d(new_n99), .o1(new_n335));
  oaib12aa1n02x5               g240(.a(new_n146), .b(new_n335), .c(new_n104), .out0(\s[4] ));
  nano22aa1n02x4               g241(.a(new_n112), .b(new_n102), .c(new_n113), .out0(new_n337));
  nanp02aa1n02x5               g242(.a(new_n146), .b(new_n337), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n112), .o1(new_n339));
  aoi022aa1n02x5               g244(.a(new_n146), .b(new_n102), .c(new_n113), .d(new_n339), .o1(new_n340));
  norb02aa1n02x5               g245(.a(new_n338), .b(new_n340), .out0(\s[5] ));
  ao0022aa1n03x5               g246(.a(new_n338), .b(new_n339), .c(new_n116), .d(new_n106), .o(new_n342));
  oaib12aa1n02x5               g247(.a(new_n342), .b(new_n117), .c(new_n338), .out0(\s[6] ));
  norb02aa1n02x5               g248(.a(new_n108), .b(new_n107), .out0(new_n344));
  aoai13aa1n02x5               g249(.a(new_n109), .b(new_n117), .c(new_n146), .d(new_n337), .o1(new_n345));
  aboi22aa1n03x5               g250(.a(new_n117), .b(new_n338), .c(\a[6] ), .d(\b[5] ), .out0(new_n346));
  oa0012aa1n02x5               g251(.a(new_n345), .b(new_n346), .c(new_n344), .o(\s[7] ));
  orn002aa1n02x5               g252(.a(\a[7] ), .b(\b[6] ), .o(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n110), .b(new_n345), .c(new_n348), .out0(\s[8] ));
  xorb03aa1n02x5               g254(.a(new_n121), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


