// Benchmark "adder" written by ABC on Thu Jul 18 00:35:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n321, new_n322, new_n324, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[2] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[1] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  tech160nm_fioaoi03aa1n02p5x5 g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n02x4               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  aoi012aa1n02x7               g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  tech160nm_fioai012aa1n05x5   g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  norp02aa1n04x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand02aa1n03x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor022aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n06x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  tech160nm_fixorc02aa1n04x5   g017(.a(\a[6] ), .b(\b[5] ), .out0(new_n113));
  tech160nm_fixorc02aa1n03p5x5 g018(.a(\a[5] ), .b(\b[4] ), .out0(new_n114));
  nano22aa1n03x7               g019(.a(new_n112), .b(new_n113), .c(new_n114), .out0(new_n115));
  norp02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  aoi112aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n117));
  norp02aa1n02x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  tech160nm_fiao0012aa1n02p5x5 g023(.a(new_n108), .b(new_n110), .c(new_n109), .o(new_n119));
  oabi12aa1n06x5               g024(.a(new_n119), .b(new_n112), .c(new_n118), .out0(new_n120));
  aoi012aa1n02x5               g025(.a(new_n120), .b(new_n115), .c(new_n107), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .c(new_n121), .o1(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xnrc02aa1n03x5               g028(.a(\b[9] ), .b(\a[10] ), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  nor042aa1n09x5               g030(.a(new_n125), .b(new_n124), .o1(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n120), .c(new_n115), .d(new_n107), .o1(new_n127));
  inv040aa1d32x5               g032(.a(\a[10] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(\b[9] ), .o1(new_n129));
  nor002aa1n03x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  oaoi03aa1n12x5               g035(.a(new_n128), .b(new_n129), .c(new_n130), .o1(new_n131));
  nor002aa1d32x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n127), .c(new_n131), .out0(\s[11] ));
  nanp02aa1n02x5               g040(.a(new_n127), .b(new_n131), .o1(new_n136));
  aoi012aa1n02x5               g041(.a(new_n132), .b(new_n136), .c(new_n133), .o1(new_n137));
  xnrb03aa1n02x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  oao003aa1n02x5               g043(.a(new_n97), .b(new_n98), .c(new_n99), .carry(new_n139));
  nano23aa1n02x5               g044(.a(new_n101), .b(new_n103), .c(new_n104), .d(new_n102), .out0(new_n140));
  aobi12aa1n06x5               g045(.a(new_n106), .b(new_n140), .c(new_n139), .out0(new_n141));
  nanb02aa1n02x5               g046(.a(new_n108), .b(new_n109), .out0(new_n142));
  nanb02aa1n02x5               g047(.a(new_n110), .b(new_n111), .out0(new_n143));
  nona23aa1n09x5               g048(.a(new_n113), .b(new_n114), .c(new_n143), .d(new_n142), .out0(new_n144));
  inv030aa1n06x5               g049(.a(new_n120), .o1(new_n145));
  tech160nm_fioai012aa1n05x5   g050(.a(new_n145), .b(new_n141), .c(new_n144), .o1(new_n146));
  nor002aa1n20x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand22aa1n12x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nano23aa1n06x5               g053(.a(new_n132), .b(new_n147), .c(new_n148), .d(new_n133), .out0(new_n149));
  nona23aa1n09x5               g054(.a(new_n148), .b(new_n133), .c(new_n132), .d(new_n147), .out0(new_n150));
  ao0012aa1n03x7               g055(.a(new_n147), .b(new_n132), .c(new_n148), .o(new_n151));
  oabi12aa1n18x5               g056(.a(new_n151), .b(new_n150), .c(new_n131), .out0(new_n152));
  aoi013aa1n02x4               g057(.a(new_n152), .b(new_n146), .c(new_n126), .d(new_n149), .o1(new_n153));
  nor042aa1n09x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  tech160nm_finand02aa1n03p5x5 g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n153), .b(new_n156), .c(new_n155), .out0(\s[13] ));
  oaoi03aa1n03x5               g062(.a(\a[13] ), .b(\b[12] ), .c(new_n153), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n16x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nand02aa1n06x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nanb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  nor042aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  tech160nm_finand02aa1n03p5x5 g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1d15x5               g069(.a(new_n154), .b(new_n163), .c(new_n164), .d(new_n156), .out0(new_n165));
  nano32aa1n03x7               g070(.a(new_n121), .b(new_n165), .c(new_n126), .d(new_n149), .out0(new_n166));
  tech160nm_fiaoi012aa1n03p5x5 g071(.a(new_n163), .b(new_n154), .c(new_n164), .o1(new_n167));
  aobi12aa1d24x5               g072(.a(new_n167), .b(new_n152), .c(new_n165), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  oabi12aa1n06x5               g074(.a(new_n162), .b(new_n166), .c(new_n169), .out0(new_n170));
  nano22aa1n02x4               g075(.a(new_n166), .b(new_n162), .c(new_n168), .out0(new_n171));
  norb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(\s[15] ));
  inv000aa1d42x5               g077(.a(new_n160), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n170), .c(new_n173), .out0(\s[16] ));
  nona23aa1n09x5               g082(.a(new_n175), .b(new_n161), .c(new_n160), .d(new_n174), .out0(new_n178));
  inv000aa1d42x5               g083(.a(new_n126), .o1(new_n179));
  nano23aa1n02x4               g084(.a(new_n160), .b(new_n174), .c(new_n175), .d(new_n161), .out0(new_n180));
  nano32aa1n03x7               g085(.a(new_n179), .b(new_n180), .c(new_n149), .d(new_n165), .out0(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n120), .c(new_n107), .d(new_n115), .o1(new_n182));
  aoi012aa1n02x5               g087(.a(new_n174), .b(new_n160), .c(new_n175), .o1(new_n183));
  oai112aa1n06x5               g088(.a(new_n182), .b(new_n183), .c(new_n168), .d(new_n178), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g090(.a(\a[18] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  oaoi03aa1n03x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n186), .out0(\s[18] ));
  nona23aa1n09x5               g095(.a(new_n165), .b(new_n126), .c(new_n178), .d(new_n150), .out0(new_n191));
  oaoi13aa1n12x5               g096(.a(new_n191), .b(new_n145), .c(new_n141), .d(new_n144), .o1(new_n192));
  oao003aa1n02x5               g097(.a(new_n128), .b(new_n129), .c(new_n130), .carry(new_n193));
  aoai13aa1n04x5               g098(.a(new_n165), .b(new_n151), .c(new_n149), .d(new_n193), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n183), .b(new_n178), .c(new_n194), .d(new_n167), .o1(new_n195));
  xroi22aa1d04x5               g100(.a(new_n187), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n196));
  tech160nm_fioai012aa1n03p5x5 g101(.a(new_n196), .b(new_n195), .c(new_n192), .o1(new_n197));
  oai022aa1n02x7               g102(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n198));
  oaib12aa1n06x5               g103(.a(new_n198), .b(new_n186), .c(\b[17] ), .out0(new_n199));
  nor002aa1n20x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand42aa1n02x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(new_n200), .b(new_n201), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  xnbna2aa1n03x5               g108(.a(new_n203), .b(new_n197), .c(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(new_n200), .o1(new_n206));
  tech160nm_fiaoi012aa1n02p5x5 g111(.a(new_n202), .b(new_n197), .c(new_n199), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand22aa1n04x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  nano22aa1n03x5               g115(.a(new_n207), .b(new_n206), .c(new_n210), .out0(new_n211));
  nanp02aa1n02x5               g116(.a(new_n188), .b(new_n187), .o1(new_n212));
  oaoi03aa1n02x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n212), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n203), .b(new_n213), .c(new_n184), .d(new_n196), .o1(new_n214));
  aoi012aa1n03x5               g119(.a(new_n210), .b(new_n214), .c(new_n206), .o1(new_n215));
  nor002aa1n02x5               g120(.a(new_n215), .b(new_n211), .o1(\s[20] ));
  nano23aa1n06x5               g121(.a(new_n200), .b(new_n208), .c(new_n209), .d(new_n201), .out0(new_n217));
  nand02aa1d04x5               g122(.a(new_n196), .b(new_n217), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  oaih12aa1n02x5               g124(.a(new_n219), .b(new_n195), .c(new_n192), .o1(new_n220));
  nona23aa1n09x5               g125(.a(new_n209), .b(new_n201), .c(new_n200), .d(new_n208), .out0(new_n221));
  aoi012aa1d18x5               g126(.a(new_n208), .b(new_n200), .c(new_n209), .o1(new_n222));
  oai012aa1d24x5               g127(.a(new_n222), .b(new_n221), .c(new_n199), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n220), .c(new_n224), .out0(\s[21] ));
  orn002aa1n24x5               g131(.a(\a[21] ), .b(\b[20] ), .o(new_n227));
  aobi12aa1n02x5               g132(.a(new_n225), .b(new_n220), .c(new_n224), .out0(new_n228));
  tech160nm_fixnrc02aa1n05x5   g133(.a(\b[21] ), .b(\a[22] ), .out0(new_n229));
  nano22aa1n02x4               g134(.a(new_n228), .b(new_n227), .c(new_n229), .out0(new_n230));
  aoai13aa1n03x5               g135(.a(new_n225), .b(new_n223), .c(new_n184), .d(new_n219), .o1(new_n231));
  aoi012aa1n03x5               g136(.a(new_n229), .b(new_n231), .c(new_n227), .o1(new_n232));
  nor002aa1n02x5               g137(.a(new_n232), .b(new_n230), .o1(\s[22] ));
  nanp02aa1n02x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  nano22aa1n06x5               g139(.a(new_n229), .b(new_n227), .c(new_n234), .out0(new_n235));
  oaoi03aa1n12x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n227), .o1(new_n236));
  tech160nm_fiaoi012aa1n04x5   g141(.a(new_n236), .b(new_n223), .c(new_n235), .o1(new_n237));
  and003aa1n02x5               g142(.a(new_n196), .b(new_n235), .c(new_n217), .o(new_n238));
  tech160nm_fioai012aa1n03p5x5 g143(.a(new_n238), .b(new_n195), .c(new_n192), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[22] ), .b(\a[23] ), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  xnbna2aa1n03x5               g146(.a(new_n241), .b(new_n239), .c(new_n237), .out0(\s[23] ));
  nor042aa1n03x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  tech160nm_fiaoi012aa1n02p5x5 g149(.a(new_n240), .b(new_n239), .c(new_n237), .o1(new_n245));
  xnrc02aa1n02x5               g150(.a(\b[23] ), .b(\a[24] ), .out0(new_n246));
  nano22aa1n02x4               g151(.a(new_n245), .b(new_n244), .c(new_n246), .out0(new_n247));
  inv000aa1n02x5               g152(.a(new_n237), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n241), .b(new_n248), .c(new_n184), .d(new_n238), .o1(new_n249));
  aoi012aa1n03x5               g154(.a(new_n246), .b(new_n249), .c(new_n244), .o1(new_n250));
  nor002aa1n02x5               g155(.a(new_n250), .b(new_n247), .o1(\s[24] ));
  nor042aa1n02x5               g156(.a(new_n246), .b(new_n240), .o1(new_n252));
  nano22aa1n02x5               g157(.a(new_n218), .b(new_n235), .c(new_n252), .out0(new_n253));
  oaih12aa1n02x5               g158(.a(new_n253), .b(new_n195), .c(new_n192), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n222), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n235), .b(new_n255), .c(new_n217), .d(new_n213), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n236), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n252), .o1(new_n258));
  oao003aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n244), .carry(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n258), .c(new_n256), .d(new_n257), .o1(new_n260));
  xnrc02aa1n12x5               g165(.a(\b[24] ), .b(\a[25] ), .out0(new_n261));
  aoib12aa1n03x5               g166(.a(new_n261), .b(new_n254), .c(new_n260), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n261), .o1(new_n263));
  aoi112aa1n02x5               g168(.a(new_n263), .b(new_n260), .c(new_n184), .d(new_n253), .o1(new_n264));
  norp02aa1n02x5               g169(.a(new_n262), .b(new_n264), .o1(\s[25] ));
  nor042aa1n03x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  nano22aa1n02x4               g173(.a(new_n262), .b(new_n267), .c(new_n268), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n263), .b(new_n260), .c(new_n184), .d(new_n253), .o1(new_n270));
  aoi012aa1n03x5               g175(.a(new_n268), .b(new_n270), .c(new_n267), .o1(new_n271));
  nor002aa1n02x5               g176(.a(new_n271), .b(new_n269), .o1(\s[26] ));
  nor042aa1n03x5               g177(.a(new_n268), .b(new_n261), .o1(new_n273));
  nano32aa1n03x7               g178(.a(new_n218), .b(new_n273), .c(new_n235), .d(new_n252), .out0(new_n274));
  oai012aa1n06x5               g179(.a(new_n274), .b(new_n195), .c(new_n192), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .c(new_n267), .carry(new_n276));
  aobi12aa1n06x5               g181(.a(new_n276), .b(new_n260), .c(new_n273), .out0(new_n277));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  nanp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  norb02aa1n02x5               g184(.a(new_n279), .b(new_n278), .out0(new_n280));
  xnbna2aa1n03x5               g185(.a(new_n280), .b(new_n275), .c(new_n277), .out0(\s[27] ));
  inv000aa1n06x5               g186(.a(new_n278), .o1(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n252), .b(new_n236), .c(new_n223), .d(new_n235), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n273), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n276), .b(new_n285), .c(new_n284), .d(new_n259), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n279), .b(new_n286), .c(new_n184), .d(new_n274), .o1(new_n287));
  aoi012aa1n02x7               g192(.a(new_n283), .b(new_n287), .c(new_n282), .o1(new_n288));
  aobi12aa1n02x7               g193(.a(new_n279), .b(new_n275), .c(new_n277), .out0(new_n289));
  nano22aa1n02x4               g194(.a(new_n289), .b(new_n282), .c(new_n283), .out0(new_n290));
  norp02aa1n03x5               g195(.a(new_n288), .b(new_n290), .o1(\s[28] ));
  nano22aa1n02x4               g196(.a(new_n283), .b(new_n282), .c(new_n279), .out0(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n286), .c(new_n184), .d(new_n274), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  aoi012aa1n03x5               g200(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n296));
  aobi12aa1n06x5               g201(.a(new_n292), .b(new_n275), .c(new_n277), .out0(new_n297));
  nano22aa1n02x4               g202(.a(new_n297), .b(new_n294), .c(new_n295), .out0(new_n298));
  nor002aa1n02x5               g203(.a(new_n296), .b(new_n298), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g205(.a(new_n280), .b(new_n295), .c(new_n283), .out0(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n286), .c(new_n184), .d(new_n274), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[29] ), .b(\a[30] ), .out0(new_n304));
  aoi012aa1n03x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  aobi12aa1n02x7               g210(.a(new_n301), .b(new_n275), .c(new_n277), .out0(new_n306));
  nano22aa1n03x5               g211(.a(new_n306), .b(new_n303), .c(new_n304), .out0(new_n307));
  norp02aa1n03x5               g212(.a(new_n305), .b(new_n307), .o1(\s[30] ));
  norb03aa1n02x5               g213(.a(new_n292), .b(new_n304), .c(new_n295), .out0(new_n309));
  aobi12aa1n02x7               g214(.a(new_n309), .b(new_n275), .c(new_n277), .out0(new_n310));
  oao003aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .c(new_n303), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[30] ), .b(\a[31] ), .out0(new_n312));
  nano22aa1n03x5               g217(.a(new_n310), .b(new_n311), .c(new_n312), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n309), .b(new_n286), .c(new_n184), .d(new_n274), .o1(new_n314));
  aoi012aa1n03x5               g219(.a(new_n312), .b(new_n314), .c(new_n311), .o1(new_n315));
  norp02aa1n03x5               g220(.a(new_n315), .b(new_n313), .o1(\s[31] ));
  xnrb03aa1n02x5               g221(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g222(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g224(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai112aa1n02x5               g225(.a(new_n106), .b(new_n114), .c(new_n105), .d(new_n100), .o1(new_n321));
  aob012aa1n02x5               g226(.a(new_n321), .b(\b[4] ), .c(\a[5] ), .out0(new_n322));
  xnrc02aa1n02x5               g227(.a(new_n322), .b(new_n113), .out0(\s[6] ));
  oao003aa1n02x5               g228(.a(\a[6] ), .b(\b[5] ), .c(new_n322), .carry(new_n324));
  xnrb03aa1n02x5               g229(.a(new_n324), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g230(.a(\a[7] ), .b(\b[6] ), .c(new_n324), .o1(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n146), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


