// Benchmark "adder" written by ABC on Wed Jul 17 15:05:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n330,
    new_n332, new_n335, new_n336, new_n337, new_n339, new_n340, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n08x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1n03x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aoi012aa1n06x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n101));
  nor002aa1n06x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand22aa1n03x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n03x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor002aa1d32x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n02x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nanb03aa1n06x5               g012(.a(new_n101), .b(new_n107), .c(new_n104), .out0(new_n108));
  tech160nm_fioai012aa1n03p5x5 g013(.a(new_n103), .b(new_n105), .c(new_n102), .o1(new_n109));
  norp02aa1n04x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanb02aa1n03x5               g016(.a(new_n110), .b(new_n111), .out0(new_n112));
  nand42aa1n16x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanb03aa1d18x5               g020(.a(new_n114), .b(new_n115), .c(new_n113), .out0(new_n116));
  nanp02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nor042aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nor002aa1d32x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  norb03aa1n06x5               g024(.a(new_n113), .b(new_n119), .c(new_n118), .out0(new_n120));
  nona23aa1n02x4               g025(.a(new_n117), .b(new_n120), .c(new_n116), .d(new_n112), .out0(new_n121));
  norp02aa1n02x5               g026(.a(new_n116), .b(new_n112), .o1(new_n122));
  inv040aa1n02x5               g027(.a(new_n119), .o1(new_n123));
  oai112aa1n03x5               g028(.a(new_n123), .b(new_n113), .c(\b[4] ), .d(\a[5] ), .o1(new_n124));
  oai012aa1n02x5               g029(.a(new_n111), .b(new_n114), .c(new_n110), .o1(new_n125));
  aobi12aa1n02x5               g030(.a(new_n125), .b(new_n122), .c(new_n124), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n121), .c(new_n108), .d(new_n109), .o1(new_n127));
  nand42aa1n06x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  aoi012aa1n02x5               g033(.a(new_n97), .b(new_n127), .c(new_n128), .o1(new_n129));
  nor042aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanp02aa1n09x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  norb02aa1n02x5               g037(.a(new_n128), .b(new_n97), .out0(new_n133));
  norb03aa1n09x5               g038(.a(new_n131), .b(new_n97), .c(new_n130), .out0(new_n134));
  aobi12aa1n02x5               g039(.a(new_n134), .b(new_n127), .c(new_n133), .out0(new_n135));
  oabi12aa1n02x5               g040(.a(new_n135), .b(new_n129), .c(new_n132), .out0(\s[10] ));
  nona23aa1n09x5               g041(.a(new_n106), .b(new_n103), .c(new_n102), .d(new_n105), .out0(new_n137));
  oaih12aa1n06x5               g042(.a(new_n109), .b(new_n137), .c(new_n101), .o1(new_n138));
  norb02aa1n03x5               g043(.a(new_n111), .b(new_n110), .out0(new_n139));
  nano23aa1n06x5               g044(.a(new_n124), .b(new_n116), .c(new_n139), .d(new_n117), .out0(new_n140));
  oai013aa1n06x5               g045(.a(new_n125), .b(new_n120), .c(new_n116), .d(new_n112), .o1(new_n141));
  nano23aa1n06x5               g046(.a(new_n97), .b(new_n130), .c(new_n131), .d(new_n128), .out0(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n141), .c(new_n138), .d(new_n140), .o1(new_n143));
  oaib12aa1n02x5               g048(.a(new_n143), .b(new_n134), .c(new_n131), .out0(new_n144));
  xorb03aa1n02x5               g049(.a(new_n144), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n04x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  aoi012aa1n02x5               g052(.a(new_n146), .b(new_n144), .c(new_n147), .o1(new_n148));
  nor042aa1n06x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nand42aa1n08x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  norb02aa1n02x5               g055(.a(new_n150), .b(new_n149), .out0(new_n151));
  norb02aa1n02x5               g056(.a(new_n147), .b(new_n146), .out0(new_n152));
  norb03aa1n03x5               g057(.a(new_n150), .b(new_n146), .c(new_n149), .out0(new_n153));
  aob012aa1n02x5               g058(.a(new_n153), .b(new_n144), .c(new_n152), .out0(new_n154));
  oai012aa1n02x5               g059(.a(new_n154), .b(new_n148), .c(new_n151), .o1(\s[12] ));
  aoi022aa1d24x5               g060(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n156));
  nona23aa1n09x5               g061(.a(new_n156), .b(new_n150), .c(new_n146), .d(new_n149), .out0(new_n157));
  nano22aa1n02x4               g062(.a(new_n157), .b(new_n133), .c(new_n132), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n141), .c(new_n138), .d(new_n140), .o1(new_n159));
  oaih12aa1n02x5               g064(.a(new_n150), .b(new_n149), .c(new_n146), .o1(new_n160));
  oai012aa1n18x5               g065(.a(new_n160), .b(new_n157), .c(new_n134), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nor022aa1n08x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  tech160nm_finand02aa1n05x5   g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  xobna2aa1n03x5               g070(.a(new_n165), .b(new_n159), .c(new_n162), .out0(\s[13] ));
  tech160nm_fiaoi012aa1n05x5   g071(.a(new_n165), .b(new_n159), .c(new_n162), .o1(new_n167));
  nor002aa1n03x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand42aa1n06x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  obai22aa1n02x7               g074(.a(new_n169), .b(new_n168), .c(new_n167), .d(new_n163), .out0(new_n170));
  norb03aa1n02x7               g075(.a(new_n169), .b(new_n163), .c(new_n168), .out0(new_n171));
  oaib12aa1n02x5               g076(.a(new_n170), .b(new_n167), .c(new_n171), .out0(\s[14] ));
  oai012aa1n02x5               g077(.a(new_n169), .b(new_n168), .c(new_n163), .o1(new_n173));
  nona23aa1n03x5               g078(.a(new_n169), .b(new_n164), .c(new_n163), .d(new_n168), .out0(new_n174));
  aoai13aa1n04x5               g079(.a(new_n173), .b(new_n174), .c(new_n159), .d(new_n162), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n04x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nor022aa1n04x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand42aa1n10x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n177), .c(new_n175), .d(new_n178), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n178), .b(new_n177), .out0(new_n183));
  norb03aa1n03x5               g088(.a(new_n180), .b(new_n177), .c(new_n179), .out0(new_n184));
  aob012aa1n02x5               g089(.a(new_n184), .b(new_n175), .c(new_n183), .out0(new_n185));
  nanp02aa1n02x5               g090(.a(new_n182), .b(new_n185), .o1(\s[16] ));
  nano23aa1n03x7               g091(.a(new_n163), .b(new_n168), .c(new_n169), .d(new_n164), .out0(new_n187));
  aoi022aa1d24x5               g092(.a(\b[14] ), .b(\a[15] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n188));
  nand03aa1n02x5               g093(.a(new_n187), .b(new_n184), .c(new_n188), .o1(new_n189));
  nano32aa1n03x7               g094(.a(new_n189), .b(new_n156), .c(new_n142), .d(new_n153), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n141), .c(new_n138), .d(new_n140), .o1(new_n191));
  nona23aa1n03x5               g096(.a(new_n188), .b(new_n180), .c(new_n177), .d(new_n179), .out0(new_n192));
  nor042aa1n02x5               g097(.a(new_n192), .b(new_n174), .o1(new_n193));
  obai22aa1n03x5               g098(.a(new_n180), .b(new_n184), .c(new_n192), .d(new_n171), .out0(new_n194));
  aoi012aa1d18x5               g099(.a(new_n194), .b(new_n161), .c(new_n193), .o1(new_n195));
  tech160nm_fixorc02aa1n04x5   g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n191), .c(new_n195), .out0(\s[17] ));
  nanp02aa1n02x5               g102(.a(new_n191), .b(new_n195), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\a[18] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[17] ), .o1(new_n201));
  nand42aa1n02x5               g106(.a(new_n201), .b(new_n200), .o1(new_n202));
  nand42aa1n03x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n202), .b(new_n203), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n204), .b(new_n199), .c(new_n198), .d(new_n196), .o1(new_n205));
  oai112aa1n03x5               g110(.a(new_n202), .b(new_n203), .c(\b[16] ), .d(\a[17] ), .o1(new_n206));
  aoai13aa1n02x5               g111(.a(new_n205), .b(new_n206), .c(new_n196), .d(new_n198), .o1(\s[18] ));
  norb02aa1n12x5               g112(.a(new_n196), .b(new_n204), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  oaoi03aa1n02x5               g114(.a(new_n200), .b(new_n201), .c(new_n199), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n209), .c(new_n191), .d(new_n195), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nanp02aa1n02x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norp02aa1n12x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand42aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanb02aa1n02x5               g122(.a(new_n216), .b(new_n217), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n214), .c(new_n211), .d(new_n215), .o1(new_n219));
  inv040aa1n08x5               g124(.a(new_n195), .o1(new_n220));
  aoai13aa1n02x5               g125(.a(new_n208), .b(new_n220), .c(new_n127), .d(new_n190), .o1(new_n221));
  nanb02aa1n02x5               g126(.a(new_n214), .b(new_n215), .out0(new_n222));
  norb03aa1n03x5               g127(.a(new_n217), .b(new_n214), .c(new_n216), .out0(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n222), .c(new_n221), .d(new_n210), .o1(new_n224));
  nanp02aa1n02x5               g129(.a(new_n219), .b(new_n224), .o1(\s[20] ));
  aoi022aa1n06x5               g130(.a(\b[18] ), .b(\a[19] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n226));
  nona23aa1n06x5               g131(.a(new_n226), .b(new_n217), .c(new_n214), .d(new_n216), .out0(new_n227));
  norb03aa1n03x5               g132(.a(new_n196), .b(new_n227), .c(new_n204), .out0(new_n228));
  inv040aa1n03x5               g133(.a(new_n228), .o1(new_n229));
  tech160nm_fioai012aa1n04x5   g134(.a(new_n217), .b(new_n216), .c(new_n214), .o1(new_n230));
  oaib12aa1n09x5               g135(.a(new_n230), .b(new_n227), .c(new_n206), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n229), .c(new_n191), .d(new_n195), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nanp02aa1n02x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  nor002aa1d32x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nand42aa1d28x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nanb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n235), .c(new_n233), .d(new_n237), .o1(new_n241));
  nanp02aa1n02x5               g146(.a(new_n233), .b(new_n237), .o1(new_n242));
  inv040aa1n09x5               g147(.a(new_n238), .o1(new_n243));
  oai112aa1n06x5               g148(.a(new_n243), .b(new_n239), .c(\b[20] ), .d(\a[21] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  nanp02aa1n02x5               g150(.a(new_n242), .b(new_n245), .o1(new_n246));
  nanp02aa1n02x5               g151(.a(new_n241), .b(new_n246), .o1(\s[22] ));
  nano23aa1n03x7               g152(.a(new_n235), .b(new_n238), .c(new_n239), .d(new_n236), .out0(new_n248));
  nano23aa1n02x4               g153(.a(new_n227), .b(new_n204), .c(new_n248), .d(new_n196), .out0(new_n249));
  inv000aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  aoi022aa1n06x5               g155(.a(new_n231), .b(new_n248), .c(new_n239), .d(new_n244), .o1(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n250), .c(new_n191), .d(new_n195), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  norp02aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nand42aa1n03x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  nanb02aa1n03x5               g162(.a(new_n256), .b(new_n257), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n254), .c(new_n252), .d(new_n255), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n249), .b(new_n220), .c(new_n127), .d(new_n190), .o1(new_n260));
  nanb02aa1n02x5               g165(.a(new_n254), .b(new_n255), .out0(new_n261));
  norb03aa1n03x5               g166(.a(new_n257), .b(new_n254), .c(new_n256), .out0(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n261), .c(new_n260), .d(new_n251), .o1(new_n263));
  nanp02aa1n03x5               g168(.a(new_n259), .b(new_n263), .o1(\s[24] ));
  inv000aa1n02x5               g169(.a(new_n254), .o1(new_n265));
  aoi022aa1n12x5               g170(.a(\b[22] ), .b(\a[23] ), .c(\a[22] ), .d(\b[21] ), .o1(new_n266));
  nano22aa1n02x4               g171(.a(new_n258), .b(new_n266), .c(new_n265), .out0(new_n267));
  nand02aa1n02x5               g172(.a(new_n267), .b(new_n248), .o1(new_n268));
  nanb02aa1n02x5               g173(.a(new_n268), .b(new_n228), .out0(new_n269));
  nanp03aa1n02x5               g174(.a(new_n206), .b(new_n223), .c(new_n226), .o1(new_n270));
  oaoi03aa1n02x5               g175(.a(\a[24] ), .b(\b[23] ), .c(new_n265), .o1(new_n271));
  aoi013aa1n06x4               g176(.a(new_n271), .b(new_n244), .c(new_n262), .d(new_n266), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n268), .c(new_n270), .d(new_n230), .o1(new_n273));
  inv000aa1n02x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n269), .c(new_n191), .d(new_n195), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  tech160nm_fixorc02aa1n05x5   g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(new_n275), .b(new_n278), .o1(new_n281));
  oabi12aa1n06x5               g186(.a(new_n279), .b(\a[25] ), .c(\b[24] ), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n281), .b(new_n283), .o1(new_n284));
  nanp02aa1n02x5               g189(.a(new_n280), .b(new_n284), .o1(\s[26] ));
  norb02aa1n02x5               g190(.a(new_n278), .b(new_n279), .out0(new_n286));
  nano32aa1n03x7               g191(.a(new_n229), .b(new_n286), .c(new_n248), .d(new_n267), .out0(new_n287));
  inv000aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[25] ), .b(\a[26] ), .o1(new_n289));
  aoi022aa1n09x5               g194(.a(new_n273), .b(new_n286), .c(new_n289), .d(new_n282), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n288), .c(new_n191), .d(new_n195), .o1(new_n291));
  xorb03aa1n03x5               g196(.a(new_n291), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  xnrc02aa1n12x5               g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n293), .c(new_n291), .d(new_n294), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n287), .b(new_n220), .c(new_n127), .d(new_n190), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n294), .o1(new_n298));
  norp02aa1n02x5               g203(.a(new_n295), .b(new_n293), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n297), .d(new_n290), .o1(new_n300));
  nanp02aa1n03x5               g205(.a(new_n296), .b(new_n300), .o1(\s[28] ));
  xorc02aa1n12x5               g206(.a(\a[29] ), .b(\b[28] ), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  norb02aa1n06x5               g208(.a(new_n294), .b(new_n295), .out0(new_n304));
  aoi012aa1n02x5               g209(.a(new_n299), .b(\a[28] ), .c(\b[27] ), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n303), .b(new_n305), .c(new_n291), .d(new_n304), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n304), .o1(new_n307));
  norp02aa1n02x5               g212(.a(new_n305), .b(new_n303), .o1(new_n308));
  aoai13aa1n02x5               g213(.a(new_n308), .b(new_n307), .c(new_n297), .d(new_n290), .o1(new_n309));
  nanp02aa1n03x5               g214(.a(new_n306), .b(new_n309), .o1(\s[29] ));
  xorb03aa1n02x5               g215(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g216(.a(new_n295), .b(new_n294), .c(new_n302), .out0(new_n312));
  nanp02aa1n03x5               g217(.a(new_n291), .b(new_n312), .o1(new_n313));
  norp02aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .o1(new_n314));
  aoi012aa1n02x5               g219(.a(new_n314), .b(new_n305), .c(new_n302), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .out0(new_n316));
  inv000aa1n02x5               g221(.a(new_n312), .o1(new_n317));
  oai012aa1n02x5               g222(.a(new_n316), .b(\b[28] ), .c(\a[29] ), .o1(new_n318));
  aoi012aa1n03x5               g223(.a(new_n318), .b(new_n305), .c(new_n302), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n317), .c(new_n297), .d(new_n290), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n316), .c(new_n313), .d(new_n315), .o1(\s[30] ));
  nano23aa1d12x5               g226(.a(new_n303), .b(new_n295), .c(new_n316), .d(new_n294), .out0(new_n322));
  aoi012aa1n02x5               g227(.a(new_n319), .b(\a[30] ), .c(\b[29] ), .o1(new_n323));
  xnrc02aa1n02x5               g228(.a(\b[30] ), .b(\a[31] ), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n323), .c(new_n291), .d(new_n322), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n322), .o1(new_n326));
  norp02aa1n02x5               g231(.a(new_n323), .b(new_n324), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n326), .c(new_n297), .d(new_n290), .o1(new_n328));
  nanp02aa1n03x5               g233(.a(new_n325), .b(new_n328), .o1(\s[31] ));
  inv000aa1d42x5               g234(.a(new_n105), .o1(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n101), .b(new_n106), .c(new_n330), .out0(\s[3] ));
  aoai13aa1n02x5               g236(.a(new_n107), .b(new_n98), .c(new_n100), .d(new_n99), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n104), .b(new_n332), .c(new_n330), .out0(\s[4] ));
  xorb03aa1n02x5               g238(.a(new_n138), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g239(.a(new_n118), .b(new_n138), .c(new_n117), .o1(new_n335));
  nanb02aa1n02x5               g240(.a(new_n118), .b(new_n117), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n120), .b(new_n336), .c(new_n108), .d(new_n109), .o1(new_n337));
  aoai13aa1n02x5               g242(.a(new_n337), .b(new_n335), .c(new_n113), .d(new_n123), .o1(\s[6] ));
  nanb02aa1n02x5               g243(.a(new_n116), .b(new_n337), .out0(new_n339));
  inv000aa1d42x5               g244(.a(new_n114), .o1(new_n340));
  aoi022aa1n02x5               g245(.a(new_n337), .b(new_n113), .c(new_n340), .d(new_n115), .o1(new_n341));
  norb02aa1n02x5               g246(.a(new_n339), .b(new_n341), .out0(\s[7] ));
  xnbna2aa1n03x5               g247(.a(new_n139), .b(new_n339), .c(new_n340), .out0(\s[8] ));
  xorb03aa1n02x5               g248(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


