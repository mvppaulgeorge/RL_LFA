// Benchmark "adder" written by ABC on Thu Jul 18 06:15:43 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n334, new_n335, new_n338, new_n339, new_n341,
    new_n342, new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  and002aa1n12x5               g002(.a(\b[1] ), .b(\a[2] ), .o(new_n98));
  nand02aa1d04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oab012aa1n06x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .out0(new_n101));
  nor022aa1n08x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  norb02aa1n02x7               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor002aa1d32x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nand22aa1n06x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb02aa1d21x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nand03aa1n03x5               g012(.a(new_n101), .b(new_n104), .c(new_n107), .o1(new_n108));
  tech160nm_fiaoi012aa1n05x5   g013(.a(new_n105), .b(new_n102), .c(new_n106), .o1(new_n109));
  nand42aa1n08x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor022aa1n06x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  norp02aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand42aa1n08x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nano23aa1n02x4               g018(.a(new_n112), .b(new_n111), .c(new_n113), .d(new_n110), .out0(new_n114));
  tech160nm_fixorc02aa1n02p5x5 g019(.a(\a[5] ), .b(\b[4] ), .out0(new_n115));
  norp02aa1n06x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nanp02aa1n12x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  norb02aa1n09x5               g022(.a(new_n117), .b(new_n116), .out0(new_n118));
  nanp03aa1n02x5               g023(.a(new_n114), .b(new_n115), .c(new_n118), .o1(new_n119));
  nano22aa1n02x4               g024(.a(new_n111), .b(new_n110), .c(new_n113), .out0(new_n120));
  oai022aa1n02x5               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  oa0012aa1n02x5               g026(.a(new_n117), .b(new_n116), .c(new_n111), .o(new_n122));
  aoi013aa1n03x5               g027(.a(new_n122), .b(new_n120), .c(new_n121), .d(new_n118), .o1(new_n123));
  aoai13aa1n06x5               g028(.a(new_n123), .b(new_n119), .c(new_n108), .d(new_n109), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoi012aa1n02x5               g030(.a(new_n97), .b(new_n124), .c(new_n125), .o1(new_n126));
  nor002aa1d32x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nanp02aa1n12x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n15x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nona22aa1n02x4               g034(.a(new_n128), .b(new_n127), .c(new_n97), .out0(new_n130));
  tech160nm_fiao0012aa1n02p5x5 g035(.a(new_n130), .b(new_n124), .c(new_n125), .o(new_n131));
  oai012aa1n02x5               g036(.a(new_n131), .b(new_n126), .c(new_n129), .o1(\s[10] ));
  nand42aa1d28x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor002aa1d24x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nano22aa1n02x4               g039(.a(new_n134), .b(new_n128), .c(new_n133), .out0(new_n135));
  inv000aa1d42x5               g040(.a(\b[10] ), .o1(new_n136));
  nanb02aa1d24x5               g041(.a(\a[11] ), .b(new_n136), .out0(new_n137));
  nanp02aa1n02x5               g042(.a(new_n137), .b(new_n133), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n128), .b(new_n130), .c(new_n124), .d(new_n125), .o1(new_n139));
  aoi022aa1n02x5               g044(.a(new_n131), .b(new_n135), .c(new_n139), .d(new_n138), .o1(\s[11] ));
  aoai13aa1n02x5               g045(.a(new_n135), .b(new_n130), .c(new_n124), .d(new_n125), .o1(new_n141));
  nor002aa1n16x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d28x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  xobna2aa1n03x5               g049(.a(new_n144), .b(new_n141), .c(new_n137), .out0(\s[12] ));
  oabi12aa1n06x5               g050(.a(new_n98), .b(new_n99), .c(new_n100), .out0(new_n146));
  nona23aa1n03x5               g051(.a(new_n106), .b(new_n103), .c(new_n102), .d(new_n105), .out0(new_n147));
  oai012aa1n12x5               g052(.a(new_n109), .b(new_n147), .c(new_n146), .o1(new_n148));
  nona23aa1n03x5               g053(.a(new_n110), .b(new_n113), .c(new_n112), .d(new_n111), .out0(new_n149));
  nano22aa1n03x7               g054(.a(new_n149), .b(new_n115), .c(new_n118), .out0(new_n150));
  nand43aa1n03x5               g055(.a(new_n120), .b(new_n118), .c(new_n121), .o1(new_n151));
  nanb02aa1n06x5               g056(.a(new_n122), .b(new_n151), .out0(new_n152));
  nano23aa1d15x5               g057(.a(new_n142), .b(new_n134), .c(new_n143), .d(new_n133), .out0(new_n153));
  nand23aa1d12x5               g058(.a(new_n153), .b(new_n125), .c(new_n129), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n152), .c(new_n148), .d(new_n150), .o1(new_n156));
  nona23aa1n03x5               g061(.a(new_n133), .b(new_n143), .c(new_n142), .d(new_n134), .out0(new_n157));
  oai112aa1n06x5               g062(.a(new_n137), .b(new_n128), .c(new_n127), .d(new_n97), .o1(new_n158));
  oaoi03aa1n09x5               g063(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .o1(new_n159));
  oabi12aa1n06x5               g064(.a(new_n159), .b(new_n157), .c(new_n158), .out0(new_n160));
  inv000aa1n02x5               g065(.a(new_n160), .o1(new_n161));
  nor042aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  tech160nm_finand02aa1n03p5x5 g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n06x4               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n156), .c(new_n161), .out0(\s[13] ));
  orn002aa1n02x5               g070(.a(\a[13] ), .b(\b[12] ), .o(new_n166));
  aoai13aa1n03x5               g071(.a(new_n164), .b(new_n160), .c(new_n124), .d(new_n155), .o1(new_n167));
  nor042aa1n04x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand22aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n03x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  xnbna2aa1n03x5               g075(.a(new_n170), .b(new_n167), .c(new_n166), .out0(\s[14] ));
  nona23aa1n09x5               g076(.a(new_n169), .b(new_n163), .c(new_n162), .d(new_n168), .out0(new_n172));
  aoi012aa1n02x5               g077(.a(new_n168), .b(new_n162), .c(new_n169), .o1(new_n173));
  aoai13aa1n06x5               g078(.a(new_n173), .b(new_n172), .c(new_n156), .d(new_n161), .o1(new_n174));
  xorb03aa1n02x5               g079(.a(new_n174), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n09x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nanp02aa1n04x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nor042aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand42aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n176), .c(new_n174), .d(new_n177), .o1(new_n181));
  aoi112aa1n03x4               g086(.a(new_n176), .b(new_n180), .c(new_n174), .d(new_n177), .o1(new_n182));
  nanb02aa1n03x5               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano23aa1n06x5               g088(.a(new_n176), .b(new_n178), .c(new_n179), .d(new_n177), .out0(new_n184));
  nano32aa1d12x5               g089(.a(new_n154), .b(new_n184), .c(new_n164), .d(new_n170), .out0(new_n185));
  aoai13aa1n12x5               g090(.a(new_n185), .b(new_n152), .c(new_n150), .d(new_n148), .o1(new_n186));
  nona23aa1n03x5               g091(.a(new_n179), .b(new_n177), .c(new_n176), .d(new_n178), .out0(new_n187));
  nor022aa1n04x5               g092(.a(new_n187), .b(new_n172), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n176), .o1(new_n189));
  aoai13aa1n06x5               g094(.a(new_n177), .b(new_n168), .c(new_n162), .d(new_n169), .o1(new_n190));
  aoi022aa1n06x5               g095(.a(new_n190), .b(new_n189), .c(\a[16] ), .d(\b[15] ), .o1(new_n191));
  aoi112aa1n09x5               g096(.a(new_n178), .b(new_n191), .c(new_n160), .d(new_n188), .o1(new_n192));
  xorc02aa1n12x5               g097(.a(\a[17] ), .b(\b[16] ), .out0(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n193), .b(new_n186), .c(new_n192), .out0(\s[17] ));
  inv000aa1d42x5               g099(.a(\a[17] ), .o1(new_n195));
  inv000aa1d42x5               g100(.a(\b[16] ), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n196), .b(new_n195), .o1(new_n197));
  inv000aa1n02x5               g102(.a(new_n158), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n188), .b(new_n159), .c(new_n198), .d(new_n153), .o1(new_n199));
  nor042aa1n02x5               g104(.a(new_n191), .b(new_n178), .o1(new_n200));
  nanp02aa1n04x5               g105(.a(new_n199), .b(new_n200), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n193), .b(new_n201), .c(new_n124), .d(new_n185), .o1(new_n202));
  nor042aa1n06x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand02aa1d06x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nanb02aa1n09x5               g109(.a(new_n203), .b(new_n204), .out0(new_n205));
  xobna2aa1n03x5               g110(.a(new_n205), .b(new_n202), .c(new_n197), .out0(\s[18] ));
  norb02aa1n02x5               g111(.a(new_n193), .b(new_n205), .out0(new_n207));
  inv000aa1n02x5               g112(.a(new_n207), .o1(new_n208));
  aoi013aa1n06x4               g113(.a(new_n203), .b(new_n204), .c(new_n195), .d(new_n196), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n208), .c(new_n186), .d(new_n192), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n16x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand42aa1n08x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nor002aa1d24x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nand42aa1d28x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  norb02aa1n15x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n213), .c(new_n210), .d(new_n214), .o1(new_n219));
  norb02aa1n06x4               g124(.a(new_n214), .b(new_n213), .out0(new_n220));
  nanp02aa1n03x5               g125(.a(new_n210), .b(new_n220), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n218), .c(new_n213), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n222), .b(new_n219), .o1(\s[20] ));
  nano23aa1n03x7               g128(.a(new_n213), .b(new_n215), .c(new_n216), .d(new_n214), .out0(new_n224));
  nanb03aa1n02x5               g129(.a(new_n205), .b(new_n224), .c(new_n193), .out0(new_n225));
  nona23aa1d18x5               g130(.a(new_n216), .b(new_n214), .c(new_n213), .d(new_n215), .out0(new_n226));
  oaih12aa1n12x5               g131(.a(new_n216), .b(new_n215), .c(new_n213), .o1(new_n227));
  oai012aa1n18x5               g132(.a(new_n227), .b(new_n226), .c(new_n209), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n225), .c(new_n186), .d(new_n192), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  tech160nm_finor002aa1n03p5x5 g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[20] ), .b(\a[21] ), .out0(new_n233));
  inv000aa1n02x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[21] ), .b(\a[22] ), .out0(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n232), .c(new_n230), .d(new_n234), .o1(new_n236));
  nanp02aa1n03x5               g141(.a(new_n230), .b(new_n234), .o1(new_n237));
  nona22aa1n02x5               g142(.a(new_n237), .b(new_n235), .c(new_n232), .out0(new_n238));
  nanp02aa1n03x5               g143(.a(new_n238), .b(new_n236), .o1(\s[22] ));
  nor002aa1n03x5               g144(.a(new_n235), .b(new_n233), .o1(new_n240));
  nona23aa1d18x5               g145(.a(new_n240), .b(new_n193), .c(new_n226), .d(new_n205), .out0(new_n241));
  aoi112aa1n03x5               g146(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n242));
  oai112aa1n06x5               g147(.a(new_n220), .b(new_n217), .c(new_n242), .d(new_n203), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(new_n235), .b(new_n234), .out0(new_n244));
  inv000aa1d42x5               g149(.a(\a[22] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\b[21] ), .o1(new_n246));
  oaoi03aa1n09x5               g151(.a(new_n245), .b(new_n246), .c(new_n232), .o1(new_n247));
  aoai13aa1n12x5               g152(.a(new_n247), .b(new_n244), .c(new_n243), .d(new_n227), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n241), .c(new_n186), .d(new_n192), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  xnrc02aa1n03x5               g158(.a(\b[23] ), .b(\a[24] ), .out0(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n252), .c(new_n250), .d(new_n253), .o1(new_n255));
  nanp02aa1n03x5               g160(.a(new_n250), .b(new_n253), .o1(new_n256));
  nona22aa1n02x5               g161(.a(new_n256), .b(new_n254), .c(new_n252), .out0(new_n257));
  nanp02aa1n03x5               g162(.a(new_n257), .b(new_n255), .o1(\s[24] ));
  norb02aa1n03x5               g163(.a(new_n253), .b(new_n254), .out0(new_n259));
  nanb03aa1n02x5               g164(.a(new_n225), .b(new_n259), .c(new_n240), .out0(new_n260));
  oaoi03aa1n02x5               g165(.a(\a[18] ), .b(\b[17] ), .c(new_n197), .o1(new_n261));
  inv040aa1n03x5               g166(.a(new_n227), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n240), .b(new_n262), .c(new_n224), .d(new_n261), .o1(new_n263));
  inv000aa1n02x5               g168(.a(new_n259), .o1(new_n264));
  inv000aa1d42x5               g169(.a(\a[24] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(\b[23] ), .o1(new_n266));
  oao003aa1n02x5               g171(.a(new_n265), .b(new_n266), .c(new_n252), .carry(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n264), .c(new_n263), .d(new_n247), .o1(new_n269));
  inv040aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n260), .c(new_n186), .d(new_n192), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  tech160nm_fixorc02aa1n04x5   g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xorc02aa1n12x5               g179(.a(\a[26] ), .b(\b[25] ), .out0(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n277));
  nanp02aa1n03x5               g182(.a(new_n271), .b(new_n274), .o1(new_n278));
  nona22aa1n02x5               g183(.a(new_n278), .b(new_n276), .c(new_n273), .out0(new_n279));
  nanp02aa1n03x5               g184(.a(new_n279), .b(new_n277), .o1(\s[26] ));
  and002aa1n12x5               g185(.a(new_n275), .b(new_n274), .o(new_n281));
  nano22aa1n03x7               g186(.a(new_n241), .b(new_n259), .c(new_n281), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n201), .c(new_n124), .d(new_n185), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(\b[25] ), .b(\a[26] ), .o1(new_n284));
  oai022aa1n02x5               g189(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n285));
  aoi022aa1n06x5               g190(.a(new_n269), .b(new_n281), .c(new_n284), .d(new_n285), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[27] ), .b(\b[26] ), .out0(new_n287));
  xnbna2aa1n03x5               g192(.a(new_n287), .b(new_n286), .c(new_n283), .out0(\s[27] ));
  aoai13aa1n04x5               g193(.a(new_n281), .b(new_n267), .c(new_n248), .d(new_n259), .o1(new_n289));
  nanp02aa1n02x5               g194(.a(new_n285), .b(new_n284), .o1(new_n290));
  nanp03aa1n03x5               g195(.a(new_n283), .b(new_n289), .c(new_n290), .o1(new_n291));
  norp02aa1n02x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  norp02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .o1(new_n293));
  nand02aa1d04x5               g198(.a(\b[27] ), .b(\a[28] ), .o1(new_n294));
  nanb02aa1n06x5               g199(.a(new_n293), .b(new_n294), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n292), .c(new_n291), .d(new_n287), .o1(new_n296));
  aobi12aa1n06x5               g201(.a(new_n282), .b(new_n186), .c(new_n192), .out0(new_n297));
  inv000aa1n02x5               g202(.a(new_n247), .o1(new_n298));
  aoai13aa1n02x7               g203(.a(new_n259), .b(new_n298), .c(new_n228), .d(new_n240), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n281), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n290), .b(new_n300), .c(new_n299), .d(new_n268), .o1(new_n301));
  oaih12aa1n02x5               g206(.a(new_n287), .b(new_n301), .c(new_n297), .o1(new_n302));
  nona22aa1n02x5               g207(.a(new_n302), .b(new_n295), .c(new_n292), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n296), .b(new_n303), .o1(\s[28] ));
  norb02aa1n03x5               g209(.a(new_n287), .b(new_n295), .out0(new_n305));
  oaih12aa1n02x5               g210(.a(new_n305), .b(new_n301), .c(new_n297), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n305), .o1(new_n307));
  aoi012aa1n02x5               g212(.a(new_n293), .b(new_n292), .c(new_n294), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n307), .c(new_n286), .d(new_n283), .o1(new_n309));
  xorc02aa1n12x5               g214(.a(\a[29] ), .b(\b[28] ), .out0(new_n310));
  norb02aa1n02x5               g215(.a(new_n308), .b(new_n310), .out0(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n306), .d(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g217(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g218(.a(new_n295), .b(new_n287), .c(new_n310), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n314), .b(new_n301), .c(new_n297), .o1(new_n315));
  inv000aa1n02x5               g220(.a(new_n314), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .carry(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n316), .c(new_n286), .d(new_n283), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n317), .b(new_n319), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n315), .d(new_n320), .o1(\s[30] ));
  nanp03aa1n02x5               g226(.a(new_n305), .b(new_n310), .c(new_n319), .o1(new_n322));
  oabi12aa1n03x5               g227(.a(new_n322), .b(new_n301), .c(new_n297), .out0(new_n323));
  xorc02aa1n02x5               g228(.a(\a[31] ), .b(\b[30] ), .out0(new_n324));
  inv000aa1d42x5               g229(.a(\a[30] ), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[29] ), .o1(new_n326));
  inv000aa1n02x5               g231(.a(new_n317), .o1(new_n327));
  oabi12aa1n02x5               g232(.a(new_n324), .b(\a[30] ), .c(\b[29] ), .out0(new_n328));
  oaoi13aa1n02x5               g233(.a(new_n328), .b(new_n327), .c(new_n325), .d(new_n326), .o1(new_n329));
  oaoi03aa1n02x5               g234(.a(new_n325), .b(new_n326), .c(new_n327), .o1(new_n330));
  aoai13aa1n02x7               g235(.a(new_n330), .b(new_n322), .c(new_n286), .d(new_n283), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n331), .b(new_n324), .c(new_n323), .d(new_n329), .o1(\s[31] ));
  xorb03aa1n02x5               g237(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g238(.a(new_n107), .o1(new_n334));
  oai112aa1n02x5               g239(.a(new_n103), .b(new_n334), .c(new_n101), .d(new_n102), .o1(new_n335));
  oai012aa1n02x5               g240(.a(new_n335), .b(new_n148), .c(new_n334), .o1(\s[4] ));
  xorb03aa1n02x5               g241(.a(new_n148), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  and002aa1n02x5               g242(.a(\b[4] ), .b(\a[5] ), .o(new_n338));
  aoi013aa1n03x5               g243(.a(new_n338), .b(new_n108), .c(new_n109), .d(new_n115), .o1(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g245(.a(\a[7] ), .o1(new_n341));
  oai012aa1n02x5               g246(.a(new_n113), .b(new_n339), .c(new_n112), .o1(new_n342));
  xorb03aa1n02x5               g247(.a(new_n342), .b(\b[6] ), .c(new_n341), .out0(\s[7] ));
  oaib12aa1n03x5               g248(.a(new_n342), .b(\b[6] ), .c(new_n341), .out0(new_n344));
  xobna2aa1n03x5               g249(.a(new_n118), .b(new_n344), .c(new_n110), .out0(\s[8] ));
  xorb03aa1n02x5               g250(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


