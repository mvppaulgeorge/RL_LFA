// Benchmark "adder" written by ABC on Wed Jul 17 17:56:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n315, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n337, new_n338,
    new_n340, new_n342, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n09x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  nor042aa1n06x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  norp02aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nor002aa1n02x5               g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanb02aa1n09x5               g007(.a(new_n99), .b(new_n102), .out0(new_n103));
  nand42aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oai112aa1n06x5               g009(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n105));
  nanp02aa1n06x5               g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n101), .b(new_n106), .c(new_n103), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand42aa1n04x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nor042aa1d18x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nanb03aa1d18x5               g015(.a(new_n110), .b(new_n108), .c(new_n109), .out0(new_n111));
  aoi022aa1d24x5               g016(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n112));
  inv030aa1d32x5               g017(.a(\a[8] ), .o1(new_n113));
  inv030aa1n06x5               g018(.a(\b[7] ), .o1(new_n114));
  nor002aa1n10x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  aoi012aa1n02x7               g020(.a(new_n115), .b(new_n113), .c(new_n114), .o1(new_n116));
  inv040aa1d32x5               g021(.a(\a[7] ), .o1(new_n117));
  inv040aa1d28x5               g022(.a(\b[6] ), .o1(new_n118));
  nand22aa1n03x5               g023(.a(new_n118), .b(new_n117), .o1(new_n119));
  nand42aa1n03x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(new_n119), .b(new_n120), .o1(new_n121));
  nano23aa1n06x5               g026(.a(new_n111), .b(new_n121), .c(new_n116), .d(new_n112), .out0(new_n122));
  nanp02aa1n02x5               g027(.a(new_n114), .b(new_n113), .o1(new_n123));
  tech160nm_finand02aa1n05x5   g028(.a(\b[5] ), .b(\a[6] ), .o1(new_n124));
  tech160nm_fioai012aa1n05x5   g029(.a(new_n124), .b(new_n115), .c(new_n110), .o1(new_n125));
  aob012aa1n02x5               g030(.a(new_n120), .b(\b[7] ), .c(\a[8] ), .out0(new_n126));
  aoai13aa1n04x5               g031(.a(new_n123), .b(new_n126), .c(new_n125), .d(new_n119), .o1(new_n127));
  tech160nm_fixorc02aa1n05x5   g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n122), .d(new_n107), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g036(.a(\a[11] ), .o1(new_n132));
  aoi113aa1n02x5               g037(.a(new_n100), .b(new_n99), .c(new_n105), .d(new_n104), .e(new_n102), .o1(new_n133));
  nano22aa1n02x4               g038(.a(new_n110), .b(new_n108), .c(new_n109), .out0(new_n134));
  inv000aa1d42x5               g039(.a(new_n112), .o1(new_n135));
  nona23aa1n02x4               g040(.a(new_n116), .b(new_n134), .c(new_n121), .d(new_n135), .out0(new_n136));
  oabi12aa1n06x5               g041(.a(new_n127), .b(new_n136), .c(new_n133), .out0(new_n137));
  nand02aa1d06x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  tech160nm_fixnrc02aa1n04x5   g043(.a(\b[9] ), .b(\a[10] ), .out0(new_n139));
  norb02aa1n02x5               g044(.a(new_n98), .b(new_n139), .out0(new_n140));
  norb02aa1n02x5               g045(.a(new_n128), .b(new_n139), .out0(new_n141));
  aboi22aa1n03x5               g046(.a(new_n140), .b(new_n138), .c(new_n137), .d(new_n141), .out0(new_n142));
  xorb03aa1n02x5               g047(.a(new_n142), .b(\b[10] ), .c(new_n132), .out0(\s[11] ));
  nor002aa1d32x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n144), .o1(new_n145));
  xorc02aa1n02x5               g050(.a(\a[11] ), .b(\b[10] ), .out0(new_n146));
  nanb02aa1n03x5               g051(.a(new_n142), .b(new_n146), .out0(new_n147));
  xorc02aa1n02x5               g052(.a(\a[12] ), .b(\b[11] ), .out0(new_n148));
  nand02aa1d24x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  inv020aa1n03x5               g054(.a(new_n149), .o1(new_n150));
  oai022aa1n02x5               g055(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n151));
  nona22aa1n02x4               g056(.a(new_n147), .b(new_n150), .c(new_n151), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n148), .c(new_n145), .d(new_n147), .o1(\s[12] ));
  nor002aa1d32x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  aoi012aa1d24x5               g059(.a(new_n154), .b(\a[11] ), .c(\b[10] ), .o1(new_n155));
  nona23aa1d18x5               g060(.a(new_n155), .b(new_n138), .c(new_n150), .d(new_n144), .out0(new_n156));
  nano22aa1n03x7               g061(.a(new_n156), .b(new_n128), .c(new_n130), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n127), .c(new_n122), .d(new_n107), .o1(new_n158));
  tech160nm_fioai012aa1n03p5x5 g063(.a(new_n149), .b(new_n154), .c(new_n144), .o1(new_n159));
  aoai13aa1n12x5               g064(.a(new_n159), .b(new_n156), .c(new_n98), .d(new_n130), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  xorc02aa1n12x5               g066(.a(\a[13] ), .b(\b[12] ), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n158), .c(new_n161), .out0(\s[13] ));
  inv000aa1d42x5               g068(.a(\a[13] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(\b[12] ), .b(new_n164), .out0(new_n165));
  aoai13aa1n03x5               g070(.a(new_n162), .b(new_n160), .c(new_n137), .d(new_n157), .o1(new_n166));
  xorc02aa1n12x5               g071(.a(\a[14] ), .b(\b[13] ), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n166), .c(new_n165), .out0(\s[14] ));
  nanp02aa1n03x5               g073(.a(new_n167), .b(new_n162), .o1(new_n169));
  inv040aa1d32x5               g074(.a(\a[14] ), .o1(new_n170));
  inv000aa1d42x5               g075(.a(\b[13] ), .o1(new_n171));
  nor002aa1n03x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  tech160nm_fioaoi03aa1n03p5x5 g077(.a(new_n170), .b(new_n171), .c(new_n172), .o1(new_n173));
  aoai13aa1n06x5               g078(.a(new_n173), .b(new_n169), .c(new_n158), .d(new_n161), .o1(new_n174));
  xorb03aa1n02x5               g079(.a(new_n174), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  xorc02aa1n12x5               g080(.a(\a[16] ), .b(\b[15] ), .out0(new_n176));
  nor002aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  xorc02aa1n12x5               g082(.a(\a[15] ), .b(\b[14] ), .out0(new_n178));
  aoi012aa1n02x5               g083(.a(new_n177), .b(new_n174), .c(new_n178), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n176), .b(new_n177), .out0(new_n180));
  aob012aa1n02x5               g085(.a(new_n180), .b(new_n174), .c(new_n178), .out0(new_n181));
  oaih12aa1n02x5               g086(.a(new_n181), .b(new_n179), .c(new_n176), .o1(\s[16] ));
  xroi22aa1d06x4               g087(.a(new_n164), .b(\b[12] ), .c(new_n170), .d(\b[13] ), .out0(new_n183));
  nand23aa1n03x5               g088(.a(new_n183), .b(new_n178), .c(new_n176), .o1(new_n184));
  nano22aa1n03x7               g089(.a(new_n169), .b(new_n178), .c(new_n176), .out0(new_n185));
  inv000aa1d42x5               g090(.a(\a[16] ), .o1(new_n186));
  inv020aa1n02x5               g091(.a(new_n177), .o1(new_n187));
  nanp02aa1n03x5               g092(.a(new_n173), .b(new_n187), .o1(new_n188));
  aoi022aa1n02x5               g093(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n188), .b(new_n189), .o1(new_n190));
  oaib12aa1n02x5               g095(.a(new_n190), .b(\b[15] ), .c(new_n186), .out0(new_n191));
  aoi012aa1d18x5               g096(.a(new_n191), .b(new_n160), .c(new_n185), .o1(new_n192));
  oaih12aa1n12x5               g097(.a(new_n192), .b(new_n158), .c(new_n184), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g099(.a(\a[17] ), .o1(new_n195));
  inv040aa1d28x5               g100(.a(\b[16] ), .o1(new_n196));
  nand42aa1n02x5               g101(.a(new_n196), .b(new_n195), .o1(new_n197));
  inv040aa1n03x5               g102(.a(new_n155), .o1(new_n198));
  nano32aa1n02x4               g103(.a(new_n198), .b(new_n145), .c(new_n149), .d(new_n138), .out0(new_n199));
  oaib12aa1n02x5               g104(.a(new_n199), .b(new_n139), .c(new_n98), .out0(new_n200));
  inv000aa1d42x5               g105(.a(\b[15] ), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n188), .b(new_n189), .c(new_n201), .d(new_n186), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n184), .c(new_n200), .d(new_n159), .o1(new_n203));
  aoi012aa1n06x5               g108(.a(new_n127), .b(new_n122), .c(new_n107), .o1(new_n204));
  nano22aa1n03x7               g109(.a(new_n204), .b(new_n157), .c(new_n185), .out0(new_n205));
  oai022aa1n02x5               g110(.a(new_n205), .b(new_n203), .c(new_n196), .d(new_n195), .o1(new_n206));
  nor042aa1n02x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nanp02aa1n04x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n206), .c(new_n197), .out0(\s[18] ));
  nanp02aa1n02x5               g115(.a(\b[16] ), .b(\a[17] ), .o1(new_n211));
  nano32aa1n03x7               g116(.a(new_n207), .b(new_n197), .c(new_n208), .d(new_n211), .out0(new_n212));
  tech160nm_fioaoi03aa1n03p5x5 g117(.a(\a[18] ), .b(\b[17] ), .c(new_n197), .o1(new_n213));
  nor002aa1d32x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand02aa1n06x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n213), .c(new_n193), .d(new_n212), .o1(new_n217));
  aoi112aa1n02x5               g122(.a(new_n216), .b(new_n213), .c(new_n193), .d(new_n212), .o1(new_n218));
  norb02aa1n03x4               g123(.a(new_n217), .b(new_n218), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n06x5               g125(.a(new_n214), .o1(new_n221));
  nor002aa1n12x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand22aa1n04x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  norb03aa1n02x5               g129(.a(new_n223), .b(new_n214), .c(new_n222), .out0(new_n225));
  nanp02aa1n03x5               g130(.a(new_n217), .b(new_n225), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n224), .c(new_n217), .d(new_n221), .o1(\s[20] ));
  nano23aa1n06x5               g132(.a(new_n214), .b(new_n222), .c(new_n223), .d(new_n215), .out0(new_n228));
  nanp02aa1n02x5               g133(.a(new_n212), .b(new_n228), .o1(new_n229));
  oabi12aa1n06x5               g134(.a(new_n229), .b(new_n205), .c(new_n203), .out0(new_n230));
  aoi013aa1n06x4               g135(.a(new_n207), .b(new_n208), .c(new_n195), .d(new_n196), .o1(new_n231));
  nona23aa1d18x5               g136(.a(new_n223), .b(new_n215), .c(new_n214), .d(new_n222), .out0(new_n232));
  tech160nm_fioaoi03aa1n03p5x5 g137(.a(\a[20] ), .b(\b[19] ), .c(new_n221), .o1(new_n233));
  oabi12aa1n18x5               g138(.a(new_n233), .b(new_n232), .c(new_n231), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  xnbna2aa1n03x5               g142(.a(new_n237), .b(new_n230), .c(new_n235), .out0(\s[21] ));
  inv000aa1n02x5               g143(.a(new_n157), .o1(new_n239));
  nona22aa1n02x4               g144(.a(new_n137), .b(new_n239), .c(new_n184), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n235), .b(new_n229), .c(new_n240), .d(new_n192), .o1(new_n241));
  nor042aa1n12x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  tech160nm_fixnrc02aa1n04x5   g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n242), .c(new_n241), .d(new_n237), .o1(new_n244));
  norp02aa1n02x5               g149(.a(new_n243), .b(new_n242), .o1(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n236), .c(new_n230), .d(new_n235), .o1(new_n246));
  nanp02aa1n03x5               g151(.a(new_n244), .b(new_n246), .o1(\s[22] ));
  nor042aa1n06x5               g152(.a(new_n243), .b(new_n236), .o1(new_n248));
  and003aa1n02x5               g153(.a(new_n248), .b(new_n212), .c(new_n228), .o(new_n249));
  oaih12aa1n02x5               g154(.a(new_n249), .b(new_n205), .c(new_n203), .o1(new_n250));
  inv020aa1d32x5               g155(.a(\a[22] ), .o1(new_n251));
  inv040aa1d32x5               g156(.a(\b[21] ), .o1(new_n252));
  oao003aa1n12x5               g157(.a(new_n251), .b(new_n252), .c(new_n242), .carry(new_n253));
  aoi012aa1n09x5               g158(.a(new_n253), .b(new_n234), .c(new_n248), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[22] ), .b(\a[23] ), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  xnbna2aa1n03x5               g161(.a(new_n256), .b(new_n250), .c(new_n254), .out0(\s[23] ));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n254), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n256), .b(new_n260), .c(new_n193), .d(new_n249), .o1(new_n261));
  tech160nm_fixorc02aa1n02p5x5 g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  nanp02aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .o1(new_n263));
  oai022aa1n02x5               g168(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n263), .b(new_n264), .out0(new_n265));
  aoai13aa1n02x5               g170(.a(new_n265), .b(new_n255), .c(new_n250), .d(new_n254), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n266), .b(new_n262), .c(new_n261), .d(new_n259), .o1(\s[24] ));
  nano32aa1n02x5               g172(.a(new_n229), .b(new_n262), .c(new_n248), .d(new_n256), .out0(new_n268));
  oai012aa1n02x5               g173(.a(new_n268), .b(new_n205), .c(new_n203), .o1(new_n269));
  aoai13aa1n06x5               g174(.a(new_n248), .b(new_n233), .c(new_n228), .d(new_n213), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n253), .o1(new_n271));
  norb02aa1n06x5               g176(.a(new_n262), .b(new_n255), .out0(new_n272));
  inv000aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  nanp02aa1n02x5               g178(.a(new_n264), .b(new_n263), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n270), .d(new_n271), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n269), .c(new_n276), .out0(\s[25] ));
  norp02aa1n02x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n277), .b(new_n275), .c(new_n193), .d(new_n268), .o1(new_n281));
  xorc02aa1n03x5               g186(.a(\a[26] ), .b(\b[25] ), .out0(new_n282));
  nanp02aa1n02x5               g187(.a(\b[25] ), .b(\a[26] ), .o1(new_n283));
  oai022aa1n02x5               g188(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n284));
  norb02aa1n02x5               g189(.a(new_n283), .b(new_n284), .out0(new_n285));
  nand42aa1n02x5               g190(.a(new_n281), .b(new_n285), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n282), .c(new_n281), .d(new_n280), .o1(\s[26] ));
  nor042aa1n03x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  and002aa1n24x5               g193(.a(\b[26] ), .b(\a[27] ), .o(new_n289));
  nor042aa1n03x5               g194(.a(new_n289), .b(new_n288), .o1(new_n290));
  and002aa1n09x5               g195(.a(new_n282), .b(new_n277), .o(new_n291));
  nano32aa1n03x7               g196(.a(new_n229), .b(new_n291), .c(new_n248), .d(new_n272), .out0(new_n292));
  tech160nm_fioai012aa1n05x5   g197(.a(new_n292), .b(new_n205), .c(new_n203), .o1(new_n293));
  aoi022aa1n06x5               g198(.a(new_n275), .b(new_n291), .c(new_n283), .d(new_n284), .o1(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n290), .b(new_n294), .c(new_n293), .out0(\s[27] ));
  inv000aa1d42x5               g200(.a(new_n289), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n272), .b(new_n253), .c(new_n234), .d(new_n248), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n291), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n284), .b(new_n283), .o1(new_n299));
  aoai13aa1n04x5               g204(.a(new_n299), .b(new_n298), .c(new_n297), .d(new_n274), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n296), .b(new_n300), .c(new_n193), .d(new_n292), .o1(new_n301));
  inv000aa1n03x5               g206(.a(new_n288), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n289), .c(new_n294), .d(new_n293), .o1(new_n303));
  xorc02aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .out0(new_n304));
  norp02aa1n02x5               g209(.a(new_n304), .b(new_n288), .o1(new_n305));
  aoi022aa1n03x5               g210(.a(new_n303), .b(new_n304), .c(new_n301), .d(new_n305), .o1(\s[28] ));
  and002aa1n03x5               g211(.a(new_n304), .b(new_n290), .o(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n300), .c(new_n193), .d(new_n292), .o1(new_n308));
  inv000aa1n02x5               g213(.a(new_n307), .o1(new_n309));
  oao003aa1n03x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n302), .carry(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n309), .c(new_n294), .d(new_n293), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n308), .d(new_n313), .o1(\s[29] ));
  nanp02aa1n02x5               g219(.a(\b[0] ), .b(\a[1] ), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g221(.a(new_n304), .b(new_n312), .c(new_n290), .o(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n300), .c(new_n193), .d(new_n292), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  oaoi03aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .o1(new_n320));
  inv000aa1n03x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n319), .c(new_n294), .d(new_n293), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(\b[28] ), .b(\a[29] ), .o(new_n324));
  oabi12aa1n02x5               g229(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n325));
  oab012aa1n02x4               g230(.a(new_n325), .b(new_n310), .c(new_n324), .out0(new_n326));
  aoi022aa1n03x5               g231(.a(new_n322), .b(new_n323), .c(new_n318), .d(new_n326), .o1(\s[30] ));
  nano22aa1n03x7               g232(.a(new_n309), .b(new_n312), .c(new_n323), .out0(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n300), .c(new_n193), .d(new_n292), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  oao003aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n331));
  norb02aa1n02x5               g236(.a(new_n331), .b(new_n330), .out0(new_n332));
  inv000aa1d42x5               g237(.a(new_n328), .o1(new_n333));
  aoai13aa1n02x7               g238(.a(new_n331), .b(new_n333), .c(new_n294), .d(new_n293), .o1(new_n334));
  aoi022aa1n03x5               g239(.a(new_n334), .b(new_n330), .c(new_n329), .d(new_n332), .o1(\s[31] ));
  xnbna2aa1n03x5               g240(.a(new_n103), .b(new_n105), .c(new_n104), .out0(\s[3] ));
  norb02aa1n02x5               g241(.a(new_n108), .b(new_n100), .out0(new_n337));
  aoi113aa1n02x5               g242(.a(new_n99), .b(new_n337), .c(new_n105), .d(new_n104), .e(new_n102), .o1(new_n338));
  aoi012aa1n02x5               g243(.a(new_n338), .b(new_n107), .c(new_n337), .o1(\s[4] ));
  nanb02aa1n02x5               g244(.a(new_n110), .b(new_n109), .out0(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n340), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  aoai13aa1n02x5               g246(.a(new_n109), .b(new_n110), .c(new_n107), .d(new_n108), .o1(new_n342));
  xnrb03aa1n02x5               g247(.a(new_n342), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n03x5               g248(.a(\a[6] ), .b(\b[5] ), .c(new_n342), .o1(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g250(.a(new_n117), .b(new_n118), .c(new_n344), .o1(new_n346));
  xorb03aa1n02x5               g251(.a(new_n346), .b(\b[7] ), .c(new_n113), .out0(\s[8] ));
  xorb03aa1n02x5               g252(.a(new_n204), .b(\b[8] ), .c(new_n97), .out0(\s[9] ));
endmodule


