// Benchmark "adder" written by ABC on Thu Jul 18 01:35:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n180, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n337, new_n340,
    new_n342, new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(new_n101), .o1(new_n102));
  nor042aa1n04x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nor042aa1n03x5               g008(.a(\b[4] ), .b(\a[5] ), .o1(new_n104));
  nor022aa1n02x5               g009(.a(new_n104), .b(new_n103), .o1(new_n105));
  nand42aa1n08x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  inv000aa1n02x5               g011(.a(new_n106), .o1(new_n107));
  nor002aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand42aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  norb02aa1n03x4               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  nor022aa1n06x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  norb02aa1n03x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nona23aa1n06x5               g018(.a(new_n113), .b(new_n110), .c(new_n105), .d(new_n107), .out0(new_n114));
  tech160nm_fioai012aa1n03p5x5 g019(.a(new_n109), .b(new_n111), .c(new_n108), .o1(new_n115));
  nand22aa1n03x5               g020(.a(new_n114), .b(new_n115), .o1(new_n116));
  nor002aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  nand42aa1n06x5               g022(.a(\b[0] ), .b(\a[1] ), .o1(new_n118));
  nand22aa1n02x5               g023(.a(\b[1] ), .b(\a[2] ), .o1(new_n119));
  tech160nm_fiaoi012aa1n05x5   g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  norp02aa1n06x5               g025(.a(\b[3] ), .b(\a[4] ), .o1(new_n121));
  tech160nm_finand02aa1n03p5x5 g026(.a(\b[3] ), .b(\a[4] ), .o1(new_n122));
  nor042aa1n04x5               g027(.a(\b[2] ), .b(\a[3] ), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(\b[2] ), .b(\a[3] ), .o1(new_n124));
  nona23aa1n09x5               g029(.a(new_n124), .b(new_n122), .c(new_n121), .d(new_n123), .out0(new_n125));
  inv000aa1d42x5               g030(.a(\a[3] ), .o1(new_n126));
  inv000aa1d42x5               g031(.a(\b[2] ), .o1(new_n127));
  aoai13aa1n04x5               g032(.a(new_n122), .b(new_n121), .c(new_n126), .d(new_n127), .o1(new_n128));
  oai012aa1n12x5               g033(.a(new_n128), .b(new_n125), .c(new_n120), .o1(new_n129));
  nona23aa1n06x5               g034(.a(new_n112), .b(new_n109), .c(new_n108), .d(new_n111), .out0(new_n130));
  norb02aa1n02x5               g035(.a(new_n106), .b(new_n103), .out0(new_n131));
  nand42aa1n02x5               g036(.a(\b[4] ), .b(\a[5] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n104), .out0(new_n133));
  nano22aa1n09x5               g038(.a(new_n130), .b(new_n131), .c(new_n133), .out0(new_n134));
  nand42aa1n08x5               g039(.a(\b[8] ), .b(\a[9] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n101), .out0(new_n136));
  aoai13aa1n06x5               g041(.a(new_n136), .b(new_n116), .c(new_n129), .d(new_n134), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n100), .b(new_n137), .c(new_n102), .out0(\s[10] ));
  oai012aa1d24x5               g043(.a(new_n98), .b(new_n101), .c(new_n97), .o1(new_n139));
  inv040aa1d32x5               g044(.a(\a[11] ), .o1(new_n140));
  inv040aa1d28x5               g045(.a(\b[10] ), .o1(new_n141));
  nand02aa1d16x5               g046(.a(new_n141), .b(new_n140), .o1(new_n142));
  nand42aa1n02x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nand02aa1n03x5               g048(.a(new_n142), .b(new_n143), .o1(new_n144));
  oaoi13aa1n04x5               g049(.a(new_n144), .b(new_n139), .c(new_n137), .d(new_n99), .o1(new_n145));
  oai112aa1n02x5               g050(.a(new_n139), .b(new_n144), .c(new_n137), .d(new_n99), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(\s[11] ));
  inv040aa1d32x5               g052(.a(\a[12] ), .o1(new_n148));
  inv030aa1d32x5               g053(.a(\b[11] ), .o1(new_n149));
  nand02aa1d28x5               g054(.a(new_n149), .b(new_n148), .o1(new_n150));
  nand02aa1n06x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nand22aa1n12x5               g056(.a(new_n150), .b(new_n151), .o1(new_n152));
  nano22aa1n02x4               g057(.a(new_n145), .b(new_n142), .c(new_n152), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n152), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n145), .c(new_n140), .d(new_n141), .o1(new_n155));
  norb02aa1n02x7               g060(.a(new_n155), .b(new_n153), .out0(\s[12] ));
  nano23aa1n06x5               g061(.a(new_n97), .b(new_n101), .c(new_n135), .d(new_n98), .out0(new_n157));
  nona22aa1d18x5               g062(.a(new_n157), .b(new_n152), .c(new_n144), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n159), .b(new_n116), .c(new_n129), .d(new_n134), .o1(new_n160));
  aoi022aa1n09x5               g065(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n161));
  inv000aa1n02x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n12x5               g067(.a(new_n150), .b(new_n162), .c(new_n139), .d(new_n142), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  nor002aa1d32x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand42aa1d28x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n160), .c(new_n164), .out0(\s[13] ));
  inv000aa1d42x5               g073(.a(new_n165), .o1(new_n169));
  oai022aa1n02x5               g074(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n170));
  nano22aa1n02x4               g075(.a(new_n130), .b(new_n170), .c(new_n106), .out0(new_n171));
  norb02aa1n02x5               g076(.a(new_n115), .b(new_n171), .out0(new_n172));
  nanp02aa1n02x5               g077(.a(new_n129), .b(new_n134), .o1(new_n173));
  nanp02aa1n06x5               g078(.a(new_n173), .b(new_n172), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n167), .b(new_n163), .c(new_n174), .d(new_n159), .o1(new_n175));
  nor022aa1n06x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  nand42aa1n16x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  xnbna2aa1n03x5               g083(.a(new_n178), .b(new_n175), .c(new_n169), .out0(\s[14] ));
  nano23aa1d15x5               g084(.a(new_n165), .b(new_n176), .c(new_n177), .d(new_n166), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  oai012aa1n03x5               g086(.a(new_n177), .b(new_n176), .c(new_n165), .o1(new_n182));
  aoai13aa1n04x5               g087(.a(new_n182), .b(new_n181), .c(new_n160), .d(new_n164), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv040aa1d32x5               g089(.a(\a[15] ), .o1(new_n185));
  inv000aa1d48x5               g090(.a(\b[14] ), .o1(new_n186));
  nand02aa1d08x5               g091(.a(new_n186), .b(new_n185), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(\b[14] ), .b(\a[15] ), .o1(new_n189));
  inv040aa1d32x5               g094(.a(\a[16] ), .o1(new_n190));
  inv040aa1d28x5               g095(.a(\b[15] ), .o1(new_n191));
  nand22aa1n09x5               g096(.a(new_n191), .b(new_n190), .o1(new_n192));
  nand22aa1n03x5               g097(.a(\b[15] ), .b(\a[16] ), .o1(new_n193));
  nand22aa1n06x5               g098(.a(new_n192), .b(new_n193), .o1(new_n194));
  inv000aa1d42x5               g099(.a(new_n194), .o1(new_n195));
  aoi112aa1n02x5               g100(.a(new_n188), .b(new_n195), .c(new_n183), .d(new_n189), .o1(new_n196));
  aoai13aa1n04x5               g101(.a(new_n195), .b(new_n188), .c(new_n183), .d(new_n189), .o1(new_n197));
  norb02aa1n02x7               g102(.a(new_n197), .b(new_n196), .out0(\s[16] ));
  xnrc02aa1n12x5               g103(.a(\b[16] ), .b(\a[17] ), .out0(new_n199));
  nand42aa1n02x5               g104(.a(new_n187), .b(new_n189), .o1(new_n200));
  nona22aa1d24x5               g105(.a(new_n180), .b(new_n200), .c(new_n194), .out0(new_n201));
  nor042aa1n09x5               g106(.a(new_n201), .b(new_n158), .o1(new_n202));
  aoai13aa1n12x5               g107(.a(new_n202), .b(new_n116), .c(new_n129), .d(new_n134), .o1(new_n203));
  nand42aa1n02x5               g108(.a(new_n182), .b(new_n187), .o1(new_n204));
  aoi022aa1n02x5               g109(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n205));
  aob012aa1n02x5               g110(.a(new_n192), .b(new_n204), .c(new_n205), .out0(new_n206));
  aoib12aa1n12x5               g111(.a(new_n206), .b(new_n163), .c(new_n201), .out0(new_n207));
  xobna2aa1n03x5               g112(.a(new_n199), .b(new_n203), .c(new_n207), .out0(\s[17] ));
  inv000aa1d42x5               g113(.a(\a[18] ), .o1(new_n209));
  norp02aa1n02x5               g114(.a(\b[16] ), .b(\a[17] ), .o1(new_n210));
  nanp02aa1n06x5               g115(.a(new_n203), .b(new_n207), .o1(new_n211));
  aoib12aa1n02x5               g116(.a(new_n210), .b(new_n211), .c(new_n199), .out0(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[17] ), .c(new_n209), .out0(\s[18] ));
  xnrc02aa1n02x5               g118(.a(\b[17] ), .b(\a[18] ), .out0(new_n214));
  nor042aa1n04x5               g119(.a(new_n214), .b(new_n199), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  nand42aa1n02x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  oai022aa1d24x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  and002aa1n02x5               g123(.a(new_n218), .b(new_n217), .o(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n216), .c(new_n203), .d(new_n207), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g127(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n02x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  nand42aa1n03x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  norp02aa1n04x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  tech160nm_finand02aa1n03p5x5 g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n227), .b(new_n226), .out0(new_n228));
  aoi112aa1n02x5               g133(.a(new_n224), .b(new_n228), .c(new_n221), .d(new_n225), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n228), .b(new_n224), .c(new_n221), .d(new_n225), .o1(new_n230));
  norb02aa1n02x7               g135(.a(new_n230), .b(new_n229), .out0(\s[20] ));
  nanb03aa1n09x5               g136(.a(new_n226), .b(new_n227), .c(new_n225), .out0(new_n232));
  nona22aa1n02x4               g137(.a(new_n215), .b(new_n224), .c(new_n232), .out0(new_n233));
  oai112aa1n06x5               g138(.a(new_n218), .b(new_n217), .c(\b[18] ), .d(\a[19] ), .o1(new_n234));
  tech160nm_fioai012aa1n04x5   g139(.a(new_n227), .b(new_n226), .c(new_n224), .o1(new_n235));
  oai012aa1n18x5               g140(.a(new_n235), .b(new_n234), .c(new_n232), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n233), .c(new_n203), .d(new_n207), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  xnrc02aa1n12x5               g145(.a(\b[20] ), .b(\a[21] ), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoi112aa1n03x5               g149(.a(new_n240), .b(new_n244), .c(new_n238), .d(new_n242), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n244), .b(new_n240), .c(new_n238), .d(new_n242), .o1(new_n246));
  norb02aa1n02x7               g151(.a(new_n246), .b(new_n245), .out0(\s[22] ));
  nor042aa1n06x5               g152(.a(new_n243), .b(new_n241), .o1(new_n248));
  nona23aa1n06x5               g153(.a(new_n215), .b(new_n248), .c(new_n232), .d(new_n224), .out0(new_n249));
  inv000aa1d42x5               g154(.a(\a[22] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[21] ), .o1(new_n251));
  oao003aa1n02x5               g156(.a(new_n250), .b(new_n251), .c(new_n240), .carry(new_n252));
  aoi012aa1n02x5               g157(.a(new_n252), .b(new_n236), .c(new_n248), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n249), .c(new_n203), .d(new_n207), .o1(new_n254));
  xorb03aa1n02x5               g159(.a(new_n254), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  tech160nm_fixorc02aa1n05x5   g161(.a(\a[23] ), .b(\b[22] ), .out0(new_n257));
  xorc02aa1n12x5               g162(.a(\a[24] ), .b(\b[23] ), .out0(new_n258));
  aoi112aa1n02x5               g163(.a(new_n256), .b(new_n258), .c(new_n254), .d(new_n257), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n258), .b(new_n256), .c(new_n254), .d(new_n257), .o1(new_n260));
  norb02aa1n03x4               g165(.a(new_n260), .b(new_n259), .out0(\s[24] ));
  nano22aa1n02x4               g166(.a(new_n226), .b(new_n225), .c(new_n227), .out0(new_n262));
  oai012aa1n02x5               g167(.a(new_n217), .b(\b[18] ), .c(\a[19] ), .o1(new_n263));
  norb02aa1n02x5               g168(.a(new_n218), .b(new_n263), .out0(new_n264));
  inv000aa1n06x5               g169(.a(new_n235), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n248), .b(new_n265), .c(new_n264), .d(new_n262), .o1(new_n266));
  inv020aa1n02x5               g171(.a(new_n252), .o1(new_n267));
  and002aa1n02x5               g172(.a(new_n258), .b(new_n257), .o(new_n268));
  inv000aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  oai022aa1n02x5               g174(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n270));
  aob012aa1n02x5               g175(.a(new_n270), .b(\b[23] ), .c(\a[24] ), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n269), .c(new_n266), .d(new_n267), .o1(new_n272));
  nano32aa1n02x4               g177(.a(new_n233), .b(new_n258), .c(new_n248), .d(new_n257), .out0(new_n273));
  tech160nm_fixorc02aa1n04x5   g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n272), .c(new_n211), .d(new_n273), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(new_n272), .b(new_n274), .c(new_n211), .d(new_n273), .o1(new_n276));
  norb02aa1n02x5               g181(.a(new_n275), .b(new_n276), .out0(\s[25] ));
  nor042aa1n03x5               g182(.a(\b[24] ), .b(\a[25] ), .o1(new_n278));
  tech160nm_fixorc02aa1n02p5x5 g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  nona22aa1n02x5               g184(.a(new_n275), .b(new_n279), .c(new_n278), .out0(new_n280));
  inv000aa1d42x5               g185(.a(new_n278), .o1(new_n281));
  aobi12aa1n06x5               g186(.a(new_n279), .b(new_n275), .c(new_n281), .out0(new_n282));
  norb02aa1n03x4               g187(.a(new_n280), .b(new_n282), .out0(\s[26] ));
  aoi022aa1n02x5               g188(.a(new_n204), .b(new_n205), .c(new_n191), .d(new_n190), .o1(new_n284));
  oaib12aa1n03x5               g189(.a(new_n284), .b(new_n201), .c(new_n163), .out0(new_n285));
  and002aa1n06x5               g190(.a(new_n279), .b(new_n274), .o(new_n286));
  nano22aa1n03x7               g191(.a(new_n249), .b(new_n268), .c(new_n286), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n287), .b(new_n285), .c(new_n174), .d(new_n202), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[26] ), .b(\b[25] ), .c(new_n281), .carry(new_n289));
  aobi12aa1n06x5               g194(.a(new_n289), .b(new_n272), .c(new_n286), .out0(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnbna2aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n288), .out0(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  inv040aa1n03x5               g198(.a(new_n293), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n291), .o1(new_n295));
  aoi012aa1n02x7               g200(.a(new_n295), .b(new_n290), .c(new_n288), .o1(new_n296));
  xnrc02aa1n12x5               g201(.a(\b[27] ), .b(\a[28] ), .out0(new_n297));
  nano22aa1n03x7               g202(.a(new_n296), .b(new_n294), .c(new_n297), .out0(new_n298));
  inv000aa1n02x5               g203(.a(new_n287), .o1(new_n299));
  aoi012aa1n06x5               g204(.a(new_n299), .b(new_n203), .c(new_n207), .o1(new_n300));
  aoai13aa1n12x5               g205(.a(new_n268), .b(new_n252), .c(new_n236), .d(new_n248), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n286), .o1(new_n302));
  aoai13aa1n06x5               g207(.a(new_n289), .b(new_n302), .c(new_n301), .d(new_n271), .o1(new_n303));
  oaih12aa1n02x5               g208(.a(new_n291), .b(new_n303), .c(new_n300), .o1(new_n304));
  aoi012aa1n03x5               g209(.a(new_n297), .b(new_n304), .c(new_n294), .o1(new_n305));
  norp02aa1n03x5               g210(.a(new_n305), .b(new_n298), .o1(\s[28] ));
  xnrc02aa1n02x5               g211(.a(\b[28] ), .b(\a[29] ), .out0(new_n307));
  norb02aa1d21x5               g212(.a(new_n291), .b(new_n297), .out0(new_n308));
  tech160nm_fioai012aa1n03p5x5 g213(.a(new_n308), .b(new_n303), .c(new_n300), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n294), .carry(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n307), .b(new_n309), .c(new_n310), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n308), .o1(new_n312));
  tech160nm_fiaoi012aa1n05x5   g217(.a(new_n312), .b(new_n290), .c(new_n288), .o1(new_n313));
  nano22aa1n03x7               g218(.a(new_n313), .b(new_n307), .c(new_n310), .out0(new_n314));
  norp02aa1n03x5               g219(.a(new_n311), .b(new_n314), .o1(\s[29] ));
  xorb03aa1n02x5               g220(.a(new_n118), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g221(.a(\b[29] ), .b(\a[30] ), .out0(new_n317));
  norb03aa1n12x5               g222(.a(new_n291), .b(new_n307), .c(new_n297), .out0(new_n318));
  oaih12aa1n02x5               g223(.a(new_n318), .b(new_n303), .c(new_n300), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .carry(new_n320));
  aoi012aa1n03x5               g225(.a(new_n317), .b(new_n319), .c(new_n320), .o1(new_n321));
  inv000aa1d42x5               g226(.a(new_n318), .o1(new_n322));
  tech160nm_fiaoi012aa1n05x5   g227(.a(new_n322), .b(new_n290), .c(new_n288), .o1(new_n323));
  nano22aa1n03x7               g228(.a(new_n323), .b(new_n317), .c(new_n320), .out0(new_n324));
  nor002aa1n02x5               g229(.a(new_n321), .b(new_n324), .o1(\s[30] ));
  xnrc02aa1n02x5               g230(.a(\b[30] ), .b(\a[31] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n318), .b(new_n317), .out0(new_n327));
  oaih12aa1n02x5               g232(.a(new_n327), .b(new_n303), .c(new_n300), .o1(new_n328));
  oao003aa1n02x5               g233(.a(\a[30] ), .b(\b[29] ), .c(new_n320), .carry(new_n329));
  aoi012aa1n03x5               g234(.a(new_n326), .b(new_n328), .c(new_n329), .o1(new_n330));
  inv000aa1n02x5               g235(.a(new_n327), .o1(new_n331));
  tech160nm_fiaoi012aa1n05x5   g236(.a(new_n331), .b(new_n290), .c(new_n288), .o1(new_n332));
  nano22aa1n03x7               g237(.a(new_n332), .b(new_n326), .c(new_n329), .out0(new_n333));
  norp02aa1n03x5               g238(.a(new_n330), .b(new_n333), .o1(\s[31] ));
  xorb03aa1n02x5               g239(.a(new_n120), .b(\b[2] ), .c(new_n126), .out0(\s[3] ));
  nona22aa1n02x4               g240(.a(new_n124), .b(new_n120), .c(new_n123), .out0(new_n336));
  aboi22aa1n03x5               g241(.a(new_n121), .b(new_n122), .c(new_n126), .d(new_n127), .out0(new_n337));
  aboi22aa1n03x5               g242(.a(new_n121), .b(new_n129), .c(new_n336), .d(new_n337), .out0(\s[4] ));
  xorb03aa1n02x5               g243(.a(new_n129), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fiao0012aa1n02p5x5 g244(.a(new_n104), .b(new_n129), .c(new_n132), .o(new_n340));
  xorb03aa1n02x5               g245(.a(new_n340), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi012aa1n06x5               g246(.a(new_n103), .b(new_n340), .c(new_n106), .o1(new_n342));
  xnrc02aa1n02x5               g247(.a(new_n342), .b(new_n113), .out0(\s[7] ));
  oaoi03aa1n02x5               g248(.a(\a[7] ), .b(\b[6] ), .c(new_n342), .o1(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g250(.a(new_n136), .b(new_n173), .c(new_n172), .out0(\s[9] ));
endmodule


