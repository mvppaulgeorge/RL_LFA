// Benchmark "adder" written by ABC on Thu Jul 18 00:21:43 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n325, new_n326,
    new_n328, new_n330, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[4] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[3] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(new_n99), .b(new_n100), .o1(new_n101));
  nor002aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanb02aa1n03x5               g008(.a(new_n102), .b(new_n103), .out0(new_n104));
  nanp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand22aa1n03x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  tech160nm_fioai012aa1n04x5   g012(.a(new_n105), .b(new_n107), .c(new_n106), .o1(new_n108));
  oaoi03aa1n09x5               g013(.a(new_n97), .b(new_n98), .c(new_n102), .o1(new_n109));
  oai013aa1n06x5               g014(.a(new_n109), .b(new_n104), .c(new_n108), .d(new_n101), .o1(new_n110));
  nor042aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand02aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  norp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nor043aa1n03x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  aoi112aa1n06x5               g023(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n119));
  nano23aa1n02x4               g024(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n120));
  and002aa1n06x5               g025(.a(\b[5] ), .b(\a[6] ), .o(new_n121));
  oai022aa1d24x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n122), .o1(new_n123));
  nona22aa1n02x4               g028(.a(new_n120), .b(new_n121), .c(new_n123), .out0(new_n124));
  nona22aa1n02x4               g029(.a(new_n124), .b(new_n119), .c(new_n111), .out0(new_n125));
  aoi012aa1n02x5               g030(.a(new_n125), .b(new_n110), .c(new_n118), .o1(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[9] ), .b(\b[8] ), .c(new_n126), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor043aa1n02x5               g033(.a(new_n108), .b(new_n104), .c(new_n101), .o1(new_n129));
  inv000aa1d42x5               g034(.a(new_n109), .o1(new_n130));
  tech160nm_fioai012aa1n05x5   g035(.a(new_n118), .b(new_n129), .c(new_n130), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n111), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n119), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n121), .o1(new_n134));
  nano22aa1n03x5               g039(.a(new_n115), .b(new_n134), .c(new_n122), .out0(new_n135));
  nano22aa1n09x5               g040(.a(new_n135), .b(new_n132), .c(new_n133), .out0(new_n136));
  nor002aa1n02x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nand22aa1n03x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  norp02aa1n04x5               g043(.a(\b[8] ), .b(\a[9] ), .o1(new_n139));
  nand42aa1n02x5               g044(.a(\b[8] ), .b(\a[9] ), .o1(new_n140));
  nona23aa1d18x5               g045(.a(new_n140), .b(new_n138), .c(new_n137), .d(new_n139), .out0(new_n141));
  oai012aa1n02x5               g046(.a(new_n138), .b(new_n139), .c(new_n137), .o1(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n141), .c(new_n131), .d(new_n136), .o1(new_n143));
  xorb03aa1n02x5               g048(.a(new_n143), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n02x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  nanp02aa1n02x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  aoi012aa1n02x5               g051(.a(new_n145), .b(new_n143), .c(new_n146), .o1(new_n147));
  xnrb03aa1n02x5               g052(.a(new_n147), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n02x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nona23aa1n02x4               g055(.a(new_n150), .b(new_n146), .c(new_n145), .d(new_n149), .out0(new_n151));
  aoi112aa1n03x5               g056(.a(new_n151), .b(new_n141), .c(new_n131), .d(new_n136), .o1(new_n152));
  tech160nm_fiao0012aa1n02p5x5 g057(.a(new_n149), .b(new_n145), .c(new_n150), .o(new_n153));
  oabi12aa1n03x5               g058(.a(new_n153), .b(new_n151), .c(new_n142), .out0(new_n154));
  nor042aa1n06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  oai112aa1n03x5               g062(.a(new_n156), .b(new_n157), .c(new_n152), .d(new_n154), .o1(new_n158));
  aoi112aa1n02x5               g063(.a(new_n152), .b(new_n154), .c(new_n157), .d(new_n156), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(\s[13] ));
  nor042aa1n02x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n158), .c(new_n156), .out0(\s[14] ));
  nor022aa1n08x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  nano23aa1n06x5               g072(.a(new_n155), .b(new_n161), .c(new_n162), .d(new_n157), .out0(new_n168));
  aoi012aa1n09x5               g073(.a(new_n161), .b(new_n155), .c(new_n162), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n170), .b(new_n154), .c(new_n168), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n141), .o1(new_n172));
  nano23aa1n06x5               g077(.a(new_n145), .b(new_n149), .c(new_n150), .d(new_n146), .out0(new_n173));
  nano32aa1n02x4               g078(.a(new_n126), .b(new_n168), .c(new_n172), .d(new_n173), .out0(new_n174));
  oaib12aa1n06x5               g079(.a(new_n167), .b(new_n174), .c(new_n171), .out0(new_n175));
  norb03aa1n02x5               g080(.a(new_n171), .b(new_n174), .c(new_n167), .out0(new_n176));
  norb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(\s[15] ));
  inv000aa1d42x5               g082(.a(new_n165), .o1(new_n178));
  norp02aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n175), .c(new_n178), .out0(\s[16] ));
  inv040aa1d32x5               g087(.a(\a[17] ), .o1(new_n183));
  and002aa1n02x5               g088(.a(\b[9] ), .b(\a[10] ), .o(new_n184));
  oab012aa1n09x5               g089(.a(new_n184), .b(new_n137), .c(new_n139), .out0(new_n185));
  aoai13aa1n09x5               g090(.a(new_n168), .b(new_n153), .c(new_n173), .d(new_n185), .o1(new_n186));
  nona23aa1n03x5               g091(.a(new_n180), .b(new_n166), .c(new_n165), .d(new_n179), .out0(new_n187));
  aoi012aa1n02x5               g092(.a(new_n179), .b(new_n165), .c(new_n180), .o1(new_n188));
  aoai13aa1n12x5               g093(.a(new_n188), .b(new_n187), .c(new_n186), .d(new_n169), .o1(new_n189));
  nona23aa1n09x5               g094(.a(new_n168), .b(new_n173), .c(new_n187), .d(new_n141), .out0(new_n190));
  aoi012aa1n12x5               g095(.a(new_n190), .b(new_n131), .c(new_n136), .o1(new_n191));
  nor042aa1n03x5               g096(.a(new_n189), .b(new_n191), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[16] ), .c(new_n183), .out0(\s[17] ));
  inv040aa1d32x5               g098(.a(\b[16] ), .o1(new_n194));
  nand42aa1n02x5               g099(.a(new_n194), .b(new_n183), .o1(new_n195));
  nor002aa1d32x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nand42aa1d28x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  and002aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o(new_n199));
  oabi12aa1n02x5               g104(.a(new_n199), .b(new_n189), .c(new_n191), .out0(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n198), .b(new_n200), .c(new_n195), .out0(\s[18] ));
  nano23aa1n03x7               g106(.a(new_n196), .b(new_n199), .c(new_n195), .d(new_n197), .out0(new_n202));
  oaih12aa1n02x5               g107(.a(new_n202), .b(new_n189), .c(new_n191), .o1(new_n203));
  aoai13aa1n12x5               g108(.a(new_n197), .b(new_n196), .c(new_n183), .d(new_n194), .o1(new_n204));
  nor042aa1n09x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanp02aa1n03x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  xobna2aa1n03x5               g112(.a(new_n207), .b(new_n203), .c(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g114(.a(new_n205), .o1(new_n210));
  aoi012aa1n02x5               g115(.a(new_n207), .b(new_n203), .c(new_n204), .o1(new_n211));
  nor042aa1n09x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand22aa1n02x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanb02aa1n02x5               g118(.a(new_n212), .b(new_n213), .out0(new_n214));
  nano22aa1n03x5               g119(.a(new_n211), .b(new_n210), .c(new_n214), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n204), .o1(new_n216));
  oaoi13aa1n02x5               g121(.a(new_n216), .b(new_n202), .c(new_n189), .d(new_n191), .o1(new_n217));
  oaoi13aa1n02x5               g122(.a(new_n214), .b(new_n210), .c(new_n217), .d(new_n207), .o1(new_n218));
  norp02aa1n02x5               g123(.a(new_n218), .b(new_n215), .o1(\s[20] ));
  inv000aa1d42x5               g124(.a(\a[21] ), .o1(new_n220));
  nona23aa1d18x5               g125(.a(new_n213), .b(new_n206), .c(new_n205), .d(new_n212), .out0(new_n221));
  nano23aa1n09x5               g126(.a(new_n221), .b(new_n199), .c(new_n195), .d(new_n198), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n212), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(new_n205), .b(new_n213), .o1(new_n224));
  oai112aa1n06x5               g129(.a(new_n224), .b(new_n223), .c(new_n221), .d(new_n204), .o1(new_n225));
  oaoi13aa1n06x5               g130(.a(new_n225), .b(new_n222), .c(new_n189), .d(new_n191), .o1(new_n226));
  xorb03aa1n02x5               g131(.a(new_n226), .b(\b[20] ), .c(new_n220), .out0(\s[21] ));
  nanb02aa1n02x5               g132(.a(\b[20] ), .b(new_n220), .out0(new_n228));
  inv000aa1n02x5               g133(.a(new_n222), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n225), .o1(new_n230));
  xnrc02aa1n03x5               g135(.a(\b[20] ), .b(\a[21] ), .out0(new_n231));
  oaoi13aa1n06x5               g136(.a(new_n231), .b(new_n230), .c(new_n192), .d(new_n229), .o1(new_n232));
  xnrc02aa1n02x5               g137(.a(\b[21] ), .b(\a[22] ), .out0(new_n233));
  nano22aa1n03x5               g138(.a(new_n232), .b(new_n228), .c(new_n233), .out0(new_n234));
  oaoi13aa1n02x7               g139(.a(new_n233), .b(new_n228), .c(new_n226), .d(new_n231), .o1(new_n235));
  norp02aa1n02x5               g140(.a(new_n235), .b(new_n234), .o1(\s[22] ));
  nor042aa1n03x5               g141(.a(new_n233), .b(new_n231), .o1(new_n237));
  oaoi03aa1n02x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n228), .o1(new_n238));
  ao0012aa1n03x7               g143(.a(new_n238), .b(new_n225), .c(new_n237), .o(new_n239));
  nanb03aa1n09x5               g144(.a(new_n221), .b(new_n237), .c(new_n202), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  oaoi13aa1n06x5               g146(.a(new_n239), .b(new_n241), .c(new_n189), .d(new_n191), .o1(new_n242));
  xnrb03aa1n03x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  oaih12aa1n02x5               g150(.a(new_n241), .b(new_n189), .c(new_n191), .o1(new_n246));
  xnrc02aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .out0(new_n247));
  aoib12aa1n03x5               g152(.a(new_n247), .b(new_n246), .c(new_n239), .out0(new_n248));
  nor042aa1n04x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  nand42aa1n04x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  norb02aa1n12x5               g155(.a(new_n250), .b(new_n249), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  nano22aa1n03x7               g157(.a(new_n248), .b(new_n245), .c(new_n252), .out0(new_n253));
  oaoi13aa1n02x5               g158(.a(new_n252), .b(new_n245), .c(new_n242), .d(new_n247), .o1(new_n254));
  norp02aa1n02x5               g159(.a(new_n254), .b(new_n253), .o1(\s[24] ));
  norb02aa1n06x4               g160(.a(new_n251), .b(new_n247), .out0(new_n256));
  nano22aa1n02x4               g161(.a(new_n229), .b(new_n237), .c(new_n256), .out0(new_n257));
  aoi122aa1n06x5               g162(.a(new_n249), .b(new_n250), .c(new_n244), .d(new_n256), .e(new_n238), .o1(new_n258));
  nand23aa1n06x5               g163(.a(new_n225), .b(new_n237), .c(new_n256), .o1(new_n259));
  nanp02aa1n09x5               g164(.a(new_n259), .b(new_n258), .o1(new_n260));
  oaoi13aa1n06x5               g165(.a(new_n260), .b(new_n257), .c(new_n189), .d(new_n191), .o1(new_n261));
  xnrb03aa1n03x5               g166(.a(new_n261), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  oaih12aa1n02x5               g169(.a(new_n257), .b(new_n189), .c(new_n191), .o1(new_n265));
  xnrc02aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .out0(new_n266));
  aoib12aa1n02x5               g171(.a(new_n266), .b(new_n265), .c(new_n260), .out0(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  nano22aa1n02x5               g173(.a(new_n267), .b(new_n264), .c(new_n268), .out0(new_n269));
  oaoi13aa1n02x5               g174(.a(new_n268), .b(new_n264), .c(new_n261), .d(new_n266), .o1(new_n270));
  norp02aa1n02x5               g175(.a(new_n270), .b(new_n269), .o1(\s[26] ));
  nor042aa1n02x5               g176(.a(new_n268), .b(new_n266), .o1(new_n272));
  nano22aa1d15x5               g177(.a(new_n240), .b(new_n256), .c(new_n272), .out0(new_n273));
  oai012aa1n04x7               g178(.a(new_n273), .b(new_n189), .c(new_n191), .o1(new_n274));
  oao003aa1n03x5               g179(.a(\a[26] ), .b(\b[25] ), .c(new_n264), .carry(new_n275));
  aobi12aa1n12x5               g180(.a(new_n275), .b(new_n260), .c(new_n272), .out0(new_n276));
  nor042aa1n03x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n278), .b(new_n277), .out0(new_n279));
  xnbna2aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n274), .out0(\s[27] ));
  inv000aa1d42x5               g185(.a(new_n277), .o1(new_n281));
  xnrc02aa1n02x5               g186(.a(\b[27] ), .b(\a[28] ), .out0(new_n282));
  nano23aa1n02x4               g187(.a(new_n165), .b(new_n179), .c(new_n180), .d(new_n166), .out0(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n170), .c(new_n154), .d(new_n168), .o1(new_n284));
  nano32aa1n02x4               g189(.a(new_n141), .b(new_n283), .c(new_n173), .d(new_n168), .out0(new_n285));
  aoai13aa1n02x5               g190(.a(new_n285), .b(new_n125), .c(new_n110), .d(new_n118), .o1(new_n286));
  nanp03aa1n02x5               g191(.a(new_n286), .b(new_n284), .c(new_n188), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n272), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n275), .b(new_n288), .c(new_n259), .d(new_n258), .o1(new_n289));
  aoai13aa1n02x7               g194(.a(new_n278), .b(new_n289), .c(new_n287), .d(new_n273), .o1(new_n290));
  aoi012aa1n02x7               g195(.a(new_n282), .b(new_n290), .c(new_n281), .o1(new_n291));
  aobi12aa1n03x5               g196(.a(new_n278), .b(new_n276), .c(new_n274), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n281), .c(new_n282), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[28] ));
  nano22aa1n02x4               g199(.a(new_n282), .b(new_n281), .c(new_n278), .out0(new_n295));
  aoai13aa1n02x5               g200(.a(new_n295), .b(new_n289), .c(new_n287), .d(new_n273), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n281), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[28] ), .b(\a[29] ), .out0(new_n298));
  aoi012aa1n02x7               g203(.a(new_n298), .b(new_n296), .c(new_n297), .o1(new_n299));
  aobi12aa1n03x5               g204(.a(new_n295), .b(new_n276), .c(new_n274), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n297), .c(new_n298), .out0(new_n301));
  nor002aa1n02x5               g206(.a(new_n299), .b(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g208(.a(new_n279), .b(new_n298), .c(new_n282), .out0(new_n304));
  aoai13aa1n02x5               g209(.a(new_n304), .b(new_n289), .c(new_n287), .d(new_n273), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[29] ), .b(\a[30] ), .out0(new_n307));
  aoi012aa1n03x5               g212(.a(new_n307), .b(new_n305), .c(new_n306), .o1(new_n308));
  aobi12aa1n03x5               g213(.a(new_n304), .b(new_n276), .c(new_n274), .out0(new_n309));
  nano22aa1n03x5               g214(.a(new_n309), .b(new_n306), .c(new_n307), .out0(new_n310));
  norp02aa1n03x5               g215(.a(new_n308), .b(new_n310), .o1(\s[30] ));
  xnrc02aa1n02x5               g216(.a(\b[30] ), .b(\a[31] ), .out0(new_n312));
  norb03aa1n02x5               g217(.a(new_n295), .b(new_n307), .c(new_n298), .out0(new_n313));
  aobi12aa1n03x5               g218(.a(new_n313), .b(new_n276), .c(new_n274), .out0(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n315));
  nano22aa1n03x5               g220(.a(new_n314), .b(new_n312), .c(new_n315), .out0(new_n316));
  aoai13aa1n02x5               g221(.a(new_n313), .b(new_n289), .c(new_n287), .d(new_n273), .o1(new_n317));
  aoi012aa1n03x5               g222(.a(new_n312), .b(new_n317), .c(new_n315), .o1(new_n318));
  norp02aa1n03x5               g223(.a(new_n318), .b(new_n316), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n108), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n108), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g228(.a(\a[5] ), .o1(new_n324));
  inv000aa1d42x5               g229(.a(\b[4] ), .o1(new_n325));
  oaoi03aa1n02x5               g230(.a(new_n324), .b(new_n325), .c(new_n110), .o1(new_n326));
  xnrb03aa1n02x5               g231(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g232(.a(\a[6] ), .b(\b[5] ), .c(new_n326), .o1(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g234(.a(new_n113), .b(new_n328), .c(new_n114), .o1(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n330), .b(new_n132), .c(new_n112), .out0(\s[8] ));
  norb02aa1n02x5               g236(.a(new_n140), .b(new_n139), .out0(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n131), .c(new_n136), .out0(\s[9] ));
endmodule


