// Benchmark "adder" written by ABC on Thu Jul 18 05:54:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n328, new_n330, new_n333,
    new_n335, new_n336, new_n338, new_n339, new_n340, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[4] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[3] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(new_n101), .b(new_n102), .o1(new_n103));
  nand02aa1n08x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanb03aa1n09x5               g011(.a(new_n105), .b(new_n106), .c(new_n104), .out0(new_n107));
  nand02aa1d04x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nor002aa1n03x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  norb03aa1n12x5               g014(.a(new_n104), .b(new_n109), .c(new_n108), .out0(new_n110));
  oaoi03aa1n09x5               g015(.a(new_n99), .b(new_n100), .c(new_n105), .o1(new_n111));
  oai013aa1d12x5               g016(.a(new_n111), .b(new_n110), .c(new_n107), .d(new_n103), .o1(new_n112));
  nor002aa1n06x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1n06x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1d18x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nor002aa1n03x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nor042aa1n03x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nand22aa1n03x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nona23aa1n02x4               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  nor042aa1n03x5               g027(.a(new_n122), .b(new_n117), .o1(new_n123));
  tech160nm_fiaoi012aa1n04x5   g028(.a(new_n120), .b(new_n118), .c(new_n121), .o1(new_n124));
  oa0012aa1n02x5               g029(.a(new_n114), .b(new_n115), .c(new_n113), .o(new_n125));
  oabi12aa1n18x5               g030(.a(new_n125), .b(new_n117), .c(new_n124), .out0(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n126), .c(new_n112), .d(new_n123), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  nor002aa1n03x5               g035(.a(new_n107), .b(new_n103), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n110), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n111), .o1(new_n133));
  aoai13aa1n06x5               g038(.a(new_n123), .b(new_n133), .c(new_n131), .d(new_n132), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n126), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(new_n129), .b(new_n127), .o1(new_n136));
  norp02aa1n02x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nanp02aa1n02x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  tech160nm_fioai012aa1n05x5   g043(.a(new_n138), .b(new_n137), .c(new_n97), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n136), .c(new_n134), .d(new_n135), .o1(new_n140));
  xorb03aa1n02x5               g045(.a(new_n140), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n09x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  nand42aa1n06x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n142), .out0(new_n145));
  nanp02aa1n03x5               g050(.a(new_n140), .b(new_n145), .o1(new_n146));
  nor042aa1n02x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  xnbna2aa1n03x5               g054(.a(new_n149), .b(new_n146), .c(new_n143), .out0(\s[12] ));
  tech160nm_fiaoi012aa1n05x5   g055(.a(new_n126), .b(new_n112), .c(new_n123), .o1(new_n151));
  nano23aa1n03x5               g056(.a(new_n142), .b(new_n147), .c(new_n148), .d(new_n144), .out0(new_n152));
  nand23aa1n03x5               g057(.a(new_n152), .b(new_n127), .c(new_n129), .o1(new_n153));
  nona23aa1n09x5               g058(.a(new_n148), .b(new_n144), .c(new_n142), .d(new_n147), .out0(new_n154));
  tech160nm_fioai012aa1n04x5   g059(.a(new_n148), .b(new_n147), .c(new_n142), .o1(new_n155));
  tech160nm_fioai012aa1n05x5   g060(.a(new_n155), .b(new_n154), .c(new_n139), .o1(new_n156));
  oabi12aa1n02x5               g061(.a(new_n156), .b(new_n151), .c(new_n153), .out0(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand02aa1n03x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nano22aa1n02x4               g065(.a(new_n159), .b(new_n157), .c(new_n160), .out0(new_n161));
  nor042aa1n04x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand22aa1n03x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n159), .c(new_n157), .d(new_n160), .o1(new_n165));
  nona22aa1n02x4               g070(.a(new_n163), .b(new_n162), .c(new_n159), .out0(new_n166));
  oai012aa1n02x5               g071(.a(new_n165), .b(new_n161), .c(new_n166), .o1(\s[14] ));
  nona23aa1n06x5               g072(.a(new_n163), .b(new_n160), .c(new_n159), .d(new_n162), .out0(new_n168));
  nano23aa1n06x5               g073(.a(new_n159), .b(new_n162), .c(new_n163), .d(new_n160), .out0(new_n169));
  aoi022aa1n02x5               g074(.a(new_n156), .b(new_n169), .c(new_n163), .d(new_n166), .o1(new_n170));
  oai013aa1n03x5               g075(.a(new_n170), .b(new_n151), .c(new_n153), .d(new_n168), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand02aa1n06x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nanb02aa1n18x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  norp02aa1n12x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand02aa1n03x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n03x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  aoai13aa1n02x5               g084(.a(new_n179), .b(new_n173), .c(new_n171), .d(new_n176), .o1(new_n180));
  nona22aa1n02x4               g085(.a(new_n178), .b(new_n177), .c(new_n173), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n180), .b(new_n181), .c(new_n176), .d(new_n171), .o1(\s[16] ));
  nona22aa1n03x5               g087(.a(new_n169), .b(new_n175), .c(new_n179), .out0(new_n183));
  nor042aa1n03x5               g088(.a(new_n153), .b(new_n183), .o1(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n126), .c(new_n112), .d(new_n123), .o1(new_n185));
  nona23aa1n02x4               g090(.a(new_n178), .b(new_n174), .c(new_n173), .d(new_n177), .out0(new_n186));
  nor042aa1n02x5               g091(.a(new_n186), .b(new_n168), .o1(new_n187));
  oai012aa1n02x5               g092(.a(new_n163), .b(new_n162), .c(new_n159), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n178), .b(new_n177), .c(new_n173), .o1(new_n189));
  tech160nm_fioai012aa1n02p5x5 g094(.a(new_n189), .b(new_n186), .c(new_n188), .o1(new_n190));
  aoi012aa1n12x5               g095(.a(new_n190), .b(new_n156), .c(new_n187), .o1(new_n191));
  xnrc02aa1n12x5               g096(.a(\b[16] ), .b(\a[17] ), .out0(new_n192));
  xobna2aa1n03x5               g097(.a(new_n192), .b(new_n185), .c(new_n191), .out0(\s[17] ));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  nona22aa1n02x4               g100(.a(new_n187), .b(new_n136), .c(new_n154), .out0(new_n196));
  aoai13aa1n09x5               g101(.a(new_n191), .b(new_n196), .c(new_n134), .d(new_n135), .o1(new_n197));
  oaoi03aa1n02x5               g102(.a(new_n194), .b(new_n195), .c(new_n197), .o1(new_n198));
  nor002aa1d32x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  tech160nm_finand02aa1n03p5x5 g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nanb02aa1n09x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  nor002aa1n12x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  norb03aa1n02x5               g107(.a(new_n200), .b(new_n202), .c(new_n199), .out0(new_n203));
  aoai13aa1n02x5               g108(.a(new_n203), .b(new_n192), .c(new_n185), .d(new_n191), .o1(new_n204));
  oaib12aa1n02x5               g109(.a(new_n204), .b(new_n198), .c(new_n201), .out0(\s[18] ));
  nor042aa1n06x5               g110(.a(new_n192), .b(new_n201), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  and002aa1n12x5               g112(.a(\b[17] ), .b(\a[18] ), .o(new_n208));
  oab012aa1d15x5               g113(.a(new_n208), .b(new_n202), .c(new_n199), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n207), .c(new_n185), .d(new_n191), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n12x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand42aa1d28x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nor042aa1n09x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand42aa1d28x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanb02aa1n02x5               g122(.a(new_n216), .b(new_n217), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n214), .c(new_n211), .d(new_n215), .o1(new_n219));
  nanp02aa1n03x5               g124(.a(new_n197), .b(new_n206), .o1(new_n220));
  nanb02aa1n02x5               g125(.a(new_n214), .b(new_n215), .out0(new_n221));
  norb03aa1n02x5               g126(.a(new_n217), .b(new_n214), .c(new_n216), .out0(new_n222));
  aoai13aa1n03x5               g127(.a(new_n222), .b(new_n221), .c(new_n220), .d(new_n210), .o1(new_n223));
  nanp02aa1n03x5               g128(.a(new_n219), .b(new_n223), .o1(\s[20] ));
  nano23aa1d15x5               g129(.a(new_n214), .b(new_n216), .c(new_n217), .d(new_n215), .out0(new_n225));
  norb03aa1n12x5               g130(.a(new_n225), .b(new_n192), .c(new_n201), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nand22aa1n09x5               g132(.a(new_n225), .b(new_n209), .o1(new_n228));
  oai012aa1d24x5               g133(.a(new_n217), .b(new_n216), .c(new_n214), .o1(new_n229));
  nand42aa1n04x5               g134(.a(new_n228), .b(new_n229), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n227), .c(new_n185), .d(new_n191), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n12x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  nand22aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n235), .b(new_n234), .out0(new_n236));
  nor042aa1n12x5               g141(.a(\b[21] ), .b(\a[22] ), .o1(new_n237));
  nand22aa1n12x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n238), .b(new_n237), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n232), .d(new_n236), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n236), .b(new_n230), .c(new_n197), .d(new_n226), .o1(new_n242));
  nona22aa1n03x5               g147(.a(new_n242), .b(new_n240), .c(new_n234), .out0(new_n243));
  nanp02aa1n02x5               g148(.a(new_n241), .b(new_n243), .o1(\s[22] ));
  nano23aa1n06x5               g149(.a(new_n234), .b(new_n237), .c(new_n238), .d(new_n235), .out0(new_n245));
  nona23aa1n02x4               g150(.a(new_n245), .b(new_n225), .c(new_n192), .d(new_n201), .out0(new_n246));
  inv000aa1n02x5               g151(.a(new_n238), .o1(new_n247));
  oab012aa1n03x5               g152(.a(new_n247), .b(new_n234), .c(new_n237), .out0(new_n248));
  tech160nm_fiaoi012aa1n03p5x5 g153(.a(new_n248), .b(new_n230), .c(new_n245), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n246), .c(new_n185), .d(new_n191), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1d32x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  nand42aa1n06x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  norb02aa1n02x5               g158(.a(new_n253), .b(new_n252), .out0(new_n254));
  nor002aa1d32x5               g159(.a(\b[23] ), .b(\a[24] ), .o1(new_n255));
  nand42aa1d28x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n02x5               g163(.a(new_n258), .b(new_n252), .c(new_n250), .d(new_n254), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(new_n250), .b(new_n254), .o1(new_n260));
  nona22aa1d36x5               g165(.a(new_n256), .b(new_n255), .c(new_n252), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(new_n260), .b(new_n262), .o1(new_n263));
  nanp02aa1n03x5               g168(.a(new_n259), .b(new_n263), .o1(\s[24] ));
  nano23aa1n09x5               g169(.a(new_n252), .b(new_n255), .c(new_n256), .d(new_n253), .out0(new_n265));
  nand22aa1n09x5               g170(.a(new_n265), .b(new_n245), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  nanp02aa1n02x5               g172(.a(new_n226), .b(new_n267), .o1(new_n268));
  aoi022aa1n12x5               g173(.a(new_n265), .b(new_n248), .c(new_n256), .d(new_n261), .o1(new_n269));
  aoai13aa1n12x5               g174(.a(new_n269), .b(new_n266), .c(new_n228), .d(new_n229), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n268), .c(new_n185), .d(new_n191), .o1(new_n272));
  xorb03aa1n02x5               g177(.a(new_n272), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  inv000aa1d42x5               g178(.a(new_n225), .o1(new_n274));
  nona32aa1n03x5               g179(.a(new_n197), .b(new_n266), .c(new_n274), .d(new_n207), .out0(new_n275));
  xnrc02aa1n12x5               g180(.a(\b[24] ), .b(\a[25] ), .out0(new_n276));
  aoi012aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n271), .o1(new_n277));
  norp02aa1n02x5               g182(.a(\b[24] ), .b(\a[25] ), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n276), .o1(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[25] ), .b(\a[26] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n278), .c(new_n272), .d(new_n279), .o1(new_n281));
  oabi12aa1n02x5               g186(.a(new_n280), .b(\a[25] ), .c(\b[24] ), .out0(new_n282));
  oai012aa1n02x5               g187(.a(new_n281), .b(new_n277), .c(new_n282), .o1(\s[26] ));
  nor002aa1n02x5               g188(.a(new_n280), .b(new_n276), .o1(new_n284));
  nano32aa1n03x7               g189(.a(new_n266), .b(new_n284), .c(new_n206), .d(new_n225), .out0(new_n285));
  inv000aa1n02x5               g190(.a(new_n285), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(\b[25] ), .b(\a[26] ), .o1(new_n287));
  aoi022aa1n06x5               g192(.a(new_n270), .b(new_n284), .c(new_n287), .d(new_n282), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n286), .c(new_n185), .d(new_n191), .o1(new_n289));
  xorb03aa1n03x5               g194(.a(new_n289), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n291), .c(new_n289), .d(new_n292), .o1(new_n294));
  nanp02aa1n03x5               g199(.a(new_n270), .b(new_n284), .o1(new_n295));
  oai012aa1n02x5               g200(.a(new_n287), .b(new_n280), .c(new_n278), .o1(new_n296));
  nanp02aa1n03x5               g201(.a(new_n295), .b(new_n296), .o1(new_n297));
  aoai13aa1n02x7               g202(.a(new_n292), .b(new_n297), .c(new_n197), .d(new_n285), .o1(new_n298));
  nona22aa1n03x5               g203(.a(new_n298), .b(new_n293), .c(new_n291), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n294), .b(new_n299), .o1(\s[28] ));
  norb02aa1n02x5               g205(.a(new_n292), .b(new_n293), .out0(new_n301));
  aoai13aa1n02x7               g206(.a(new_n301), .b(new_n297), .c(new_n197), .d(new_n285), .o1(new_n302));
  tech160nm_fixorc02aa1n03p5x5 g207(.a(\a[29] ), .b(\b[28] ), .out0(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  inv000aa1d42x5               g209(.a(\a[28] ), .o1(new_n305));
  inv000aa1d42x5               g210(.a(\b[27] ), .o1(new_n306));
  oao003aa1n02x5               g211(.a(new_n305), .b(new_n306), .c(new_n291), .carry(new_n307));
  nona22aa1n03x5               g212(.a(new_n302), .b(new_n304), .c(new_n307), .out0(new_n308));
  aoai13aa1n02x7               g213(.a(new_n304), .b(new_n307), .c(new_n289), .d(new_n301), .o1(new_n309));
  nanp02aa1n03x5               g214(.a(new_n309), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g215(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g216(.a(new_n293), .b(new_n292), .c(new_n303), .out0(new_n312));
  inv000aa1n03x5               g217(.a(new_n307), .o1(new_n313));
  oaoi03aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .o1(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[29] ), .b(\a[30] ), .out0(new_n315));
  aoai13aa1n02x7               g220(.a(new_n315), .b(new_n314), .c(new_n289), .d(new_n312), .o1(new_n316));
  aoai13aa1n02x7               g221(.a(new_n312), .b(new_n297), .c(new_n197), .d(new_n285), .o1(new_n317));
  nona22aa1n02x4               g222(.a(new_n317), .b(new_n314), .c(new_n315), .out0(new_n318));
  nanp02aa1n03x5               g223(.a(new_n316), .b(new_n318), .o1(\s[30] ));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nano23aa1n02x4               g225(.a(new_n315), .b(new_n293), .c(new_n292), .d(new_n303), .out0(new_n321));
  and002aa1n02x5               g226(.a(\b[29] ), .b(\a[30] ), .o(new_n322));
  oab012aa1n02x4               g227(.a(new_n322), .b(new_n314), .c(new_n315), .out0(new_n323));
  aoai13aa1n02x7               g228(.a(new_n320), .b(new_n323), .c(new_n289), .d(new_n321), .o1(new_n324));
  aoai13aa1n02x7               g229(.a(new_n321), .b(new_n297), .c(new_n197), .d(new_n285), .o1(new_n325));
  nona22aa1n02x4               g230(.a(new_n325), .b(new_n323), .c(new_n320), .out0(new_n326));
  nanp02aa1n03x5               g231(.a(new_n324), .b(new_n326), .o1(\s[31] ));
  oai012aa1n02x5               g232(.a(new_n104), .b(new_n109), .c(new_n108), .o1(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g234(.a(\a[3] ), .b(\b[2] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g236(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n04x7               g237(.a(new_n119), .b(new_n112), .c(new_n118), .o1(new_n333));
  xnrb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g239(.a(new_n115), .b(new_n116), .out0(new_n335));
  nanb03aa1n03x5               g240(.a(new_n120), .b(new_n333), .c(new_n121), .out0(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n335), .b(new_n336), .c(new_n121), .out0(\s[7] ));
  nona22aa1n02x4               g242(.a(new_n114), .b(new_n115), .c(new_n113), .out0(new_n338));
  nano22aa1n02x4               g243(.a(new_n115), .b(new_n116), .c(new_n121), .out0(new_n339));
  nanb02aa1n02x5               g244(.a(new_n113), .b(new_n114), .out0(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n115), .c(new_n336), .d(new_n339), .o1(new_n341));
  aoai13aa1n02x5               g246(.a(new_n341), .b(new_n338), .c(new_n339), .d(new_n336), .o1(\s[8] ));
  xnbna2aa1n03x5               g247(.a(new_n127), .b(new_n134), .c(new_n135), .out0(\s[9] ));
endmodule


