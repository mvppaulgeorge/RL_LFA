// Benchmark "adder" written by ABC on Wed Jul 17 15:54:11 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n320, new_n323, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  tech160nm_finor002aa1n03p5x5 g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  tech160nm_fiaoi012aa1n05x5   g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor002aa1n06x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1d06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  tech160nm_fiaoi012aa1n04x5   g012(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n108));
  oai012aa1n06x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nor022aa1n08x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand42aa1n04x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nor002aa1n12x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n09x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .d(new_n110), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  nor043aa1n02x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  inv040aa1d32x5               g022(.a(\a[5] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[4] ), .o1(new_n119));
  nand42aa1n04x5               g024(.a(new_n119), .b(new_n118), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[6] ), .b(\b[5] ), .c(new_n120), .o1(new_n121));
  aoi012aa1n02x7               g026(.a(new_n110), .b(new_n113), .c(new_n111), .o1(new_n122));
  oaib12aa1n06x5               g027(.a(new_n122), .b(new_n114), .c(new_n121), .out0(new_n123));
  nand42aa1n04x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n97), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n126));
  nor002aa1d32x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n20x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  nor042aa1n04x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nand42aa1n06x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n127), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n128), .o1(new_n135));
  aoai13aa1n06x5               g040(.a(new_n134), .b(new_n135), .c(new_n126), .d(new_n98), .o1(new_n136));
  nano23aa1n03x5               g041(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n137));
  nanb02aa1n02x5               g042(.a(new_n102), .b(new_n137), .out0(new_n138));
  nano23aa1n03x5               g043(.a(new_n113), .b(new_n110), .c(new_n111), .d(new_n112), .out0(new_n139));
  nona22aa1n02x4               g044(.a(new_n139), .b(new_n115), .c(new_n116), .out0(new_n140));
  aobi12aa1n02x7               g045(.a(new_n122), .b(new_n139), .c(new_n121), .out0(new_n141));
  aoai13aa1n04x5               g046(.a(new_n141), .b(new_n140), .c(new_n138), .d(new_n108), .o1(new_n142));
  norp02aa1n06x5               g047(.a(new_n127), .b(new_n97), .o1(new_n143));
  inv040aa1n04x5               g048(.a(new_n143), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n128), .b(new_n144), .c(new_n142), .d(new_n125), .o1(new_n145));
  mtn022aa1n02x5               g050(.a(new_n136), .b(new_n145), .sa(new_n133), .o1(\s[11] ));
  xorc02aa1n12x5               g051(.a(\a[12] ), .b(\b[11] ), .out0(new_n147));
  aoi112aa1n02x5               g052(.a(new_n147), .b(new_n131), .c(new_n136), .d(new_n133), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n147), .b(new_n131), .c(new_n136), .d(new_n132), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(\s[12] ));
  nano22aa1d15x5               g055(.a(new_n131), .b(new_n128), .c(new_n132), .out0(new_n151));
  norb03aa1d15x5               g056(.a(new_n124), .b(new_n97), .c(new_n127), .out0(new_n152));
  nand23aa1n09x5               g057(.a(new_n151), .b(new_n147), .c(new_n152), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n155));
  nand23aa1n06x5               g060(.a(new_n151), .b(new_n147), .c(new_n144), .o1(new_n156));
  aoi112aa1n03x5               g061(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n157));
  oab012aa1n06x5               g062(.a(new_n157), .b(\a[12] ), .c(\b[11] ), .out0(new_n158));
  nand22aa1n09x5               g063(.a(new_n156), .b(new_n158), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  xorc02aa1n12x5               g065(.a(\a[13] ), .b(\b[12] ), .out0(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n155), .c(new_n160), .out0(\s[13] ));
  orn002aa1n24x5               g067(.a(\a[13] ), .b(\b[12] ), .o(new_n163));
  xnrc02aa1n02x5               g068(.a(\b[12] ), .b(\a[13] ), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n163), .b(new_n164), .c(new_n155), .d(new_n160), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xorc02aa1n12x5               g071(.a(\a[14] ), .b(\b[13] ), .out0(new_n167));
  nand02aa1d06x5               g072(.a(new_n167), .b(new_n161), .o1(new_n168));
  oaoi03aa1n12x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n169));
  inv000aa1n02x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n168), .c(new_n155), .d(new_n160), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  xorc02aa1n12x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  xorc02aa1n12x5               g079(.a(\a[16] ), .b(\b[15] ), .out0(new_n175));
  aoi112aa1n02x5               g080(.a(new_n173), .b(new_n175), .c(new_n171), .d(new_n174), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n175), .b(new_n173), .c(new_n171), .d(new_n174), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(\s[16] ));
  tech160nm_finand02aa1n05x5   g083(.a(new_n175), .b(new_n174), .o1(new_n179));
  nor043aa1d12x5               g084(.a(new_n153), .b(new_n168), .c(new_n179), .o1(new_n180));
  aoai13aa1n06x5               g085(.a(new_n180), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n181));
  nano22aa1n02x5               g086(.a(new_n168), .b(new_n174), .c(new_n175), .out0(new_n182));
  inv000aa1d42x5               g087(.a(new_n173), .o1(new_n183));
  tech160nm_fioaoi03aa1n03p5x5 g088(.a(\a[16] ), .b(\b[15] ), .c(new_n183), .o1(new_n184));
  oabi12aa1n06x5               g089(.a(new_n184), .b(new_n179), .c(new_n170), .out0(new_n185));
  aoi012aa1n12x5               g090(.a(new_n185), .b(new_n159), .c(new_n182), .o1(new_n186));
  nand02aa1d08x5               g091(.a(new_n181), .b(new_n186), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[16] ), .o1(new_n191));
  oaoi03aa1n02x5               g096(.a(new_n190), .b(new_n191), .c(new_n187), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(new_n189), .out0(\s[18] ));
  xroi22aa1d06x4               g098(.a(new_n190), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n194));
  oai022aa1d18x5               g099(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n195));
  oaib12aa1n06x5               g100(.a(new_n195), .b(new_n189), .c(\b[17] ), .out0(new_n196));
  inv000aa1n06x5               g101(.a(new_n196), .o1(new_n197));
  nor002aa1d32x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand22aa1n12x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n201));
  aoi112aa1n02x5               g106(.a(new_n200), .b(new_n197), .c(new_n187), .d(new_n194), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n201), .b(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n06x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand22aa1n09x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  nona22aa1n03x5               g112(.a(new_n201), .b(new_n207), .c(new_n198), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n198), .o1(new_n209));
  aobi12aa1n06x5               g114(.a(new_n207), .b(new_n201), .c(new_n209), .out0(new_n210));
  norb02aa1n03x4               g115(.a(new_n208), .b(new_n210), .out0(\s[20] ));
  nano23aa1n06x5               g116(.a(new_n198), .b(new_n205), .c(new_n206), .d(new_n199), .out0(new_n212));
  nand22aa1n04x5               g117(.a(new_n194), .b(new_n212), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nona23aa1n03x5               g119(.a(new_n206), .b(new_n199), .c(new_n198), .d(new_n205), .out0(new_n215));
  aoi012aa1n02x7               g120(.a(new_n205), .b(new_n198), .c(new_n206), .o1(new_n216));
  tech160nm_fioai012aa1n05x5   g121(.a(new_n216), .b(new_n215), .c(new_n196), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n217), .c(new_n187), .d(new_n214), .o1(new_n219));
  aoi112aa1n02x5               g124(.a(new_n218), .b(new_n217), .c(new_n187), .d(new_n214), .o1(new_n220));
  norb02aa1n02x5               g125(.a(new_n219), .b(new_n220), .out0(\s[21] ));
  xnrc02aa1n02x5               g126(.a(\b[21] ), .b(\a[22] ), .out0(new_n222));
  oai112aa1n03x5               g127(.a(new_n219), .b(new_n222), .c(\b[20] ), .d(\a[21] ), .o1(new_n223));
  oaoi13aa1n06x5               g128(.a(new_n222), .b(new_n219), .c(\a[21] ), .d(\b[20] ), .o1(new_n224));
  norb02aa1n03x4               g129(.a(new_n223), .b(new_n224), .out0(\s[22] ));
  inv000aa1d42x5               g130(.a(\a[21] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  and003aa1n02x5               g133(.a(new_n194), .b(new_n228), .c(new_n212), .o(new_n229));
  inv020aa1n03x5               g134(.a(new_n216), .o1(new_n230));
  aoai13aa1n06x5               g135(.a(new_n228), .b(new_n230), .c(new_n212), .d(new_n197), .o1(new_n231));
  inv040aa1d32x5               g136(.a(\b[21] ), .o1(new_n232));
  nor042aa1n03x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  oao003aa1n02x5               g138(.a(new_n227), .b(new_n232), .c(new_n233), .carry(new_n234));
  inv030aa1n02x5               g139(.a(new_n234), .o1(new_n235));
  nanp02aa1n02x5               g140(.a(new_n231), .b(new_n235), .o1(new_n236));
  xorc02aa1n02x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n236), .c(new_n187), .d(new_n229), .o1(new_n238));
  aoi112aa1n02x5               g143(.a(new_n237), .b(new_n236), .c(new_n187), .d(new_n229), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(\s[23] ));
  xorc02aa1n02x5               g145(.a(\a[24] ), .b(\b[23] ), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  oai112aa1n03x5               g147(.a(new_n238), .b(new_n242), .c(\b[22] ), .d(\a[23] ), .o1(new_n243));
  oaoi13aa1n06x5               g148(.a(new_n242), .b(new_n238), .c(\a[23] ), .d(\b[22] ), .o1(new_n244));
  norb02aa1n03x4               g149(.a(new_n243), .b(new_n244), .out0(\s[24] ));
  xnrc02aa1n02x5               g150(.a(\b[14] ), .b(\a[15] ), .out0(new_n246));
  nona23aa1n02x4               g151(.a(new_n175), .b(new_n167), .c(new_n164), .d(new_n246), .out0(new_n247));
  aoi013aa1n02x4               g152(.a(new_n184), .b(new_n169), .c(new_n174), .d(new_n175), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n247), .c(new_n156), .d(new_n158), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\a[23] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\a[24] ), .o1(new_n251));
  xroi22aa1d06x4               g156(.a(new_n250), .b(\b[22] ), .c(new_n251), .d(\b[23] ), .out0(new_n252));
  nano22aa1n03x7               g157(.a(new_n213), .b(new_n228), .c(new_n252), .out0(new_n253));
  aoai13aa1n02x5               g158(.a(new_n253), .b(new_n249), .c(new_n142), .d(new_n180), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n252), .o1(new_n255));
  aoi112aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n256));
  aoib12aa1n06x5               g161(.a(new_n256), .b(new_n251), .c(\b[23] ), .out0(new_n257));
  aoai13aa1n12x5               g162(.a(new_n257), .b(new_n255), .c(new_n231), .d(new_n235), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[24] ), .b(\a[25] ), .out0(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n254), .c(new_n259), .out0(\s[25] ));
  nor042aa1n03x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aoai13aa1n04x5               g169(.a(new_n261), .b(new_n258), .c(new_n187), .d(new_n253), .o1(new_n265));
  xnrc02aa1n06x5               g170(.a(\b[25] ), .b(\a[26] ), .out0(new_n266));
  nand03aa1n02x5               g171(.a(new_n265), .b(new_n264), .c(new_n266), .o1(new_n267));
  aoi012aa1n02x7               g172(.a(new_n266), .b(new_n265), .c(new_n264), .o1(new_n268));
  norb02aa1n02x7               g173(.a(new_n267), .b(new_n268), .out0(\s[26] ));
  nor042aa1n06x5               g174(.a(new_n266), .b(new_n260), .o1(new_n270));
  nano32aa1n03x7               g175(.a(new_n213), .b(new_n270), .c(new_n228), .d(new_n252), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n249), .c(new_n142), .d(new_n180), .o1(new_n272));
  nand02aa1d10x5               g177(.a(new_n258), .b(new_n270), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .c(new_n264), .carry(new_n274));
  xorc02aa1n12x5               g179(.a(\a[27] ), .b(\b[26] ), .out0(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoi013aa1n06x4               g181(.a(new_n276), .b(new_n272), .c(new_n273), .d(new_n274), .o1(new_n277));
  aobi12aa1n06x5               g182(.a(new_n271), .b(new_n181), .c(new_n186), .out0(new_n278));
  aoai13aa1n03x5               g183(.a(new_n252), .b(new_n234), .c(new_n217), .d(new_n228), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n270), .o1(new_n280));
  aoai13aa1n04x5               g185(.a(new_n274), .b(new_n280), .c(new_n279), .d(new_n257), .o1(new_n281));
  norp03aa1n02x5               g186(.a(new_n281), .b(new_n278), .c(new_n275), .o1(new_n282));
  nor002aa1n02x5               g187(.a(new_n277), .b(new_n282), .o1(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  xnrc02aa1n12x5               g190(.a(\b[27] ), .b(\a[28] ), .out0(new_n286));
  nano22aa1n03x7               g191(.a(new_n277), .b(new_n285), .c(new_n286), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n275), .b(new_n281), .c(new_n278), .o1(new_n288));
  aoi012aa1n02x5               g193(.a(new_n286), .b(new_n288), .c(new_n285), .o1(new_n289));
  norp02aa1n03x5               g194(.a(new_n289), .b(new_n287), .o1(\s[28] ));
  norb02aa1d21x5               g195(.a(new_n275), .b(new_n286), .out0(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoi013aa1n02x5               g197(.a(new_n292), .b(new_n272), .c(new_n273), .d(new_n274), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  nano22aa1n03x5               g200(.a(new_n293), .b(new_n294), .c(new_n295), .out0(new_n296));
  tech160nm_fioai012aa1n03p5x5 g201(.a(new_n291), .b(new_n281), .c(new_n278), .o1(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n295), .b(new_n297), .c(new_n294), .o1(new_n298));
  norp02aa1n03x5               g203(.a(new_n298), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g205(.a(new_n275), .b(new_n295), .c(new_n286), .out0(new_n301));
  oai012aa1n02x5               g206(.a(new_n301), .b(new_n281), .c(new_n278), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[29] ), .b(\a[30] ), .out0(new_n304));
  aoi012aa1n02x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n301), .o1(new_n306));
  aoi013aa1n02x5               g211(.a(new_n306), .b(new_n272), .c(new_n273), .d(new_n274), .o1(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n304), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n305), .b(new_n308), .o1(\s[30] ));
  norb02aa1n02x5               g214(.a(new_n301), .b(new_n304), .out0(new_n310));
  inv000aa1n02x5               g215(.a(new_n310), .o1(new_n311));
  aoi013aa1n02x5               g216(.a(new_n311), .b(new_n272), .c(new_n273), .d(new_n274), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .c(new_n303), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[30] ), .b(\a[31] ), .out0(new_n314));
  nano22aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n314), .out0(new_n315));
  oai012aa1n02x7               g220(.a(new_n310), .b(new_n281), .c(new_n278), .o1(new_n316));
  aoi012aa1n02x5               g221(.a(new_n314), .b(new_n316), .c(new_n313), .o1(new_n317));
  norp02aa1n03x5               g222(.a(new_n317), .b(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g223(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g224(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g226(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g227(.a(new_n118), .b(new_n119), .c(new_n109), .o1(new_n323));
  xnrb03aa1n02x5               g228(.a(new_n323), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g229(.a(\a[6] ), .b(\b[5] ), .c(new_n323), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g231(.a(new_n113), .b(new_n325), .c(new_n112), .o1(new_n327));
  xnrb03aa1n02x5               g232(.a(new_n327), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n142), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


