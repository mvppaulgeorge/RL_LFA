// Benchmark "adder" written by ABC on Thu Jul 18 12:08:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n320, new_n323, new_n324, new_n325, new_n326,
    new_n328, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1d32x5               g002(.a(\b[6] ), .b(\a[7] ), .o1(new_n98));
  inv030aa1n04x5               g003(.a(new_n98), .o1(new_n99));
  oaoi03aa1n03x5               g004(.a(\a[8] ), .b(\b[7] ), .c(new_n99), .o1(new_n100));
  nor042aa1n03x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  nor042aa1n06x5               g006(.a(\b[4] ), .b(\a[5] ), .o1(new_n102));
  nand22aa1n06x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  aoi012aa1n06x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nanp02aa1n04x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nanp02aa1n06x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nona23aa1d18x5               g012(.a(new_n106), .b(new_n107), .c(new_n98), .d(new_n105), .out0(new_n108));
  oabi12aa1n18x5               g013(.a(new_n100), .b(new_n108), .c(new_n104), .out0(new_n109));
  inv040aa1n02x5               g014(.a(new_n109), .o1(new_n110));
  inv040aa1d32x5               g015(.a(\a[4] ), .o1(new_n111));
  inv040aa1n18x5               g016(.a(\b[3] ), .o1(new_n112));
  nanp02aa1n06x5               g017(.a(new_n112), .b(new_n111), .o1(new_n113));
  nand22aa1n09x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nand02aa1d08x5               g019(.a(new_n113), .b(new_n114), .o1(new_n115));
  nor002aa1d32x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  tech160nm_fioaoi03aa1n03p5x5 g021(.a(new_n111), .b(new_n112), .c(new_n116), .o1(new_n117));
  nor042aa1n04x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  nand22aa1n09x5               g023(.a(\b[0] ), .b(\a[1] ), .o1(new_n119));
  nand22aa1n12x5               g024(.a(\b[1] ), .b(\a[2] ), .o1(new_n120));
  aoi012aa1d24x5               g025(.a(new_n118), .b(new_n119), .c(new_n120), .o1(new_n121));
  nanp02aa1n06x5               g026(.a(\b[2] ), .b(\a[3] ), .o1(new_n122));
  nanb02aa1n12x5               g027(.a(new_n116), .b(new_n122), .out0(new_n123));
  oai013aa1d12x5               g028(.a(new_n117), .b(new_n121), .c(new_n123), .d(new_n115), .o1(new_n124));
  xnrc02aa1n12x5               g029(.a(\b[5] ), .b(\a[6] ), .out0(new_n125));
  nand42aa1n02x5               g030(.a(\b[4] ), .b(\a[5] ), .o1(new_n126));
  nanb02aa1n09x5               g031(.a(new_n102), .b(new_n126), .out0(new_n127));
  nor043aa1d12x5               g032(.a(new_n108), .b(new_n127), .c(new_n125), .o1(new_n128));
  nand42aa1n02x5               g033(.a(new_n124), .b(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(new_n129), .b(new_n110), .o1(new_n130));
  nand02aa1d28x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  aoi012aa1n02x5               g036(.a(new_n97), .b(new_n130), .c(new_n131), .o1(new_n132));
  xnrb03aa1n02x5               g037(.a(new_n132), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nand42aa1d28x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  aoi012aa1d24x5               g040(.a(new_n134), .b(new_n97), .c(new_n135), .o1(new_n136));
  nona23aa1n09x5               g041(.a(new_n135), .b(new_n131), .c(new_n97), .d(new_n134), .out0(new_n137));
  aoai13aa1n03x5               g042(.a(new_n136), .b(new_n137), .c(new_n129), .d(new_n110), .o1(new_n138));
  xorb03aa1n02x5               g043(.a(new_n138), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g044(.a(\a[12] ), .o1(new_n140));
  nor002aa1d32x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nand42aa1d28x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  aoi012aa1n03x5               g047(.a(new_n141), .b(new_n138), .c(new_n142), .o1(new_n143));
  xorb03aa1n02x5               g048(.a(new_n143), .b(\b[11] ), .c(new_n140), .out0(\s[12] ));
  nor002aa1d32x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand02aa1d28x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  aoi012aa1n12x5               g051(.a(new_n145), .b(new_n141), .c(new_n146), .o1(new_n147));
  nona23aa1d18x5               g052(.a(new_n146), .b(new_n142), .c(new_n141), .d(new_n145), .out0(new_n148));
  oai012aa1d24x5               g053(.a(new_n147), .b(new_n148), .c(new_n136), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nor002aa1n02x5               g055(.a(new_n148), .b(new_n137), .o1(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n109), .c(new_n124), .d(new_n128), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(new_n152), .b(new_n150), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g059(.a(\a[14] ), .o1(new_n155));
  nor002aa1d32x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1d28x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n156), .b(new_n153), .c(new_n157), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(new_n155), .out0(\s[14] ));
  nor002aa1d32x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1d28x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  aoi012aa1d24x5               g066(.a(new_n160), .b(new_n156), .c(new_n161), .o1(new_n162));
  nona23aa1d18x5               g067(.a(new_n161), .b(new_n157), .c(new_n156), .d(new_n160), .out0(new_n163));
  aoai13aa1n06x5               g068(.a(new_n162), .b(new_n163), .c(new_n152), .d(new_n150), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  tech160nm_fixorc02aa1n05x5   g071(.a(\a[15] ), .b(\b[14] ), .out0(new_n167));
  xnrc02aa1n12x5               g072(.a(\b[15] ), .b(\a[16] ), .out0(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n166), .c(new_n164), .d(new_n167), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(new_n164), .b(new_n167), .o1(new_n170));
  nona22aa1n02x5               g075(.a(new_n170), .b(new_n168), .c(new_n166), .out0(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n169), .o1(\s[16] ));
  xnrc02aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .out0(new_n173));
  inv040aa1n02x5               g078(.a(new_n166), .o1(new_n174));
  oao003aa1n03x5               g079(.a(\a[16] ), .b(\b[15] ), .c(new_n174), .carry(new_n175));
  oai013aa1n06x5               g080(.a(new_n175), .b(new_n168), .c(new_n173), .d(new_n162), .o1(new_n176));
  nor043aa1n09x5               g081(.a(new_n163), .b(new_n168), .c(new_n173), .o1(new_n177));
  aoi012aa1d24x5               g082(.a(new_n176), .b(new_n149), .c(new_n177), .o1(new_n178));
  nano23aa1n03x5               g083(.a(new_n97), .b(new_n134), .c(new_n135), .d(new_n131), .out0(new_n179));
  nano23aa1n06x5               g084(.a(new_n141), .b(new_n145), .c(new_n146), .d(new_n142), .out0(new_n180));
  nano23aa1n03x7               g085(.a(new_n156), .b(new_n160), .c(new_n161), .d(new_n157), .out0(new_n181));
  xorc02aa1n03x5               g086(.a(\a[16] ), .b(\b[15] ), .out0(new_n182));
  nand23aa1n02x5               g087(.a(new_n181), .b(new_n167), .c(new_n182), .o1(new_n183));
  nano22aa1n03x7               g088(.a(new_n183), .b(new_n179), .c(new_n180), .out0(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n109), .c(new_n124), .d(new_n128), .o1(new_n185));
  xorc02aa1n12x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n178), .out0(\s[17] ));
  nand22aa1n03x5               g092(.a(new_n177), .b(new_n151), .o1(new_n188));
  aoai13aa1n12x5               g093(.a(new_n178), .b(new_n188), .c(new_n129), .d(new_n110), .o1(new_n189));
  nor042aa1d18x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  tech160nm_fiaoi012aa1n05x5   g095(.a(new_n190), .b(new_n189), .c(new_n186), .o1(new_n191));
  inv040aa1d32x5               g096(.a(\a[18] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[17] ), .o1(new_n193));
  nand42aa1n10x5               g098(.a(new_n193), .b(new_n192), .o1(new_n194));
  nand02aa1d28x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n191), .b(new_n195), .c(new_n194), .out0(\s[18] ));
  aob012aa1d18x5               g101(.a(new_n194), .b(new_n190), .c(new_n195), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  inv000aa1n09x5               g103(.a(new_n186), .o1(new_n199));
  nano22aa1d15x5               g104(.a(new_n199), .b(new_n194), .c(new_n195), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n06x5               g106(.a(new_n198), .b(new_n201), .c(new_n185), .d(new_n178), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n12x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand02aa1n04x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nor042aa1n12x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nand02aa1d28x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n12x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n205), .c(new_n202), .d(new_n206), .o1(new_n211));
  norb02aa1n03x5               g116(.a(new_n206), .b(new_n205), .out0(new_n212));
  aoai13aa1n03x5               g117(.a(new_n212), .b(new_n197), .c(new_n189), .d(new_n200), .o1(new_n213));
  nona22aa1n03x5               g118(.a(new_n213), .b(new_n210), .c(new_n205), .out0(new_n214));
  nanp02aa1n03x5               g119(.a(new_n211), .b(new_n214), .o1(\s[20] ));
  aoi012aa1n12x5               g120(.a(new_n207), .b(new_n205), .c(new_n208), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  nano23aa1n06x5               g122(.a(new_n205), .b(new_n207), .c(new_n208), .d(new_n206), .out0(new_n218));
  aoi012aa1n06x5               g123(.a(new_n217), .b(new_n218), .c(new_n197), .o1(new_n219));
  nand02aa1d06x5               g124(.a(new_n200), .b(new_n218), .o1(new_n220));
  aoai13aa1n06x5               g125(.a(new_n219), .b(new_n220), .c(new_n185), .d(new_n178), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nand02aa1d24x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  nor002aa1n20x5               g130(.a(\b[21] ), .b(\a[22] ), .o1(new_n226));
  nand02aa1d28x5               g131(.a(\b[21] ), .b(\a[22] ), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n227), .b(new_n226), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n229), .b(new_n223), .c(new_n221), .d(new_n225), .o1(new_n230));
  inv030aa1n03x5               g135(.a(new_n219), .o1(new_n231));
  inv000aa1n02x5               g136(.a(new_n220), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n225), .b(new_n231), .c(new_n189), .d(new_n232), .o1(new_n233));
  nona22aa1n03x5               g138(.a(new_n233), .b(new_n229), .c(new_n223), .out0(new_n234));
  nanp02aa1n03x5               g139(.a(new_n230), .b(new_n234), .o1(\s[22] ));
  aoi012aa1n06x5               g140(.a(new_n226), .b(new_n223), .c(new_n227), .o1(new_n236));
  inv020aa1n03x5               g141(.a(new_n236), .o1(new_n237));
  nano23aa1d15x5               g142(.a(new_n223), .b(new_n226), .c(new_n227), .d(new_n224), .out0(new_n238));
  aoi012aa1d18x5               g143(.a(new_n237), .b(new_n231), .c(new_n238), .o1(new_n239));
  nano22aa1n06x5               g144(.a(new_n201), .b(new_n218), .c(new_n238), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n239), .b(new_n241), .c(new_n185), .d(new_n178), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  nand22aa1n09x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  norp02aa1n09x5               g151(.a(\b[23] ), .b(\a[24] ), .o1(new_n247));
  nand22aa1n12x5               g152(.a(\b[23] ), .b(\a[24] ), .o1(new_n248));
  nanb02aa1n02x5               g153(.a(new_n247), .b(new_n248), .out0(new_n249));
  aoai13aa1n02x5               g154(.a(new_n249), .b(new_n244), .c(new_n242), .d(new_n246), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n239), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n246), .b(new_n251), .c(new_n189), .d(new_n240), .o1(new_n252));
  nona22aa1n03x5               g157(.a(new_n252), .b(new_n249), .c(new_n244), .out0(new_n253));
  nanp02aa1n03x5               g158(.a(new_n250), .b(new_n253), .o1(\s[24] ));
  nanp03aa1n06x5               g159(.a(new_n197), .b(new_n212), .c(new_n209), .o1(new_n255));
  tech160nm_fiao0012aa1n02p5x5 g160(.a(new_n247), .b(new_n244), .c(new_n248), .o(new_n256));
  nano23aa1n09x5               g161(.a(new_n244), .b(new_n247), .c(new_n248), .d(new_n245), .out0(new_n257));
  tech160nm_fiaoi012aa1n05x5   g162(.a(new_n256), .b(new_n257), .c(new_n237), .o1(new_n258));
  nand22aa1n03x5               g163(.a(new_n257), .b(new_n238), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n258), .b(new_n259), .c(new_n255), .d(new_n216), .o1(new_n260));
  inv030aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  nano32aa1n02x4               g166(.a(new_n201), .b(new_n257), .c(new_n218), .d(new_n238), .out0(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n04x5               g168(.a(new_n261), .b(new_n263), .c(new_n185), .d(new_n178), .o1(new_n264));
  xorb03aa1n02x5               g169(.a(new_n264), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor002aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  xorc02aa1n12x5               g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  tech160nm_fixnrc02aa1n04x5   g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  aoai13aa1n02x5               g173(.a(new_n268), .b(new_n266), .c(new_n264), .d(new_n267), .o1(new_n269));
  aoai13aa1n03x5               g174(.a(new_n267), .b(new_n260), .c(new_n189), .d(new_n262), .o1(new_n270));
  nona22aa1n03x5               g175(.a(new_n270), .b(new_n268), .c(new_n266), .out0(new_n271));
  nanp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[26] ));
  inv000aa1d42x5               g177(.a(\a[26] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\b[25] ), .o1(new_n274));
  oaoi03aa1n02x5               g179(.a(new_n273), .b(new_n274), .c(new_n266), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  norb02aa1n02x5               g181(.a(new_n267), .b(new_n268), .out0(new_n277));
  aoi012aa1n06x5               g182(.a(new_n276), .b(new_n260), .c(new_n277), .o1(new_n278));
  nanb02aa1n02x5               g183(.a(new_n268), .b(new_n267), .out0(new_n279));
  nona22aa1n02x4               g184(.a(new_n232), .b(new_n259), .c(new_n279), .out0(new_n280));
  aoai13aa1n04x5               g185(.a(new_n278), .b(new_n280), .c(new_n185), .d(new_n178), .o1(new_n281));
  xorb03aa1n03x5               g186(.a(new_n281), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  xorc02aa1n12x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  xnrc02aa1n02x5               g189(.a(\b[27] ), .b(\a[28] ), .out0(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n283), .c(new_n281), .d(new_n284), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(new_n260), .b(new_n277), .o1(new_n287));
  nand22aa1n03x5               g192(.a(new_n287), .b(new_n275), .o1(new_n288));
  nano32aa1n03x7               g193(.a(new_n220), .b(new_n277), .c(new_n238), .d(new_n257), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n284), .b(new_n288), .c(new_n189), .d(new_n289), .o1(new_n290));
  nona22aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n283), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n286), .b(new_n291), .o1(\s[28] ));
  inv000aa1d42x5               g197(.a(\a[28] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  oaoi03aa1n09x5               g199(.a(new_n293), .b(new_n294), .c(new_n283), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  norb02aa1n02x5               g201(.a(new_n284), .b(new_n285), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n288), .c(new_n189), .d(new_n289), .o1(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .out0(new_n299));
  nona22aa1n03x5               g204(.a(new_n298), .b(new_n299), .c(new_n296), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n299), .b(new_n296), .c(new_n281), .d(new_n297), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n301), .b(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n119), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  tech160nm_fioaoi03aa1n03p5x5 g208(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .o1(new_n304));
  norb03aa1n02x5               g209(.a(new_n284), .b(new_n299), .c(new_n285), .out0(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n304), .c(new_n281), .d(new_n305), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n305), .b(new_n288), .c(new_n189), .d(new_n289), .o1(new_n308));
  nona22aa1n03x5               g213(.a(new_n308), .b(new_n306), .c(new_n304), .out0(new_n309));
  nanp02aa1n03x5               g214(.a(new_n307), .b(new_n309), .o1(\s[30] ));
  nanb02aa1n02x5               g215(.a(new_n306), .b(new_n304), .out0(new_n311));
  oai012aa1n02x5               g216(.a(new_n311), .b(\b[29] ), .c(\a[30] ), .o1(new_n312));
  norb02aa1n02x5               g217(.a(new_n305), .b(new_n306), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n288), .c(new_n189), .d(new_n289), .o1(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  nona22aa1n03x5               g220(.a(new_n314), .b(new_n315), .c(new_n312), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n315), .b(new_n312), .c(new_n281), .d(new_n313), .o1(new_n317));
  nanp02aa1n03x5               g222(.a(new_n317), .b(new_n316), .o1(\s[31] ));
  xnrb03aa1n02x5               g223(.a(new_n121), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g224(.a(\a[3] ), .b(\b[2] ), .c(new_n121), .o1(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g226(.a(new_n124), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n02x5               g227(.a(new_n125), .b(new_n102), .c(new_n124), .d(new_n126), .o1(new_n323));
  and002aa1n02x5               g228(.a(\b[5] ), .b(\a[6] ), .o(new_n324));
  nanb02aa1n02x5               g229(.a(new_n127), .b(new_n124), .out0(new_n325));
  nona32aa1n03x5               g230(.a(new_n325), .b(new_n324), .c(new_n102), .d(new_n101), .out0(new_n326));
  nanp02aa1n02x5               g231(.a(new_n326), .b(new_n323), .o1(\s[6] ));
  nona23aa1n02x4               g232(.a(new_n326), .b(new_n107), .c(new_n98), .d(new_n324), .out0(new_n328));
  aoi022aa1n02x5               g233(.a(new_n326), .b(new_n103), .c(new_n99), .d(new_n107), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n328), .b(new_n329), .out0(\s[7] ));
  aoi013aa1n02x4               g235(.a(new_n98), .b(new_n326), .c(new_n107), .d(new_n103), .o1(new_n331));
  xnrb03aa1n03x5               g236(.a(new_n331), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g237(.a(new_n130), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


