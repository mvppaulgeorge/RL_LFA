// Benchmark "adder" written by ABC on Wed Jul 17 18:59:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n341, new_n343, new_n345, new_n347,
    new_n349, new_n351, new_n352, new_n353;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  nor002aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1n03x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aob012aa1n02x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  nor042aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n02x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor042aa1n03x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n06x4               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nand23aa1n03x5               g014(.a(new_n103), .b(new_n106), .c(new_n109), .o1(new_n110));
  tech160nm_fioai012aa1n03p5x5 g015(.a(new_n105), .b(new_n107), .c(new_n104), .o1(new_n111));
  norp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand22aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor002aa1n03x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n03x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  norp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand42aa1n03x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  norp02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nano23aa1n02x4               g025(.a(new_n117), .b(new_n119), .c(new_n120), .d(new_n118), .out0(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n116), .o1(new_n122));
  norb02aa1n06x4               g027(.a(new_n115), .b(new_n114), .out0(new_n123));
  oai022aa1n03x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  aoi022aa1n06x5               g029(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  tech160nm_fiao0012aa1n02p5x5 g030(.a(new_n112), .b(new_n114), .c(new_n113), .o(new_n126));
  aoi013aa1n09x5               g031(.a(new_n126), .b(new_n123), .c(new_n124), .d(new_n125), .o1(new_n127));
  aoai13aa1n12x5               g032(.a(new_n127), .b(new_n122), .c(new_n110), .d(new_n111), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  nand22aa1n03x5               g034(.a(new_n128), .b(new_n129), .o1(new_n130));
  xorc02aa1n12x5               g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  oai022aa1d18x5               g037(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nand02aa1n02x5               g039(.a(new_n130), .b(new_n134), .o1(new_n135));
  nand42aa1n03x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nor042aa1d18x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  tech160nm_fiaoi012aa1n04x5   g042(.a(new_n137), .b(\a[10] ), .c(\b[9] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n138), .b(new_n136), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n139), .b(new_n135), .out0(new_n140));
  norb02aa1n02x5               g045(.a(new_n136), .b(new_n137), .out0(new_n141));
  aoi022aa1n02x5               g046(.a(new_n130), .b(new_n134), .c(\b[9] ), .d(\a[10] ), .o1(new_n142));
  oa0012aa1n03x5               g047(.a(new_n140), .b(new_n142), .c(new_n141), .o(\s[11] ));
  inv000aa1d42x5               g048(.a(new_n137), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n139), .c(new_n130), .d(new_n134), .o1(new_n145));
  nor042aa1n03x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  aoib12aa1n02x5               g053(.a(new_n137), .b(new_n147), .c(new_n146), .out0(new_n149));
  aoi022aa1n02x5               g054(.a(new_n140), .b(new_n149), .c(new_n145), .d(new_n148), .o1(\s[12] ));
  aoi012aa1n02x5               g055(.a(new_n99), .b(new_n101), .c(new_n102), .o1(new_n151));
  nona23aa1n09x5               g056(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n152));
  tech160nm_fioai012aa1n04x5   g057(.a(new_n111), .b(new_n152), .c(new_n151), .o1(new_n153));
  nanb02aa1n06x5               g058(.a(new_n122), .b(new_n153), .out0(new_n154));
  nano23aa1n09x5               g059(.a(new_n146), .b(new_n137), .c(new_n147), .d(new_n136), .out0(new_n155));
  nand23aa1n09x5               g060(.a(new_n155), .b(new_n129), .c(new_n131), .o1(new_n156));
  aoi022aa1n02x5               g061(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n157));
  nand03aa1n02x5               g062(.a(new_n138), .b(new_n133), .c(new_n157), .o1(new_n158));
  tech160nm_fiaoi012aa1n05x5   g063(.a(new_n146), .b(new_n137), .c(new_n147), .o1(new_n159));
  nanp02aa1n12x5               g064(.a(new_n158), .b(new_n159), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n02x7               g066(.a(new_n161), .b(new_n156), .c(new_n154), .d(new_n127), .o1(new_n162));
  nor042aa1n03x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  inv000aa1d42x5               g070(.a(new_n156), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n165), .b(new_n160), .c(new_n128), .d(new_n166), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n162), .c(new_n165), .o1(\s[13] ));
  nor042aa1n02x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand42aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  aoai13aa1n02x7               g076(.a(new_n171), .b(new_n163), .c(new_n162), .d(new_n164), .o1(new_n172));
  aoi112aa1n02x5               g077(.a(new_n163), .b(new_n171), .c(new_n162), .d(new_n165), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(\s[14] ));
  nano23aa1n06x5               g079(.a(new_n163), .b(new_n169), .c(new_n170), .d(new_n164), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n160), .c(new_n128), .d(new_n166), .o1(new_n176));
  tech160nm_fiaoi012aa1n04x5   g081(.a(new_n169), .b(new_n163), .c(new_n170), .o1(new_n177));
  nor042aa1n09x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nand42aa1n03x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  norb02aa1n09x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n176), .c(new_n177), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(new_n177), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n180), .b(new_n182), .c(new_n162), .d(new_n175), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n178), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n180), .o1(new_n185));
  aoai13aa1n03x5               g090(.a(new_n184), .b(new_n185), .c(new_n176), .d(new_n177), .o1(new_n186));
  nor002aa1n04x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nand42aa1n03x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  norb02aa1n02x5               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  aoib12aa1n02x5               g094(.a(new_n178), .b(new_n188), .c(new_n187), .out0(new_n190));
  aoi022aa1n02x5               g095(.a(new_n186), .b(new_n189), .c(new_n183), .d(new_n190), .o1(\s[16] ));
  nona23aa1n02x4               g096(.a(new_n170), .b(new_n164), .c(new_n163), .d(new_n169), .out0(new_n192));
  nano22aa1n03x7               g097(.a(new_n192), .b(new_n180), .c(new_n189), .out0(new_n193));
  nanb02aa1n03x5               g098(.a(new_n156), .b(new_n193), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n179), .b(new_n169), .c(new_n163), .d(new_n170), .o1(new_n195));
  aoi022aa1n02x5               g100(.a(new_n195), .b(new_n184), .c(\a[16] ), .d(\b[15] ), .o1(new_n196));
  aoi112aa1n06x5               g101(.a(new_n196), .b(new_n187), .c(new_n193), .d(new_n160), .o1(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n194), .c(new_n154), .d(new_n127), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g104(.a(\a[17] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(\b[16] ), .b(new_n200), .out0(new_n201));
  nano32aa1n03x7               g106(.a(new_n156), .b(new_n189), .c(new_n175), .d(new_n180), .out0(new_n202));
  nand42aa1n04x5               g107(.a(new_n193), .b(new_n160), .o1(new_n203));
  nona22aa1n09x5               g108(.a(new_n203), .b(new_n196), .c(new_n187), .out0(new_n204));
  xorc02aa1n02x5               g109(.a(\a[17] ), .b(\b[16] ), .out0(new_n205));
  aoai13aa1n02x5               g110(.a(new_n205), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n206));
  nor042aa1d18x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nand22aa1n12x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  norb02aa1n03x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n206), .c(new_n201), .out0(\s[18] ));
  and002aa1n02x5               g115(.a(new_n205), .b(new_n209), .o(new_n211));
  aoai13aa1n04x5               g116(.a(new_n211), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n212));
  nor042aa1n06x5               g117(.a(\b[16] ), .b(\a[17] ), .o1(new_n213));
  aoi012aa1n09x5               g118(.a(new_n207), .b(new_n213), .c(new_n208), .o1(new_n214));
  nor042aa1d18x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand02aa1n10x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g124(.a(new_n214), .o1(new_n220));
  aoai13aa1n04x5               g125(.a(new_n217), .b(new_n220), .c(new_n198), .d(new_n211), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n215), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n216), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n222), .b(new_n223), .c(new_n212), .d(new_n214), .o1(new_n224));
  nor042aa1n02x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand42aa1n03x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  norp02aa1n02x5               g132(.a(new_n227), .b(new_n215), .o1(new_n228));
  aoi022aa1n02x5               g133(.a(new_n224), .b(new_n227), .c(new_n221), .d(new_n228), .o1(\s[20] ));
  nano23aa1n02x5               g134(.a(new_n215), .b(new_n225), .c(new_n226), .d(new_n216), .out0(new_n230));
  and003aa1n02x5               g135(.a(new_n230), .b(new_n209), .c(new_n205), .o(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n232));
  nand02aa1n04x5               g137(.a(new_n213), .b(new_n208), .o1(new_n233));
  nona22aa1n09x5               g138(.a(new_n233), .b(new_n215), .c(new_n207), .out0(new_n234));
  aoai13aa1n12x5               g139(.a(new_n226), .b(new_n225), .c(new_n234), .d(new_n216), .o1(new_n235));
  nor042aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nand42aa1n03x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  xnbna2aa1n03x5               g143(.a(new_n238), .b(new_n232), .c(new_n235), .out0(\s[21] ));
  inv000aa1d42x5               g144(.a(new_n235), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n238), .b(new_n240), .c(new_n198), .d(new_n231), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n236), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n238), .o1(new_n243));
  aoai13aa1n02x5               g148(.a(new_n242), .b(new_n243), .c(new_n232), .d(new_n235), .o1(new_n244));
  norp02aa1n04x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  tech160nm_finand02aa1n05x5   g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  norb02aa1n02x5               g151(.a(new_n246), .b(new_n245), .out0(new_n247));
  aoib12aa1n02x5               g152(.a(new_n236), .b(new_n246), .c(new_n245), .out0(new_n248));
  aoi022aa1n03x5               g153(.a(new_n244), .b(new_n247), .c(new_n241), .d(new_n248), .o1(\s[22] ));
  nona23aa1n06x5               g154(.a(new_n246), .b(new_n237), .c(new_n236), .d(new_n245), .out0(new_n250));
  nano32aa1n02x4               g155(.a(new_n250), .b(new_n230), .c(new_n209), .d(new_n205), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n252));
  tech160nm_fiaoi012aa1n05x5   g157(.a(new_n245), .b(new_n236), .c(new_n246), .o1(new_n253));
  oa0012aa1n06x5               g158(.a(new_n253), .b(new_n235), .c(new_n250), .o(new_n254));
  nanp02aa1n02x5               g159(.a(new_n252), .b(new_n254), .o1(new_n255));
  nor042aa1d18x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  nand42aa1n08x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  norb02aa1n06x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  oai112aa1n02x5               g164(.a(new_n253), .b(new_n259), .c(new_n235), .d(new_n250), .o1(new_n260));
  aboi22aa1n03x5               g165(.a(new_n260), .b(new_n252), .c(new_n255), .d(new_n258), .out0(\s[23] ));
  inv040aa1d30x5               g166(.a(new_n254), .o1(new_n262));
  aoai13aa1n02x5               g167(.a(new_n258), .b(new_n262), .c(new_n198), .d(new_n251), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n256), .o1(new_n264));
  aoai13aa1n02x5               g169(.a(new_n264), .b(new_n259), .c(new_n252), .d(new_n254), .o1(new_n265));
  nor002aa1n02x5               g170(.a(\b[23] ), .b(\a[24] ), .o1(new_n266));
  nand42aa1n03x5               g171(.a(\b[23] ), .b(\a[24] ), .o1(new_n267));
  norb02aa1n06x4               g172(.a(new_n267), .b(new_n266), .out0(new_n268));
  aoib12aa1n02x5               g173(.a(new_n256), .b(new_n267), .c(new_n266), .out0(new_n269));
  aoi022aa1n02x5               g174(.a(new_n265), .b(new_n268), .c(new_n263), .d(new_n269), .o1(\s[24] ));
  nano23aa1n02x5               g175(.a(new_n236), .b(new_n245), .c(new_n246), .d(new_n237), .out0(new_n271));
  nanp03aa1n06x5               g176(.a(new_n271), .b(new_n258), .c(new_n268), .o1(new_n272));
  nano32aa1n02x5               g177(.a(new_n272), .b(new_n230), .c(new_n209), .d(new_n205), .out0(new_n273));
  aoai13aa1n04x5               g178(.a(new_n273), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n274));
  nand22aa1n03x5               g179(.a(new_n253), .b(new_n264), .o1(new_n275));
  aoai13aa1n12x5               g180(.a(new_n267), .b(new_n266), .c(new_n275), .d(new_n257), .o1(new_n276));
  oai012aa1d24x5               g181(.a(new_n276), .b(new_n235), .c(new_n272), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  nanp02aa1n02x5               g183(.a(new_n274), .b(new_n278), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[25] ), .b(\b[24] ), .out0(new_n280));
  oaoi03aa1n02x5               g185(.a(\a[19] ), .b(\b[18] ), .c(new_n214), .o1(new_n281));
  nano22aa1n03x7               g186(.a(new_n250), .b(new_n258), .c(new_n268), .out0(new_n282));
  oai112aa1n02x5               g187(.a(new_n282), .b(new_n226), .c(new_n281), .d(new_n225), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n280), .o1(new_n284));
  and003aa1n02x5               g189(.a(new_n283), .b(new_n284), .c(new_n276), .o(new_n285));
  aoi022aa1n02x5               g190(.a(new_n279), .b(new_n280), .c(new_n274), .d(new_n285), .o1(\s[25] ));
  aoai13aa1n03x5               g191(.a(new_n280), .b(new_n277), .c(new_n198), .d(new_n273), .o1(new_n287));
  norp02aa1n02x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n284), .c(new_n274), .d(new_n278), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[26] ), .b(\b[25] ), .out0(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n288), .o1(new_n292));
  aoi022aa1n02x5               g197(.a(new_n290), .b(new_n291), .c(new_n287), .d(new_n292), .o1(\s[26] ));
  nand02aa1n03x5               g198(.a(new_n291), .b(new_n280), .o1(new_n294));
  nano32aa1n03x7               g199(.a(new_n294), .b(new_n211), .c(new_n282), .d(new_n230), .out0(new_n295));
  aoai13aa1n04x5               g200(.a(new_n295), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n296));
  nanp02aa1n02x5               g201(.a(\b[25] ), .b(\a[26] ), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n294), .o1(new_n298));
  oai022aa1n02x5               g203(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n299));
  aoi022aa1d18x5               g204(.a(new_n277), .b(new_n298), .c(new_n297), .d(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  xnbna2aa1n06x5               g206(.a(new_n301), .b(new_n296), .c(new_n300), .out0(\s[27] ));
  nanp02aa1n02x5               g207(.a(new_n299), .b(new_n297), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n294), .c(new_n283), .d(new_n276), .o1(new_n304));
  aoai13aa1n02x5               g209(.a(new_n301), .b(new_n304), .c(new_n198), .d(new_n295), .o1(new_n305));
  norp02aa1n02x5               g210(.a(\b[26] ), .b(\a[27] ), .o1(new_n306));
  inv000aa1n03x5               g211(.a(new_n306), .o1(new_n307));
  inv000aa1n02x5               g212(.a(new_n301), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n307), .b(new_n308), .c(new_n296), .d(new_n300), .o1(new_n309));
  tech160nm_fixorc02aa1n03p5x5 g214(.a(\a[28] ), .b(\b[27] ), .out0(new_n310));
  norp02aa1n02x5               g215(.a(new_n310), .b(new_n306), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n305), .d(new_n311), .o1(\s[28] ));
  and002aa1n02x5               g217(.a(new_n310), .b(new_n301), .o(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n304), .c(new_n198), .d(new_n295), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .c(new_n307), .carry(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n296), .d(new_n300), .o1(new_n317));
  tech160nm_fixorc02aa1n02p5x5 g222(.a(\a[29] ), .b(\b[28] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n316), .b(new_n318), .out0(new_n319));
  aoi022aa1n03x5               g224(.a(new_n317), .b(new_n318), .c(new_n314), .d(new_n319), .o1(\s[29] ));
  xorb03aa1n02x5               g225(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g226(.a(new_n308), .b(new_n310), .c(new_n318), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n304), .c(new_n198), .d(new_n295), .o1(new_n323));
  inv000aa1d42x5               g228(.a(new_n322), .o1(new_n324));
  oaoi03aa1n02x5               g229(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .o1(new_n325));
  inv000aa1n03x5               g230(.a(new_n325), .o1(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n324), .c(new_n296), .d(new_n300), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .out0(new_n328));
  and002aa1n02x5               g233(.a(\b[28] ), .b(\a[29] ), .o(new_n329));
  oabi12aa1n02x5               g234(.a(new_n328), .b(\a[29] ), .c(\b[28] ), .out0(new_n330));
  oab012aa1n02x4               g235(.a(new_n330), .b(new_n316), .c(new_n329), .out0(new_n331));
  aoi022aa1n03x5               g236(.a(new_n327), .b(new_n328), .c(new_n323), .d(new_n331), .o1(\s[30] ));
  nano32aa1n06x5               g237(.a(new_n308), .b(new_n328), .c(new_n310), .d(new_n318), .out0(new_n333));
  aoai13aa1n03x5               g238(.a(new_n333), .b(new_n304), .c(new_n198), .d(new_n295), .o1(new_n334));
  xorc02aa1n02x5               g239(.a(\a[31] ), .b(\b[30] ), .out0(new_n335));
  oao003aa1n02x5               g240(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n336));
  norb02aa1n02x5               g241(.a(new_n336), .b(new_n335), .out0(new_n337));
  inv000aa1d42x5               g242(.a(new_n333), .o1(new_n338));
  aoai13aa1n03x5               g243(.a(new_n336), .b(new_n338), .c(new_n296), .d(new_n300), .o1(new_n339));
  aoi022aa1n03x5               g244(.a(new_n339), .b(new_n335), .c(new_n334), .d(new_n337), .o1(\s[31] ));
  aoi112aa1n02x5               g245(.a(new_n109), .b(new_n99), .c(new_n101), .d(new_n102), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n341), .b(new_n103), .c(new_n109), .o1(\s[3] ));
  aoi112aa1n02x5               g247(.a(new_n107), .b(new_n106), .c(new_n103), .d(new_n108), .o1(new_n343));
  aoib12aa1n02x5               g248(.a(new_n343), .b(new_n153), .c(new_n104), .out0(\s[4] ));
  norb02aa1n02x5               g249(.a(new_n120), .b(new_n119), .out0(new_n345));
  xnbna2aa1n03x5               g250(.a(new_n345), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  aoi012aa1n02x5               g251(.a(new_n119), .b(new_n153), .c(new_n120), .o1(new_n347));
  xnrb03aa1n02x5               g252(.a(new_n347), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g253(.a(new_n124), .b(new_n153), .c(new_n345), .o(new_n349));
  xobna2aa1n03x5               g254(.a(new_n123), .b(new_n349), .c(new_n118), .out0(\s[7] ));
  norb02aa1n02x5               g255(.a(new_n113), .b(new_n112), .out0(new_n351));
  aoi013aa1n02x4               g256(.a(new_n114), .b(new_n349), .c(new_n118), .d(new_n115), .o1(new_n352));
  aoi113aa1n02x5               g257(.a(new_n114), .b(new_n351), .c(new_n349), .d(new_n118), .e(new_n123), .o1(new_n353));
  aoib12aa1n02x5               g258(.a(new_n353), .b(new_n351), .c(new_n352), .out0(\s[8] ));
  xnbna2aa1n03x5               g259(.a(new_n129), .b(new_n154), .c(new_n127), .out0(\s[9] ));
endmodule


