// Benchmark "adder" written by ABC on Thu Jul 18 11:19:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n337, new_n339, new_n340,
    new_n342, new_n343, new_n345, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  and002aa1n06x5               g002(.a(\b[0] ), .b(\a[1] ), .o(new_n98));
  oaoi03aa1n12x5               g003(.a(\a[2] ), .b(\b[1] ), .c(new_n98), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nand42aa1n06x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nano23aa1n09x5               g008(.a(new_n100), .b(new_n102), .c(new_n103), .d(new_n101), .out0(new_n104));
  tech160nm_fiao0012aa1n05x5   g009(.a(new_n100), .b(new_n102), .c(new_n101), .o(new_n105));
  aoi012aa1n02x5               g010(.a(new_n105), .b(new_n104), .c(new_n99), .o1(new_n106));
  norp02aa1n12x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand42aa1n08x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nor042aa1d18x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nand42aa1n03x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nano23aa1n06x5               g015(.a(new_n107), .b(new_n109), .c(new_n110), .d(new_n108), .out0(new_n111));
  nand42aa1n03x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor042aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  norb02aa1n06x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  xorc02aa1n02x5               g019(.a(\a[8] ), .b(\b[7] ), .out0(new_n115));
  nand23aa1n03x5               g020(.a(new_n111), .b(new_n114), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[8] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\b[7] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(new_n107), .o1(new_n119));
  aoai13aa1n06x5               g024(.a(new_n108), .b(new_n113), .c(new_n109), .d(new_n112), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(new_n117), .b(new_n118), .c(new_n121), .o1(new_n122));
  oai012aa1n06x5               g027(.a(new_n122), .b(new_n106), .c(new_n116), .o1(new_n123));
  nand42aa1n10x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  aoi012aa1n02x5               g029(.a(new_n97), .b(new_n123), .c(new_n124), .o1(new_n125));
  xnrb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1d28x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nanp02aa1n12x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(\a[11] ), .o1(new_n129));
  nanb02aa1d36x5               g034(.a(\b[10] ), .b(new_n129), .out0(new_n130));
  nand02aa1d06x5               g035(.a(new_n130), .b(new_n128), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n124), .b(new_n97), .out0(new_n132));
  nor042aa1n09x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norp02aa1n02x5               g038(.a(new_n97), .b(new_n133), .o1(new_n134));
  aob012aa1n02x5               g039(.a(new_n134), .b(new_n123), .c(new_n132), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n131), .b(new_n135), .c(new_n127), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n130), .o1(new_n137));
  nano22aa1n02x4               g042(.a(new_n137), .b(new_n127), .c(new_n128), .out0(new_n138));
  tech160nm_fixnrc02aa1n04x5   g043(.a(\b[11] ), .b(\a[12] ), .out0(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n137), .c(new_n135), .d(new_n138), .o1(new_n140));
  aoi112aa1n02x7               g045(.a(new_n139), .b(new_n137), .c(new_n135), .d(new_n138), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(\s[12] ));
  nand02aa1n03x5               g047(.a(new_n104), .b(new_n99), .o1(new_n143));
  inv040aa1n02x5               g048(.a(new_n105), .o1(new_n144));
  nand42aa1n02x5               g049(.a(new_n143), .b(new_n144), .o1(new_n145));
  inv030aa1n02x5               g050(.a(new_n116), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(new_n118), .b(new_n117), .o1(new_n147));
  and002aa1n02x5               g052(.a(\b[7] ), .b(\a[8] ), .o(new_n148));
  aoai13aa1n06x5               g053(.a(new_n147), .b(new_n148), .c(new_n120), .d(new_n119), .o1(new_n149));
  nano23aa1d15x5               g054(.a(new_n133), .b(new_n97), .c(new_n124), .d(new_n127), .out0(new_n150));
  nona22aa1d36x5               g055(.a(new_n150), .b(new_n139), .c(new_n131), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n03x5               g057(.a(new_n152), .b(new_n149), .c(new_n146), .d(new_n145), .o1(new_n153));
  inv000aa1d42x5               g058(.a(\a[12] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(\b[11] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n155), .b(new_n154), .o1(new_n156));
  and002aa1n02x5               g061(.a(\b[11] ), .b(\a[12] ), .o(new_n157));
  aoai13aa1n12x5               g062(.a(new_n128), .b(new_n133), .c(new_n97), .d(new_n127), .o1(new_n158));
  aoai13aa1n12x5               g063(.a(new_n156), .b(new_n157), .c(new_n158), .d(new_n130), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nor002aa1d32x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nand02aa1d04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(new_n161), .b(new_n162), .out0(new_n163));
  xobna2aa1n03x5               g068(.a(new_n163), .b(new_n153), .c(new_n160), .out0(\s[13] ));
  inv000aa1d42x5               g069(.a(new_n161), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n163), .c(new_n153), .d(new_n160), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand02aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nona23aa1d18x5               g074(.a(new_n169), .b(new_n162), .c(new_n161), .d(new_n168), .out0(new_n170));
  inv040aa1n02x5               g075(.a(new_n170), .o1(new_n171));
  aoai13aa1n02x5               g076(.a(new_n171), .b(new_n159), .c(new_n123), .d(new_n152), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n168), .b(new_n161), .c(new_n169), .o1(new_n173));
  nor022aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nand42aa1n08x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nanb02aa1n12x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n172), .c(new_n173), .out0(\s[15] ));
  aoai13aa1n06x5               g083(.a(new_n173), .b(new_n170), .c(new_n153), .d(new_n160), .o1(new_n179));
  nor002aa1n02x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nand42aa1n03x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n174), .c(new_n179), .d(new_n175), .o1(new_n183));
  nand42aa1n03x5               g088(.a(new_n179), .b(new_n177), .o1(new_n184));
  nona22aa1n02x4               g089(.a(new_n184), .b(new_n182), .c(new_n174), .out0(new_n185));
  nanp02aa1n02x5               g090(.a(new_n185), .b(new_n183), .o1(\s[16] ));
  nano23aa1n02x5               g091(.a(new_n174), .b(new_n180), .c(new_n181), .d(new_n175), .out0(new_n187));
  nano22aa1n12x5               g092(.a(new_n151), .b(new_n171), .c(new_n187), .out0(new_n188));
  aoai13aa1n12x5               g093(.a(new_n188), .b(new_n149), .c(new_n146), .d(new_n145), .o1(new_n189));
  norp03aa1n09x5               g094(.a(new_n170), .b(new_n176), .c(new_n182), .o1(new_n190));
  aoai13aa1n06x5               g095(.a(new_n175), .b(new_n168), .c(new_n161), .d(new_n169), .o1(new_n191));
  tech160nm_fioai012aa1n03p5x5 g096(.a(new_n191), .b(\b[14] ), .c(\a[15] ), .o1(new_n192));
  tech160nm_fiao0012aa1n02p5x5 g097(.a(new_n180), .b(new_n192), .c(new_n181), .o(new_n193));
  aoi012aa1d18x5               g098(.a(new_n193), .b(new_n159), .c(new_n190), .o1(new_n194));
  nand02aa1d08x5               g099(.a(new_n189), .b(new_n194), .o1(new_n195));
  nor042aa1n09x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nand42aa1n20x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  aoi112aa1n02x5               g103(.a(new_n193), .b(new_n198), .c(new_n159), .d(new_n190), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n195), .b(new_n198), .c(new_n199), .d(new_n189), .o1(\s[17] ));
  inv000aa1d42x5               g105(.a(\a[18] ), .o1(new_n201));
  tech160nm_fiaoi012aa1n05x5   g106(.a(new_n196), .b(new_n195), .c(new_n198), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[17] ), .c(new_n201), .out0(\s[18] ));
  nor042aa1n06x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nand42aa1n20x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nano23aa1d15x5               g110(.a(new_n196), .b(new_n204), .c(new_n205), .d(new_n197), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  oa0012aa1n02x5               g112(.a(new_n205), .b(new_n204), .c(new_n196), .o(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n207), .c(new_n189), .d(new_n194), .o1(new_n210));
  nor042aa1n04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand42aa1n03x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n09x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  aoi112aa1n03x4               g118(.a(new_n213), .b(new_n208), .c(new_n195), .d(new_n206), .o1(new_n214));
  aoi012aa1n02x5               g119(.a(new_n214), .b(new_n210), .c(new_n213), .o1(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1n06x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n06x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n211), .c(new_n210), .d(new_n212), .o1(new_n220));
  nand02aa1d04x5               g125(.a(new_n210), .b(new_n213), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n219), .c(new_n211), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n222), .b(new_n220), .o1(\s[20] ));
  nanb03aa1d24x5               g128(.a(new_n219), .b(new_n206), .c(new_n213), .out0(new_n224));
  nanb03aa1n12x5               g129(.a(new_n217), .b(new_n218), .c(new_n212), .out0(new_n225));
  orn002aa1n02x5               g130(.a(\a[19] ), .b(\b[18] ), .o(new_n226));
  oai112aa1n06x5               g131(.a(new_n226), .b(new_n205), .c(new_n204), .d(new_n196), .o1(new_n227));
  aoi012aa1d24x5               g132(.a(new_n217), .b(new_n211), .c(new_n218), .o1(new_n228));
  oai012aa1d24x5               g133(.a(new_n228), .b(new_n227), .c(new_n225), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n224), .c(new_n189), .d(new_n194), .o1(new_n231));
  nor042aa1n03x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n224), .o1(new_n235));
  aoi112aa1n03x4               g140(.a(new_n234), .b(new_n229), .c(new_n195), .d(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n231), .c(new_n234), .o1(\s[21] ));
  nor042aa1n02x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nanp02aa1n04x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n238), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n241), .b(new_n232), .c(new_n231), .d(new_n234), .o1(new_n242));
  nand42aa1n04x5               g147(.a(new_n231), .b(new_n234), .o1(new_n243));
  nona22aa1n02x4               g148(.a(new_n243), .b(new_n241), .c(new_n232), .out0(new_n244));
  nanp02aa1n03x5               g149(.a(new_n244), .b(new_n242), .o1(\s[22] ));
  nano23aa1n06x5               g150(.a(new_n232), .b(new_n238), .c(new_n239), .d(new_n233), .out0(new_n246));
  nanp03aa1n02x5               g151(.a(new_n195), .b(new_n235), .c(new_n246), .o1(new_n247));
  nona23aa1n02x4               g152(.a(new_n246), .b(new_n213), .c(new_n207), .d(new_n219), .out0(new_n248));
  nano22aa1n02x4               g153(.a(new_n217), .b(new_n212), .c(new_n218), .out0(new_n249));
  oai012aa1n02x5               g154(.a(new_n205), .b(\b[18] ), .c(\a[19] ), .o1(new_n250));
  oab012aa1n02x4               g155(.a(new_n250), .b(new_n196), .c(new_n204), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n228), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n246), .b(new_n252), .c(new_n251), .d(new_n249), .o1(new_n253));
  aoi012aa1d18x5               g158(.a(new_n238), .b(new_n232), .c(new_n239), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(new_n253), .b(new_n254), .o1(new_n255));
  inv000aa1n02x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n248), .c(new_n189), .d(new_n194), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[23] ), .b(\b[22] ), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n254), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(new_n258), .b(new_n259), .c(new_n229), .d(new_n246), .o1(new_n260));
  aoi022aa1n02x5               g165(.a(new_n247), .b(new_n260), .c(new_n257), .d(new_n258), .o1(\s[23] ));
  norp02aa1n02x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  xnrc02aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .out0(new_n263));
  aoai13aa1n03x5               g168(.a(new_n263), .b(new_n262), .c(new_n257), .d(new_n258), .o1(new_n264));
  nand42aa1n02x5               g169(.a(new_n257), .b(new_n258), .o1(new_n265));
  nona22aa1n03x5               g170(.a(new_n265), .b(new_n263), .c(new_n262), .out0(new_n266));
  nanp02aa1n03x5               g171(.a(new_n266), .b(new_n264), .o1(\s[24] ));
  norb02aa1n02x7               g172(.a(new_n258), .b(new_n263), .out0(new_n268));
  nanb03aa1n03x5               g173(.a(new_n224), .b(new_n268), .c(new_n246), .out0(new_n269));
  inv000aa1n02x5               g174(.a(new_n268), .o1(new_n270));
  orn002aa1n02x5               g175(.a(\a[23] ), .b(\b[22] ), .o(new_n271));
  oao003aa1n02x5               g176(.a(\a[24] ), .b(\b[23] ), .c(new_n271), .carry(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n270), .c(new_n253), .d(new_n254), .o1(new_n273));
  inv040aa1n03x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n269), .c(new_n189), .d(new_n194), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  tech160nm_fixnrc02aa1n05x5   g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  nand42aa1n02x5               g185(.a(new_n275), .b(new_n278), .o1(new_n281));
  nona22aa1n03x5               g186(.a(new_n281), .b(new_n279), .c(new_n277), .out0(new_n282));
  nanp02aa1n03x5               g187(.a(new_n282), .b(new_n280), .o1(\s[26] ));
  tech160nm_finand02aa1n03p5x5 g188(.a(new_n159), .b(new_n190), .o1(new_n284));
  aoi012aa1n02x5               g189(.a(new_n180), .b(new_n192), .c(new_n181), .o1(new_n285));
  nanp02aa1n03x5               g190(.a(new_n284), .b(new_n285), .o1(new_n286));
  norb02aa1n03x4               g191(.a(new_n278), .b(new_n279), .out0(new_n287));
  inv000aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nano23aa1d15x5               g193(.a(new_n288), .b(new_n224), .c(new_n268), .d(new_n246), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n286), .c(new_n123), .d(new_n188), .o1(new_n290));
  inv000aa1d42x5               g195(.a(\a[26] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\b[25] ), .o1(new_n292));
  tech160nm_fioaoi03aa1n03p5x5 g197(.a(new_n291), .b(new_n292), .c(new_n277), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  aoi012aa1n12x5               g199(.a(new_n294), .b(new_n273), .c(new_n287), .o1(new_n295));
  xorc02aa1n12x5               g200(.a(\a[27] ), .b(\b[26] ), .out0(new_n296));
  xnbna2aa1n03x5               g201(.a(new_n296), .b(new_n295), .c(new_n290), .out0(\s[27] ));
  xnrc02aa1n02x5               g202(.a(\b[27] ), .b(\a[28] ), .out0(new_n298));
  norp02aa1n02x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  inv000aa1n03x5               g204(.a(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n296), .o1(new_n301));
  aoai13aa1n04x5               g206(.a(new_n300), .b(new_n301), .c(new_n295), .d(new_n290), .o1(new_n302));
  nand02aa1n02x5               g207(.a(new_n302), .b(new_n298), .o1(new_n303));
  aoai13aa1n06x5               g208(.a(new_n268), .b(new_n259), .c(new_n229), .d(new_n246), .o1(new_n304));
  aoai13aa1n04x5               g209(.a(new_n293), .b(new_n288), .c(new_n304), .d(new_n272), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n296), .b(new_n305), .c(new_n195), .d(new_n289), .o1(new_n306));
  nona22aa1n03x5               g211(.a(new_n306), .b(new_n298), .c(new_n299), .out0(new_n307));
  nanp02aa1n03x5               g212(.a(new_n303), .b(new_n307), .o1(\s[28] ));
  norb02aa1n02x5               g213(.a(new_n296), .b(new_n298), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n195), .d(new_n289), .o1(new_n310));
  tech160nm_fixorc02aa1n02p5x5 g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  oao003aa1n02x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n300), .carry(new_n312));
  norb02aa1n02x5               g217(.a(new_n312), .b(new_n311), .out0(new_n313));
  inv000aa1n02x5               g218(.a(new_n309), .o1(new_n314));
  aoai13aa1n02x7               g219(.a(new_n312), .b(new_n314), .c(new_n295), .d(new_n290), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n310), .d(new_n313), .o1(\s[29] ));
  xnrb03aa1n02x5               g221(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g222(.a(new_n298), .b(new_n296), .c(new_n311), .out0(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n305), .c(new_n195), .d(new_n289), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .out0(new_n320));
  oao003aa1n03x5               g225(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .carry(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(new_n322));
  inv000aa1d42x5               g227(.a(new_n318), .o1(new_n323));
  aoai13aa1n02x7               g228(.a(new_n321), .b(new_n323), .c(new_n295), .d(new_n290), .o1(new_n324));
  aoi022aa1n03x5               g229(.a(new_n324), .b(new_n320), .c(new_n319), .d(new_n322), .o1(\s[30] ));
  nano22aa1n06x5               g230(.a(new_n314), .b(new_n311), .c(new_n320), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n305), .c(new_n195), .d(new_n289), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[31] ), .b(\b[30] ), .out0(new_n328));
  oao003aa1n02x5               g233(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n329));
  norb02aa1n02x5               g234(.a(new_n329), .b(new_n328), .out0(new_n330));
  inv000aa1d42x5               g235(.a(new_n326), .o1(new_n331));
  aoai13aa1n02x7               g236(.a(new_n329), .b(new_n331), .c(new_n295), .d(new_n290), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n332), .b(new_n328), .c(new_n327), .d(new_n330), .o1(\s[31] ));
  xorb03aa1n02x5               g238(.a(new_n99), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oai012aa1n02x5               g239(.a(new_n103), .b(new_n99), .c(new_n102), .o1(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  norb02aa1n02x5               g241(.a(new_n110), .b(new_n109), .out0(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n337), .b(new_n143), .c(new_n144), .out0(\s[5] ));
  inv000aa1d42x5               g243(.a(new_n109), .o1(new_n339));
  aoai13aa1n02x5               g244(.a(new_n337), .b(new_n105), .c(new_n104), .d(new_n99), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n114), .b(new_n340), .c(new_n339), .out0(\s[6] ));
  aobi12aa1n02x5               g246(.a(new_n114), .b(new_n340), .c(new_n339), .out0(new_n342));
  norp02aa1n02x5               g247(.a(new_n342), .b(new_n113), .o1(new_n343));
  xnrb03aa1n02x5               g248(.a(new_n343), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oai013aa1n02x4               g249(.a(new_n108), .b(new_n342), .c(new_n113), .d(new_n107), .o1(new_n345));
  xorb03aa1n02x5               g250(.a(new_n345), .b(\b[7] ), .c(new_n117), .out0(\s[8] ));
  aoi112aa1n02x5               g251(.a(new_n149), .b(new_n132), .c(new_n146), .d(new_n145), .o1(new_n347));
  aoi012aa1n02x5               g252(.a(new_n347), .b(new_n123), .c(new_n132), .o1(\s[9] ));
endmodule


