// Benchmark "adder" written by ABC on Thu Jul 18 00:51:55 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n337, new_n340,
    new_n342, new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n12x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand02aa1n03x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nona23aa1n09x5               g007(.a(new_n102), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n103));
  tech160nm_finor002aa1n03p5x5 g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nor022aa1n04x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nona23aa1n02x4               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  nor042aa1n03x5               g013(.a(new_n108), .b(new_n103), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[1] ), .b(\a[2] ), .o1(new_n110));
  nand22aa1n03x5               g015(.a(\b[0] ), .b(\a[1] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[1] ), .b(\a[2] ), .o1(new_n112));
  tech160nm_fiaoi012aa1n05x5   g017(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n113));
  inv040aa1d32x5               g018(.a(\a[4] ), .o1(new_n114));
  inv040aa1d32x5               g019(.a(\b[3] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(new_n115), .b(new_n114), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n116), .b(new_n117), .o1(new_n118));
  nor022aa1n16x5               g023(.a(\b[2] ), .b(\a[3] ), .o1(new_n119));
  nand42aa1n02x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  nanb02aa1n02x5               g025(.a(new_n119), .b(new_n120), .out0(new_n121));
  oaoi03aa1n12x5               g026(.a(new_n114), .b(new_n115), .c(new_n119), .o1(new_n122));
  oai013aa1n06x5               g027(.a(new_n122), .b(new_n113), .c(new_n121), .d(new_n118), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n99), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(new_n101), .b(new_n100), .o1(new_n125));
  oaih12aa1n02x5               g030(.a(new_n105), .b(new_n106), .c(new_n104), .o1(new_n126));
  oai112aa1n04x5               g031(.a(new_n124), .b(new_n125), .c(new_n103), .d(new_n126), .o1(new_n127));
  nanp02aa1n09x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n97), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n127), .c(new_n123), .d(new_n109), .o1(new_n130));
  nor042aa1n04x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nand42aa1n06x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n133), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  norp03aa1n02x5               g039(.a(new_n113), .b(new_n121), .c(new_n118), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n122), .o1(new_n136));
  tech160nm_fioai012aa1n05x5   g041(.a(new_n109), .b(new_n135), .c(new_n136), .o1(new_n137));
  norp02aa1n02x5               g042(.a(new_n103), .b(new_n126), .o1(new_n138));
  nano22aa1n02x5               g043(.a(new_n138), .b(new_n124), .c(new_n125), .out0(new_n139));
  nano23aa1d15x5               g044(.a(new_n97), .b(new_n131), .c(new_n132), .d(new_n128), .out0(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  tech160nm_fioai012aa1n05x5   g046(.a(new_n132), .b(new_n131), .c(new_n97), .o1(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n141), .c(new_n137), .d(new_n139), .o1(new_n143));
  xorb03aa1n02x5               g048(.a(new_n143), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  nanp02aa1n04x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  aoi012aa1n03x5               g051(.a(new_n145), .b(new_n143), .c(new_n146), .o1(new_n147));
  nor002aa1n16x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nanp02aa1n04x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n147), .b(new_n150), .c(new_n149), .out0(\s[12] ));
  nanp02aa1n02x5               g056(.a(new_n145), .b(new_n150), .o1(new_n152));
  nona23aa1d18x5               g057(.a(new_n150), .b(new_n146), .c(new_n145), .d(new_n148), .out0(new_n153));
  oai112aa1n06x5               g058(.a(new_n152), .b(new_n149), .c(new_n153), .d(new_n142), .o1(new_n154));
  aoi112aa1n03x5               g059(.a(new_n153), .b(new_n141), .c(new_n137), .d(new_n139), .o1(new_n155));
  nor042aa1d18x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand02aa1n03x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nanb02aa1n02x5               g062(.a(new_n156), .b(new_n157), .out0(new_n158));
  oabi12aa1n06x5               g063(.a(new_n158), .b(new_n155), .c(new_n154), .out0(new_n159));
  inv040aa1n03x5               g064(.a(new_n156), .o1(new_n160));
  aoi112aa1n02x5               g065(.a(new_n155), .b(new_n154), .c(new_n160), .d(new_n157), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n159), .b(new_n161), .out0(\s[13] ));
  nor042aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  xobna2aa1n03x5               g070(.a(new_n165), .b(new_n159), .c(new_n160), .out0(\s[14] ));
  nano23aa1n06x5               g071(.a(new_n156), .b(new_n163), .c(new_n164), .d(new_n157), .out0(new_n167));
  oaoi03aa1n02x7               g072(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n168), .b(new_n154), .c(new_n167), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(new_n137), .b(new_n139), .o1(new_n170));
  nona23aa1n02x4               g075(.a(new_n164), .b(new_n157), .c(new_n156), .d(new_n163), .out0(new_n171));
  nona32aa1n02x4               g076(.a(new_n170), .b(new_n171), .c(new_n153), .d(new_n141), .out0(new_n172));
  nor042aa1d18x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n16x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n172), .c(new_n169), .out0(\s[15] ));
  inv000aa1d42x5               g081(.a(new_n173), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n175), .o1(new_n178));
  aoai13aa1n02x5               g083(.a(new_n177), .b(new_n178), .c(new_n172), .d(new_n169), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nano23aa1n06x5               g085(.a(new_n145), .b(new_n148), .c(new_n150), .d(new_n146), .out0(new_n181));
  nor042aa1n04x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand42aa1n16x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nano23aa1d15x5               g088(.a(new_n173), .b(new_n182), .c(new_n183), .d(new_n174), .out0(new_n184));
  nand02aa1d04x5               g089(.a(new_n184), .b(new_n167), .o1(new_n185));
  nano22aa1n03x7               g090(.a(new_n185), .b(new_n140), .c(new_n181), .out0(new_n186));
  aoai13aa1n12x5               g091(.a(new_n186), .b(new_n127), .c(new_n123), .d(new_n109), .o1(new_n187));
  aoi122aa1n12x5               g092(.a(new_n182), .b(new_n183), .c(new_n173), .d(new_n184), .e(new_n168), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n184), .o1(new_n189));
  nona32aa1n09x5               g094(.a(new_n154), .b(new_n189), .c(new_n165), .d(new_n158), .out0(new_n190));
  nand23aa1d12x5               g095(.a(new_n187), .b(new_n188), .c(new_n190), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[16] ), .o1(new_n194));
  tech160nm_fioaoi03aa1n03p5x5 g099(.a(new_n193), .b(new_n194), .c(new_n191), .o1(new_n195));
  nor002aa1d32x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nand42aa1n08x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nanb02aa1n02x5               g102(.a(new_n196), .b(new_n197), .out0(new_n198));
  tech160nm_fixorc02aa1n02p5x5 g103(.a(new_n195), .b(new_n198), .out0(\s[18] ));
  inv000aa1n06x5               g104(.a(new_n188), .o1(new_n200));
  aoi013aa1n06x4               g105(.a(new_n200), .b(new_n154), .c(new_n167), .d(new_n184), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(new_n194), .b(new_n193), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  nano22aa1n12x5               g108(.a(new_n198), .b(new_n202), .c(new_n203), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  aoai13aa1n12x5               g110(.a(new_n197), .b(new_n196), .c(new_n193), .d(new_n194), .o1(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n205), .c(new_n201), .d(new_n187), .o1(new_n207));
  xorb03aa1n03x5               g112(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n16x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nand42aa1n02x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanb02aa1n12x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  inv000aa1d42x5               g118(.a(\b[19] ), .o1(new_n214));
  nanb02aa1n18x5               g119(.a(\a[20] ), .b(new_n214), .out0(new_n215));
  nanp02aa1n03x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand02aa1d06x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoi112aa1n03x5               g123(.a(new_n210), .b(new_n218), .c(new_n207), .d(new_n213), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n210), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n206), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n213), .b(new_n221), .c(new_n191), .d(new_n204), .o1(new_n222));
  aoi012aa1n03x5               g127(.a(new_n217), .b(new_n222), .c(new_n220), .o1(new_n223));
  norp02aa1n03x5               g128(.a(new_n223), .b(new_n219), .o1(\s[20] ));
  nona22aa1d24x5               g129(.a(new_n204), .b(new_n212), .c(new_n217), .out0(new_n225));
  nanp02aa1n02x5               g130(.a(new_n210), .b(new_n216), .o1(new_n226));
  nor043aa1n03x5               g131(.a(new_n206), .b(new_n212), .c(new_n217), .o1(new_n227));
  nano22aa1n02x4               g132(.a(new_n227), .b(new_n215), .c(new_n226), .out0(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n225), .c(new_n201), .d(new_n187), .o1(new_n229));
  xorb03aa1n02x5               g134(.a(new_n229), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  xorc02aa1n06x5               g136(.a(\a[21] ), .b(\b[20] ), .out0(new_n232));
  xorc02aa1n12x5               g137(.a(\a[22] ), .b(\b[21] ), .out0(new_n233));
  aoi112aa1n03x5               g138(.a(new_n231), .b(new_n233), .c(new_n229), .d(new_n232), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n231), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n225), .o1(new_n236));
  norp02aa1n02x5               g141(.a(\b[19] ), .b(\a[20] ), .o1(new_n237));
  nona23aa1n02x4               g142(.a(new_n216), .b(new_n211), .c(new_n210), .d(new_n237), .out0(new_n238));
  oai112aa1n06x5               g143(.a(new_n226), .b(new_n215), .c(new_n238), .d(new_n206), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n232), .b(new_n239), .c(new_n191), .d(new_n236), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n233), .o1(new_n241));
  tech160nm_fiaoi012aa1n02p5x5 g146(.a(new_n241), .b(new_n240), .c(new_n235), .o1(new_n242));
  nor002aa1n02x5               g147(.a(new_n242), .b(new_n234), .o1(\s[22] ));
  nano22aa1n03x7               g148(.a(new_n225), .b(new_n232), .c(new_n233), .out0(new_n244));
  inv020aa1n02x5               g149(.a(new_n244), .o1(new_n245));
  and002aa1n02x5               g150(.a(new_n233), .b(new_n232), .o(new_n246));
  tech160nm_fioaoi03aa1n03p5x5 g151(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .o1(new_n247));
  aoi012aa1n09x5               g152(.a(new_n247), .b(new_n239), .c(new_n246), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n245), .c(new_n201), .d(new_n187), .o1(new_n249));
  xorb03aa1n02x5               g154(.a(new_n249), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor022aa1n16x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  nand42aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  nor042aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(\b[23] ), .b(\a[24] ), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n255), .b(new_n254), .out0(new_n256));
  aoi112aa1n03x4               g161(.a(new_n251), .b(new_n256), .c(new_n249), .d(new_n253), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n251), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n248), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n253), .b(new_n259), .c(new_n191), .d(new_n244), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n256), .o1(new_n261));
  aoi012aa1n03x5               g166(.a(new_n261), .b(new_n260), .c(new_n258), .o1(new_n262));
  norp02aa1n03x5               g167(.a(new_n262), .b(new_n257), .o1(\s[24] ));
  nano23aa1n06x5               g168(.a(new_n251), .b(new_n254), .c(new_n255), .d(new_n252), .out0(new_n264));
  nano32aa1n03x7               g169(.a(new_n225), .b(new_n264), .c(new_n232), .d(new_n233), .out0(new_n265));
  inv000aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  aoi112aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n267));
  nand42aa1n04x5               g172(.a(new_n264), .b(new_n247), .o1(new_n268));
  nona22aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n254), .out0(new_n269));
  nand23aa1n06x5               g174(.a(new_n264), .b(new_n232), .c(new_n233), .o1(new_n270));
  inv040aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  aoi012aa1n09x5               g176(.a(new_n269), .b(new_n239), .c(new_n271), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n266), .c(new_n201), .d(new_n187), .o1(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  aoi112aa1n03x4               g182(.a(new_n275), .b(new_n277), .c(new_n273), .d(new_n276), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n275), .o1(new_n279));
  inv000aa1n02x5               g184(.a(new_n272), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n276), .b(new_n280), .c(new_n191), .d(new_n265), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n277), .o1(new_n282));
  tech160nm_fiaoi012aa1n02p5x5 g187(.a(new_n282), .b(new_n281), .c(new_n279), .o1(new_n283));
  nor002aa1n02x5               g188(.a(new_n283), .b(new_n278), .o1(\s[26] ));
  nona23aa1n02x4               g189(.a(new_n140), .b(new_n184), .c(new_n171), .d(new_n153), .out0(new_n285));
  tech160nm_fiaoi012aa1n05x5   g190(.a(new_n285), .b(new_n137), .c(new_n139), .o1(new_n286));
  nanp02aa1n06x5               g191(.a(new_n190), .b(new_n188), .o1(new_n287));
  and002aa1n02x5               g192(.a(new_n277), .b(new_n276), .o(new_n288));
  nano32aa1d12x5               g193(.a(new_n225), .b(new_n288), .c(new_n246), .d(new_n264), .out0(new_n289));
  oai012aa1n06x5               g194(.a(new_n289), .b(new_n287), .c(new_n286), .o1(new_n290));
  norp02aa1n02x5               g195(.a(\b[25] ), .b(\a[26] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoi112aa1n02x7               g197(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n293));
  inv000aa1n02x5               g198(.a(new_n293), .o1(new_n294));
  aoi112aa1n06x5               g199(.a(new_n267), .b(new_n254), .c(new_n264), .d(new_n247), .o1(new_n295));
  inv000aa1n02x5               g200(.a(new_n288), .o1(new_n296));
  oaoi13aa1n03x5               g201(.a(new_n296), .b(new_n295), .c(new_n228), .d(new_n270), .o1(new_n297));
  nano22aa1n03x7               g202(.a(new_n297), .b(new_n292), .c(new_n294), .out0(new_n298));
  xorc02aa1n02x5               g203(.a(\a[27] ), .b(\b[26] ), .out0(new_n299));
  xnbna2aa1n03x5               g204(.a(new_n299), .b(new_n290), .c(new_n298), .out0(\s[27] ));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  inv040aa1n03x5               g206(.a(new_n301), .o1(new_n302));
  aobi12aa1n02x5               g207(.a(new_n299), .b(new_n290), .c(new_n298), .out0(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[27] ), .b(\a[28] ), .out0(new_n304));
  nano22aa1n02x4               g209(.a(new_n303), .b(new_n302), .c(new_n304), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n288), .b(new_n269), .c(new_n239), .d(new_n271), .o1(new_n306));
  nona22aa1n03x5               g211(.a(new_n306), .b(new_n293), .c(new_n291), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n299), .b(new_n307), .c(new_n191), .d(new_n289), .o1(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n304), .b(new_n308), .c(new_n302), .o1(new_n309));
  nor002aa1n02x5               g214(.a(new_n309), .b(new_n305), .o1(\s[28] ));
  norb02aa1n02x5               g215(.a(new_n299), .b(new_n304), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n307), .c(new_n191), .d(new_n289), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[28] ), .b(\b[27] ), .c(new_n302), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .out0(new_n314));
  aoi012aa1n02x7               g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  aobi12aa1n02x7               g220(.a(new_n311), .b(new_n290), .c(new_n298), .out0(new_n316));
  nano22aa1n03x5               g221(.a(new_n316), .b(new_n313), .c(new_n314), .out0(new_n317));
  norp02aa1n03x5               g222(.a(new_n315), .b(new_n317), .o1(\s[29] ));
  xorb03aa1n02x5               g223(.a(new_n111), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g224(.a(new_n299), .b(new_n314), .c(new_n304), .out0(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n307), .c(new_n191), .d(new_n289), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .carry(new_n322));
  xnrc02aa1n02x5               g227(.a(\b[29] ), .b(\a[30] ), .out0(new_n323));
  tech160nm_fiaoi012aa1n02p5x5 g228(.a(new_n323), .b(new_n321), .c(new_n322), .o1(new_n324));
  aobi12aa1n02x7               g229(.a(new_n320), .b(new_n290), .c(new_n298), .out0(new_n325));
  nano22aa1n02x4               g230(.a(new_n325), .b(new_n322), .c(new_n323), .out0(new_n326));
  norp02aa1n03x5               g231(.a(new_n324), .b(new_n326), .o1(\s[30] ));
  norb02aa1n02x5               g232(.a(new_n320), .b(new_n323), .out0(new_n328));
  aobi12aa1n02x7               g233(.a(new_n328), .b(new_n290), .c(new_n298), .out0(new_n329));
  oao003aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .c(new_n322), .carry(new_n330));
  xnrc02aa1n02x5               g235(.a(\b[30] ), .b(\a[31] ), .out0(new_n331));
  nano22aa1n03x5               g236(.a(new_n329), .b(new_n330), .c(new_n331), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n328), .b(new_n307), .c(new_n191), .d(new_n289), .o1(new_n333));
  aoi012aa1n03x5               g238(.a(new_n331), .b(new_n333), .c(new_n330), .o1(new_n334));
  nor002aa1n02x5               g239(.a(new_n334), .b(new_n332), .o1(\s[31] ));
  xnrb03aa1n02x5               g240(.a(new_n113), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g241(.a(\a[3] ), .b(\b[2] ), .c(new_n113), .o1(new_n337));
  xorb03aa1n02x5               g242(.a(new_n337), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g243(.a(new_n123), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g244(.a(new_n106), .b(new_n123), .c(new_n107), .o1(new_n340));
  xnrb03aa1n02x5               g245(.a(new_n340), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaib12aa1n02x5               g246(.a(new_n126), .b(new_n108), .c(new_n123), .out0(new_n342));
  xorb03aa1n02x5               g247(.a(new_n342), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g248(.a(new_n101), .b(new_n342), .c(new_n102), .o1(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n344), .b(new_n124), .c(new_n100), .out0(\s[8] ));
  xnbna2aa1n03x5               g250(.a(new_n129), .b(new_n137), .c(new_n139), .out0(\s[9] ));
endmodule


