// Benchmark "adder" written by ABC on Thu Jul 18 03:09:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n338, new_n339, new_n341,
    new_n342, new_n344, new_n345;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n09x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n09x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  inv040aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nor002aa1d24x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand02aa1n02x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oao003aa1n02x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .carry(new_n105));
  nand02aa1n03x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nor022aa1n08x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  norp02aa1n04x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nano23aa1n02x4               g014(.a(new_n108), .b(new_n107), .c(new_n109), .d(new_n106), .out0(new_n110));
  inv030aa1n02x5               g015(.a(new_n107), .o1(new_n111));
  aob012aa1n03x5               g016(.a(new_n111), .b(new_n108), .c(new_n106), .out0(new_n112));
  aoi012aa1n02x5               g017(.a(new_n112), .b(new_n110), .c(new_n105), .o1(new_n113));
  nor042aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand02aa1n03x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor002aa1n03x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nano23aa1n03x5               g022(.a(new_n117), .b(new_n114), .c(new_n115), .d(new_n116), .out0(new_n118));
  norp02aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  tech160nm_finand02aa1n05x5   g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nanb02aa1n09x5               g025(.a(new_n119), .b(new_n120), .out0(new_n121));
  xnrc02aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .out0(new_n122));
  nona22aa1n02x4               g027(.a(new_n118), .b(new_n122), .c(new_n121), .out0(new_n123));
  aoi112aa1n02x5               g028(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n124));
  nona23aa1n03x5               g029(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n125));
  oai022aa1n02x5               g030(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n126));
  nano22aa1n03x5               g031(.a(new_n125), .b(new_n120), .c(new_n126), .out0(new_n127));
  nor003aa1n03x5               g032(.a(new_n127), .b(new_n124), .c(new_n114), .o1(new_n128));
  tech160nm_fioai012aa1n03p5x5 g033(.a(new_n128), .b(new_n123), .c(new_n113), .o1(new_n129));
  xorc02aa1n06x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  aoi012aa1n02x5               g035(.a(new_n101), .b(new_n129), .c(new_n130), .o1(new_n131));
  xnrc02aa1n02x5               g036(.a(new_n131), .b(new_n100), .out0(\s[10] ));
  nanp03aa1n02x5               g037(.a(new_n129), .b(new_n100), .c(new_n130), .o1(new_n133));
  aoi012aa1n02x5               g038(.a(new_n97), .b(new_n101), .c(new_n98), .o1(new_n134));
  xorc02aa1n12x5               g039(.a(\a[11] ), .b(\b[10] ), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  orn002aa1n12x5               g041(.a(\a[11] ), .b(\b[10] ), .o(new_n137));
  inv000aa1d42x5               g042(.a(new_n135), .o1(new_n138));
  aoai13aa1n03x5               g043(.a(new_n137), .b(new_n138), .c(new_n133), .d(new_n134), .o1(new_n139));
  xorb03aa1n02x5               g044(.a(new_n139), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  tech160nm_fioaoi03aa1n03p5x5 g045(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n141));
  nona23aa1n02x4               g046(.a(new_n106), .b(new_n109), .c(new_n108), .d(new_n107), .out0(new_n142));
  oabi12aa1n06x5               g047(.a(new_n112), .b(new_n142), .c(new_n141), .out0(new_n143));
  nor043aa1n02x5               g048(.a(new_n125), .b(new_n121), .c(new_n122), .o1(new_n144));
  nand22aa1n02x5               g049(.a(new_n143), .b(new_n144), .o1(new_n145));
  xnrc02aa1n02x5               g050(.a(\b[11] ), .b(\a[12] ), .out0(new_n146));
  nona23aa1n09x5               g051(.a(new_n135), .b(new_n130), .c(new_n146), .d(new_n99), .out0(new_n147));
  inv000aa1d42x5               g052(.a(\a[12] ), .o1(new_n148));
  inv000aa1d42x5               g053(.a(\b[11] ), .o1(new_n149));
  nand42aa1n06x5               g054(.a(new_n149), .b(new_n148), .o1(new_n150));
  and002aa1n12x5               g055(.a(\b[11] ), .b(\a[12] ), .o(new_n151));
  nand02aa1d04x5               g056(.a(\b[10] ), .b(\a[11] ), .o1(new_n152));
  aoai13aa1n12x5               g057(.a(new_n152), .b(new_n97), .c(new_n101), .d(new_n98), .o1(new_n153));
  aoai13aa1n12x5               g058(.a(new_n150), .b(new_n151), .c(new_n153), .d(new_n137), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n147), .c(new_n128), .d(new_n145), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d28x5               g062(.a(\a[14] ), .o1(new_n158));
  nor042aa1d18x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  tech160nm_fixorc02aa1n02p5x5 g064(.a(\a[13] ), .b(\b[12] ), .out0(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n156), .c(new_n160), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(new_n158), .out0(\s[14] ));
  nand03aa1n02x5               g067(.a(new_n118), .b(new_n120), .c(new_n126), .o1(new_n163));
  nona22aa1n06x5               g068(.a(new_n163), .b(new_n124), .c(new_n114), .out0(new_n164));
  nano32aa1n03x5               g069(.a(new_n146), .b(new_n100), .c(new_n130), .d(new_n135), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n164), .c(new_n143), .d(new_n144), .o1(new_n166));
  xorc02aa1n03x5               g071(.a(\a[14] ), .b(\b[13] ), .out0(new_n167));
  nand42aa1n03x5               g072(.a(new_n167), .b(new_n160), .o1(new_n168));
  inv020aa1d28x5               g073(.a(\b[13] ), .o1(new_n169));
  oaoi03aa1n12x5               g074(.a(new_n158), .b(new_n169), .c(new_n159), .o1(new_n170));
  aoai13aa1n02x7               g075(.a(new_n170), .b(new_n168), .c(new_n166), .d(new_n155), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  xorc02aa1n02x5               g079(.a(\a[16] ), .b(\b[15] ), .out0(new_n175));
  aoi112aa1n02x5               g080(.a(new_n173), .b(new_n175), .c(new_n171), .d(new_n174), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n173), .o1(new_n177));
  inv000aa1d42x5               g082(.a(\a[13] ), .o1(new_n178));
  xroi22aa1d04x5               g083(.a(new_n178), .b(\b[12] ), .c(new_n158), .d(\b[13] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n170), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n174), .b(new_n173), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n180), .c(new_n156), .d(new_n179), .o1(new_n182));
  aobi12aa1n03x5               g087(.a(new_n175), .b(new_n182), .c(new_n177), .out0(new_n183));
  norp02aa1n02x5               g088(.a(new_n183), .b(new_n176), .o1(\s[16] ));
  nor042aa1n02x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nand42aa1n08x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nano23aa1n03x5               g091(.a(new_n173), .b(new_n185), .c(new_n186), .d(new_n174), .out0(new_n187));
  nano22aa1n03x7               g092(.a(new_n147), .b(new_n179), .c(new_n187), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n164), .c(new_n143), .d(new_n144), .o1(new_n189));
  norb02aa1n03x5               g094(.a(new_n187), .b(new_n168), .out0(new_n190));
  norp02aa1n02x5               g095(.a(new_n185), .b(new_n173), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n170), .c(\a[15] ), .d(\b[14] ), .o1(new_n192));
  aoi022aa1d18x5               g097(.a(new_n190), .b(new_n154), .c(new_n192), .d(new_n186), .o1(new_n193));
  xnrc02aa1n02x5               g098(.a(\b[16] ), .b(\a[17] ), .out0(new_n194));
  xobna2aa1n03x5               g099(.a(new_n194), .b(new_n189), .c(new_n193), .out0(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n165), .b(new_n190), .o1(new_n197));
  aoai13aa1n06x5               g102(.a(new_n193), .b(new_n197), .c(new_n145), .d(new_n128), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  aoib12aa1n06x5               g104(.a(new_n199), .b(new_n198), .c(new_n194), .out0(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n196), .out0(\s[18] ));
  inv020aa1d32x5               g106(.a(\a[17] ), .o1(new_n202));
  xroi22aa1d06x4               g107(.a(new_n202), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\b[17] ), .o1(new_n205));
  oao003aa1n02x5               g110(.a(new_n196), .b(new_n205), .c(new_n199), .carry(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n207), .b(new_n204), .c(new_n189), .d(new_n193), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g115(.a(\a[19] ), .o1(new_n211));
  inv030aa1d32x5               g116(.a(\b[18] ), .o1(new_n212));
  nand22aa1n09x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  tech160nm_finand02aa1n03p5x5 g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nor022aa1n12x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand42aa1n06x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  aoi112aa1n02x5               g123(.a(new_n214), .b(new_n218), .c(new_n208), .d(new_n215), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[19] ), .b(\b[18] ), .out0(new_n220));
  aoai13aa1n03x5               g125(.a(new_n220), .b(new_n206), .c(new_n198), .d(new_n203), .o1(new_n221));
  aobi12aa1n03x5               g126(.a(new_n218), .b(new_n221), .c(new_n213), .out0(new_n222));
  nor002aa1n02x5               g127(.a(new_n222), .b(new_n219), .o1(\s[20] ));
  nanb03aa1n09x5               g128(.a(new_n216), .b(new_n217), .c(new_n215), .out0(new_n224));
  nona22aa1n03x5               g129(.a(new_n203), .b(new_n214), .c(new_n224), .out0(new_n225));
  nand42aa1n02x5               g130(.a(\b[17] ), .b(\a[18] ), .o1(new_n226));
  oaih22aa1n04x5               g131(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n227));
  nand23aa1n03x5               g132(.a(new_n227), .b(new_n213), .c(new_n226), .o1(new_n228));
  aoai13aa1n04x5               g133(.a(new_n217), .b(new_n216), .c(new_n211), .d(new_n212), .o1(new_n229));
  oai012aa1n18x5               g134(.a(new_n229), .b(new_n228), .c(new_n224), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n225), .c(new_n189), .d(new_n193), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[21] ), .b(\a[22] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoi112aa1n02x5               g143(.a(new_n234), .b(new_n238), .c(new_n232), .d(new_n236), .o1(new_n239));
  inv000aa1n02x5               g144(.a(new_n225), .o1(new_n240));
  aoai13aa1n04x5               g145(.a(new_n236), .b(new_n230), .c(new_n198), .d(new_n240), .o1(new_n241));
  oaoi13aa1n06x5               g146(.a(new_n237), .b(new_n241), .c(\a[21] ), .d(\b[20] ), .o1(new_n242));
  norp02aa1n03x5               g147(.a(new_n242), .b(new_n239), .o1(\s[22] ));
  nor042aa1n06x5               g148(.a(new_n237), .b(new_n235), .o1(new_n244));
  nona23aa1d18x5               g149(.a(new_n203), .b(new_n244), .c(new_n224), .d(new_n214), .out0(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oao003aa1n12x5               g152(.a(new_n246), .b(new_n247), .c(new_n234), .carry(new_n248));
  aoi012aa1d18x5               g153(.a(new_n248), .b(new_n230), .c(new_n244), .o1(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n245), .c(new_n189), .d(new_n193), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  xorc02aa1n12x5               g158(.a(\a[24] ), .b(\b[23] ), .out0(new_n254));
  aoi112aa1n02x5               g159(.a(new_n252), .b(new_n254), .c(new_n250), .d(new_n253), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n252), .o1(new_n256));
  inv040aa1n03x5               g161(.a(new_n245), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n249), .o1(new_n258));
  aoai13aa1n03x5               g163(.a(new_n253), .b(new_n258), .c(new_n198), .d(new_n257), .o1(new_n259));
  aobi12aa1n03x5               g164(.a(new_n254), .b(new_n259), .c(new_n256), .out0(new_n260));
  nor002aa1n02x5               g165(.a(new_n260), .b(new_n255), .o1(\s[24] ));
  nano32aa1n03x7               g166(.a(new_n225), .b(new_n254), .c(new_n244), .d(new_n253), .out0(new_n262));
  inv020aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  nano22aa1n02x4               g168(.a(new_n216), .b(new_n215), .c(new_n217), .out0(new_n264));
  oai012aa1n02x5               g169(.a(new_n226), .b(\b[18] ), .c(\a[19] ), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n227), .b(new_n265), .out0(new_n266));
  inv000aa1n02x5               g171(.a(new_n229), .o1(new_n267));
  aoai13aa1n04x5               g172(.a(new_n244), .b(new_n267), .c(new_n266), .d(new_n264), .o1(new_n268));
  inv000aa1n02x5               g173(.a(new_n248), .o1(new_n269));
  and002aa1n02x5               g174(.a(new_n254), .b(new_n253), .o(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .carry(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n268), .d(new_n269), .o1(new_n273));
  inv040aa1n03x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n04x5               g179(.a(new_n274), .b(new_n263), .c(new_n189), .d(new_n193), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  xorc02aa1n03x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  xorc02aa1n03x5               g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  aoi112aa1n02x5               g184(.a(new_n277), .b(new_n279), .c(new_n275), .d(new_n278), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n277), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n278), .b(new_n273), .c(new_n198), .d(new_n262), .o1(new_n282));
  aobi12aa1n03x5               g187(.a(new_n279), .b(new_n282), .c(new_n281), .out0(new_n283));
  nor002aa1n02x5               g188(.a(new_n283), .b(new_n280), .o1(\s[26] ));
  nanp02aa1n02x5               g189(.a(new_n192), .b(new_n186), .o1(new_n285));
  aob012aa1n03x5               g190(.a(new_n285), .b(new_n190), .c(new_n154), .out0(new_n286));
  and002aa1n02x5               g191(.a(new_n279), .b(new_n278), .o(new_n287));
  nano22aa1d15x5               g192(.a(new_n245), .b(new_n270), .c(new_n287), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n286), .c(new_n129), .d(new_n188), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[26] ), .b(\b[25] ), .c(new_n281), .carry(new_n290));
  aobi12aa1n06x5               g195(.a(new_n290), .b(new_n273), .c(new_n287), .out0(new_n291));
  xorc02aa1n12x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  xnbna2aa1n03x5               g197(.a(new_n292), .b(new_n291), .c(new_n289), .out0(\s[27] ));
  norp02aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv040aa1n03x5               g199(.a(new_n294), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n292), .o1(new_n296));
  aoi012aa1n02x7               g201(.a(new_n296), .b(new_n291), .c(new_n289), .o1(new_n297));
  xnrc02aa1n12x5               g202(.a(\b[27] ), .b(\a[28] ), .out0(new_n298));
  nano22aa1n03x5               g203(.a(new_n297), .b(new_n295), .c(new_n298), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n270), .b(new_n248), .c(new_n230), .d(new_n244), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n287), .o1(new_n301));
  aoai13aa1n04x5               g206(.a(new_n290), .b(new_n301), .c(new_n300), .d(new_n272), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n292), .b(new_n302), .c(new_n198), .d(new_n288), .o1(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n298), .b(new_n303), .c(new_n295), .o1(new_n304));
  norp02aa1n03x5               g209(.a(new_n304), .b(new_n299), .o1(\s[28] ));
  xnrc02aa1n02x5               g210(.a(\b[28] ), .b(\a[29] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n292), .b(new_n298), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n302), .c(new_n198), .d(new_n288), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n309));
  aoi012aa1n03x5               g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  inv000aa1n02x5               g215(.a(new_n307), .o1(new_n311));
  aoi012aa1n02x7               g216(.a(new_n311), .b(new_n291), .c(new_n289), .o1(new_n312));
  nano22aa1n02x4               g217(.a(new_n312), .b(new_n306), .c(new_n309), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n310), .b(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g220(.a(new_n292), .b(new_n306), .c(new_n298), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n302), .c(new_n198), .d(new_n288), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .carry(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .out0(new_n319));
  aoi012aa1n02x7               g224(.a(new_n319), .b(new_n317), .c(new_n318), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n316), .o1(new_n321));
  aoi012aa1n02x7               g226(.a(new_n321), .b(new_n291), .c(new_n289), .o1(new_n322));
  nano22aa1n02x4               g227(.a(new_n322), .b(new_n318), .c(new_n319), .out0(new_n323));
  norp02aa1n03x5               g228(.a(new_n320), .b(new_n323), .o1(\s[30] ));
  norb02aa1n09x5               g229(.a(new_n316), .b(new_n319), .out0(new_n325));
  inv000aa1n02x5               g230(.a(new_n325), .o1(new_n326));
  aoi012aa1n02x7               g231(.a(new_n326), .b(new_n291), .c(new_n289), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n318), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  nano22aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n329), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n325), .b(new_n302), .c(new_n198), .d(new_n288), .o1(new_n331));
  aoi012aa1n02x7               g236(.a(new_n329), .b(new_n331), .c(new_n328), .o1(new_n332));
  norp02aa1n03x5               g237(.a(new_n332), .b(new_n330), .o1(\s[31] ));
  xnrb03aa1n02x5               g238(.a(new_n141), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi122aa1n02x5               g239(.a(new_n108), .b(new_n106), .c(new_n111), .d(new_n105), .e(new_n109), .o1(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n111), .c(new_n143), .o1(\s[4] ));
  xorb03aa1n02x5               g241(.a(new_n143), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g242(.a(new_n121), .o1(new_n338));
  oao003aa1n03x5               g243(.a(\a[5] ), .b(\b[4] ), .c(new_n113), .carry(new_n339));
  xnrc02aa1n02x5               g244(.a(new_n339), .b(new_n338), .out0(\s[6] ));
  norb02aa1n02x5               g245(.a(new_n116), .b(new_n117), .out0(new_n341));
  nanp02aa1n02x5               g246(.a(new_n339), .b(new_n338), .o1(new_n342));
  xobna2aa1n03x5               g247(.a(new_n341), .b(new_n342), .c(new_n120), .out0(\s[7] ));
  orn002aa1n02x5               g248(.a(\a[8] ), .b(\b[7] ), .o(new_n344));
  aoi013aa1n03x5               g249(.a(new_n117), .b(new_n342), .c(new_n120), .d(new_n116), .o1(new_n345));
  xnbna2aa1n03x5               g250(.a(new_n345), .b(new_n344), .c(new_n115), .out0(\s[8] ));
  xnbna2aa1n03x5               g251(.a(new_n130), .b(new_n128), .c(new_n145), .out0(\s[9] ));
endmodule


