// Benchmark "adder" written by ABC on Thu Jul 18 06:47:07 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n353, new_n354, new_n357, new_n359, new_n360, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor022aa1n16x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nand22aa1n09x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand02aa1n08x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  norp02aa1n12x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nano23aa1n03x7               g006(.a(new_n101), .b(new_n98), .c(new_n99), .d(new_n100), .out0(new_n102));
  nand42aa1n02x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nanb02aa1n06x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  inv040aa1d32x5               g010(.a(\a[5] ), .o1(new_n106));
  inv040aa1d28x5               g011(.a(\b[4] ), .o1(new_n107));
  nand02aa1d24x5               g012(.a(new_n107), .b(new_n106), .o1(new_n108));
  nand42aa1n03x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nanp02aa1n04x5               g014(.a(new_n108), .b(new_n109), .o1(new_n110));
  nona22aa1n02x4               g015(.a(new_n102), .b(new_n105), .c(new_n110), .out0(new_n111));
  nor042aa1n06x5               g016(.a(\b[1] ), .b(\a[2] ), .o1(new_n112));
  inv000aa1n02x5               g017(.a(new_n112), .o1(new_n113));
  nand22aa1n04x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nand02aa1d04x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  aob012aa1n02x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .out0(new_n116));
  nand02aa1n06x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  nor002aa1n03x5               g022(.a(\b[3] ), .b(\a[4] ), .o1(new_n118));
  norb02aa1n02x5               g023(.a(new_n117), .b(new_n118), .out0(new_n119));
  nor042aa1n02x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  nand42aa1n02x5               g025(.a(\b[2] ), .b(\a[3] ), .o1(new_n121));
  norb02aa1n06x4               g026(.a(new_n121), .b(new_n120), .out0(new_n122));
  nanp03aa1n03x5               g027(.a(new_n116), .b(new_n119), .c(new_n122), .o1(new_n123));
  aoi012aa1n09x5               g028(.a(new_n118), .b(new_n120), .c(new_n117), .o1(new_n124));
  oaoi03aa1n12x5               g029(.a(\a[6] ), .b(\b[5] ), .c(new_n108), .o1(new_n125));
  tech160nm_fiao0012aa1n04x5   g030(.a(new_n98), .b(new_n101), .c(new_n99), .o(new_n126));
  aoi012aa1n06x5               g031(.a(new_n126), .b(new_n102), .c(new_n125), .o1(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n111), .c(new_n123), .d(new_n124), .o1(new_n128));
  tech160nm_fixorc02aa1n02p5x5 g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  aoi012aa1n02x5               g034(.a(new_n97), .b(new_n128), .c(new_n129), .o1(new_n130));
  xnrb03aa1n02x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nona23aa1d18x5               g036(.a(new_n100), .b(new_n99), .c(new_n101), .d(new_n98), .out0(new_n132));
  nor043aa1d12x5               g037(.a(new_n132), .b(new_n105), .c(new_n110), .o1(new_n133));
  aoi012aa1n09x5               g038(.a(new_n112), .b(new_n114), .c(new_n115), .o1(new_n134));
  inv000aa1d42x5               g039(.a(\b[3] ), .o1(new_n135));
  nanb02aa1n12x5               g040(.a(\a[4] ), .b(new_n135), .out0(new_n136));
  nand02aa1n03x5               g041(.a(new_n136), .b(new_n117), .o1(new_n137));
  inv040aa1d32x5               g042(.a(\a[3] ), .o1(new_n138));
  inv000aa1d42x5               g043(.a(\b[2] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n139), .b(new_n138), .o1(new_n140));
  nand42aa1n02x5               g045(.a(new_n140), .b(new_n121), .o1(new_n141));
  oai013aa1n06x5               g046(.a(new_n124), .b(new_n134), .c(new_n137), .d(new_n141), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n125), .o1(new_n143));
  oabi12aa1n18x5               g048(.a(new_n126), .b(new_n143), .c(new_n132), .out0(new_n144));
  aoai13aa1n03x5               g049(.a(new_n129), .b(new_n144), .c(new_n142), .d(new_n133), .o1(new_n145));
  nor042aa1n06x5               g050(.a(\b[9] ), .b(\a[10] ), .o1(new_n146));
  norp02aa1n02x5               g051(.a(new_n146), .b(new_n97), .o1(new_n147));
  aoi022aa1n06x5               g052(.a(new_n145), .b(new_n147), .c(\b[9] ), .d(\a[10] ), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n12x5               g054(.a(\b[10] ), .b(\a[11] ), .o1(new_n150));
  nand42aa1n03x5               g055(.a(\b[10] ), .b(\a[11] ), .o1(new_n151));
  xorc02aa1n12x5               g056(.a(\a[12] ), .b(\b[11] ), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n150), .c(new_n148), .d(new_n151), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n152), .b(new_n150), .c(new_n148), .d(new_n151), .o1(new_n154));
  norb02aa1n02x7               g059(.a(new_n153), .b(new_n154), .out0(\s[12] ));
  nor003aa1n02x5               g060(.a(new_n134), .b(new_n137), .c(new_n141), .o1(new_n156));
  inv020aa1n02x5               g061(.a(new_n124), .o1(new_n157));
  tech160nm_fioai012aa1n05x5   g062(.a(new_n133), .b(new_n156), .c(new_n157), .o1(new_n158));
  nand42aa1n03x5               g063(.a(\b[9] ), .b(\a[10] ), .o1(new_n159));
  nano23aa1n03x5               g064(.a(new_n146), .b(new_n150), .c(new_n151), .d(new_n159), .out0(new_n160));
  nand23aa1n03x5               g065(.a(new_n160), .b(new_n129), .c(new_n152), .o1(new_n161));
  inv000aa1d42x5               g066(.a(\b[11] ), .o1(new_n162));
  inv000aa1n02x5               g067(.a(new_n150), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(\a[12] ), .b(new_n162), .out0(new_n164));
  aoi022aa1d24x5               g069(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n165));
  oai012aa1n04x7               g070(.a(new_n165), .b(new_n146), .c(new_n97), .o1(new_n166));
  nand43aa1n02x5               g071(.a(new_n166), .b(new_n163), .c(new_n164), .o1(new_n167));
  oaib12aa1n06x5               g072(.a(new_n167), .b(new_n162), .c(\a[12] ), .out0(new_n168));
  aoai13aa1n06x5               g073(.a(new_n168), .b(new_n161), .c(new_n158), .d(new_n127), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n16x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nand02aa1n03x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  xnrb03aa1n02x5               g078(.a(new_n173), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nona23aa1n02x4               g079(.a(new_n151), .b(new_n159), .c(new_n146), .d(new_n150), .out0(new_n175));
  nano22aa1n02x4               g080(.a(new_n175), .b(new_n129), .c(new_n152), .out0(new_n176));
  aoai13aa1n03x5               g081(.a(new_n176), .b(new_n144), .c(new_n142), .d(new_n133), .o1(new_n177));
  nor042aa1d18x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nanp02aa1n04x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nona23aa1n03x5               g084(.a(new_n179), .b(new_n172), .c(new_n171), .d(new_n178), .out0(new_n180));
  oa0012aa1n02x5               g085(.a(new_n179), .b(new_n178), .c(new_n171), .o(new_n181));
  inv000aa1n02x5               g086(.a(new_n181), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n180), .c(new_n177), .d(new_n168), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  nano23aa1n06x5               g091(.a(new_n171), .b(new_n178), .c(new_n179), .d(new_n172), .out0(new_n187));
  nand22aa1n12x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  nanb02aa1d36x5               g093(.a(new_n185), .b(new_n188), .out0(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  aoai13aa1n03x5               g095(.a(new_n190), .b(new_n181), .c(new_n169), .d(new_n187), .o1(new_n191));
  nor042aa1n06x5               g096(.a(\b[15] ), .b(\a[16] ), .o1(new_n192));
  nand22aa1n09x5               g097(.a(\b[15] ), .b(\a[16] ), .o1(new_n193));
  nanb02aa1d24x5               g098(.a(new_n192), .b(new_n193), .out0(new_n194));
  tech160nm_fiaoi012aa1n05x5   g099(.a(new_n194), .b(new_n191), .c(new_n186), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n194), .o1(new_n196));
  aoi112aa1n03x4               g101(.a(new_n185), .b(new_n196), .c(new_n183), .d(new_n188), .o1(new_n197));
  norp02aa1n02x5               g102(.a(new_n195), .b(new_n197), .o1(\s[16] ));
  nona22aa1n09x5               g103(.a(new_n187), .b(new_n189), .c(new_n194), .out0(new_n199));
  nor042aa1n06x5               g104(.a(new_n161), .b(new_n199), .o1(new_n200));
  aoai13aa1n12x5               g105(.a(new_n200), .b(new_n144), .c(new_n142), .d(new_n133), .o1(new_n201));
  and002aa1n02x5               g106(.a(\b[11] ), .b(\a[12] ), .o(new_n202));
  aoi013aa1n06x4               g107(.a(new_n202), .b(new_n166), .c(new_n163), .d(new_n164), .o1(new_n203));
  nor043aa1n03x5               g108(.a(new_n180), .b(new_n189), .c(new_n194), .o1(new_n204));
  oai112aa1n02x5               g109(.a(new_n179), .b(new_n188), .c(new_n178), .d(new_n171), .o1(new_n205));
  nona22aa1n03x5               g110(.a(new_n205), .b(new_n192), .c(new_n185), .out0(new_n206));
  aoi022aa1n12x5               g111(.a(new_n203), .b(new_n204), .c(new_n193), .d(new_n206), .o1(new_n207));
  xorc02aa1n12x5               g112(.a(\a[17] ), .b(\b[16] ), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n201), .c(new_n207), .out0(\s[17] ));
  nor002aa1d32x5               g114(.a(\b[16] ), .b(\a[17] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(new_n206), .b(new_n193), .o1(new_n212));
  tech160nm_fioai012aa1n04x5   g117(.a(new_n212), .b(new_n168), .c(new_n199), .o1(new_n213));
  aoai13aa1n02x5               g118(.a(new_n208), .b(new_n213), .c(new_n128), .d(new_n200), .o1(new_n214));
  xnrc02aa1n12x5               g119(.a(\b[17] ), .b(\a[18] ), .out0(new_n215));
  xobna2aa1n03x5               g120(.a(new_n215), .b(new_n214), .c(new_n211), .out0(\s[18] ));
  inv000aa1d42x5               g121(.a(\a[17] ), .o1(new_n217));
  inv040aa1d32x5               g122(.a(\a[18] ), .o1(new_n218));
  xroi22aa1d04x5               g123(.a(new_n217), .b(\b[16] ), .c(new_n218), .d(\b[17] ), .out0(new_n219));
  inv030aa1n02x5               g124(.a(new_n219), .o1(new_n220));
  oaoi03aa1n12x5               g125(.a(\a[18] ), .b(\b[17] ), .c(new_n211), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n222), .b(new_n220), .c(new_n201), .d(new_n207), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g130(.a(\b[18] ), .b(\a[19] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nanp02aa1n02x5               g132(.a(new_n176), .b(new_n204), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n207), .b(new_n228), .c(new_n158), .d(new_n127), .o1(new_n229));
  nand02aa1n20x5               g134(.a(\b[18] ), .b(\a[19] ), .o1(new_n230));
  nanb02aa1d36x5               g135(.a(new_n226), .b(new_n230), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n221), .c(new_n229), .d(new_n219), .o1(new_n233));
  xnrc02aa1n06x5               g138(.a(\b[19] ), .b(\a[20] ), .out0(new_n234));
  tech160nm_fiaoi012aa1n02p5x5 g139(.a(new_n234), .b(new_n233), .c(new_n227), .o1(new_n235));
  inv040aa1n02x5               g140(.a(new_n234), .o1(new_n236));
  aoi112aa1n03x4               g141(.a(new_n226), .b(new_n236), .c(new_n223), .d(new_n230), .o1(new_n237));
  norp02aa1n03x5               g142(.a(new_n235), .b(new_n237), .o1(\s[20] ));
  nona23aa1d24x5               g143(.a(new_n236), .b(new_n208), .c(new_n215), .d(new_n231), .out0(new_n239));
  norp02aa1n06x5               g144(.a(\b[17] ), .b(\a[18] ), .o1(new_n240));
  nanp02aa1n02x5               g145(.a(\b[17] ), .b(\a[18] ), .o1(new_n241));
  oai112aa1n04x5               g146(.a(new_n241), .b(new_n230), .c(new_n240), .d(new_n210), .o1(new_n242));
  oab012aa1n06x5               g147(.a(new_n226), .b(\a[20] ), .c(\b[19] ), .out0(new_n243));
  aoi022aa1n12x5               g148(.a(new_n242), .b(new_n243), .c(\b[19] ), .d(\a[20] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n239), .c(new_n201), .d(new_n207), .o1(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n16x5               g152(.a(\b[20] ), .b(\a[21] ), .o1(new_n248));
  inv040aa1n03x5               g153(.a(new_n248), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n239), .o1(new_n250));
  nanp02aa1n04x5               g155(.a(\b[20] ), .b(\a[21] ), .o1(new_n251));
  norb02aa1n02x5               g156(.a(new_n251), .b(new_n248), .out0(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n244), .c(new_n229), .d(new_n250), .o1(new_n253));
  inv040aa1d32x5               g158(.a(\a[22] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\b[21] ), .o1(new_n255));
  nand22aa1n09x5               g160(.a(new_n255), .b(new_n254), .o1(new_n256));
  nand02aa1d06x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  nand22aa1n12x5               g162(.a(new_n256), .b(new_n257), .o1(new_n258));
  tech160nm_fiaoi012aa1n02p5x5 g163(.a(new_n258), .b(new_n253), .c(new_n249), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n258), .o1(new_n260));
  aoi112aa1n03x4               g165(.a(new_n248), .b(new_n260), .c(new_n246), .d(new_n252), .o1(new_n261));
  nor002aa1n02x5               g166(.a(new_n259), .b(new_n261), .o1(\s[22] ));
  nano22aa1n03x7               g167(.a(new_n258), .b(new_n249), .c(new_n251), .out0(new_n263));
  nano32aa1n02x4               g168(.a(new_n220), .b(new_n263), .c(new_n232), .d(new_n236), .out0(new_n264));
  inv020aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  nanp02aa1n06x5               g170(.a(new_n242), .b(new_n243), .o1(new_n266));
  nand42aa1n02x5               g171(.a(\b[19] ), .b(\a[20] ), .o1(new_n267));
  nano32aa1n09x5               g172(.a(new_n258), .b(new_n249), .c(new_n251), .d(new_n267), .out0(new_n268));
  oaoi03aa1n09x5               g173(.a(new_n254), .b(new_n255), .c(new_n248), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  aoi012aa1n09x5               g175(.a(new_n270), .b(new_n266), .c(new_n268), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n265), .c(new_n201), .d(new_n207), .o1(new_n272));
  xorb03aa1n02x5               g177(.a(new_n272), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g178(.a(\b[22] ), .b(\a[23] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n274), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n271), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[23] ), .b(\b[22] ), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n276), .c(new_n229), .d(new_n264), .o1(new_n278));
  xorc02aa1n12x5               g183(.a(\a[24] ), .b(\b[23] ), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n278), .c(new_n275), .o1(new_n281));
  aoi112aa1n03x4               g186(.a(new_n274), .b(new_n279), .c(new_n272), .d(new_n277), .o1(new_n282));
  nor002aa1n02x5               g187(.a(new_n281), .b(new_n282), .o1(\s[24] ));
  nano32aa1n02x5               g188(.a(new_n239), .b(new_n279), .c(new_n263), .d(new_n277), .out0(new_n284));
  inv000aa1n02x5               g189(.a(new_n284), .o1(new_n285));
  nor002aa1n02x5               g190(.a(new_n240), .b(new_n210), .o1(new_n286));
  nano22aa1n02x5               g191(.a(new_n286), .b(new_n241), .c(new_n230), .out0(new_n287));
  inv040aa1n03x5               g192(.a(new_n243), .o1(new_n288));
  oai012aa1n06x5               g193(.a(new_n268), .b(new_n287), .c(new_n288), .o1(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[22] ), .b(\a[23] ), .out0(new_n290));
  norb02aa1n12x5               g195(.a(new_n279), .b(new_n290), .out0(new_n291));
  inv000aa1n06x5               g196(.a(new_n291), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[24] ), .b(\b[23] ), .c(new_n275), .carry(new_n293));
  aoai13aa1n06x5               g198(.a(new_n293), .b(new_n292), .c(new_n289), .d(new_n269), .o1(new_n294));
  inv040aa1n02x5               g199(.a(new_n294), .o1(new_n295));
  aoai13aa1n04x5               g200(.a(new_n295), .b(new_n285), .c(new_n201), .d(new_n207), .o1(new_n296));
  xorb03aa1n02x5               g201(.a(new_n296), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g202(.a(\b[24] ), .b(\a[25] ), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n298), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[25] ), .b(\b[24] ), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n294), .c(new_n229), .d(new_n284), .o1(new_n301));
  xorc02aa1n12x5               g206(.a(\a[26] ), .b(\b[25] ), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n301), .c(new_n299), .o1(new_n304));
  aoi112aa1n03x4               g209(.a(new_n298), .b(new_n302), .c(new_n296), .d(new_n300), .o1(new_n305));
  nor002aa1n02x5               g210(.a(new_n304), .b(new_n305), .o1(\s[26] ));
  nand02aa1d08x5               g211(.a(new_n302), .b(new_n300), .o1(new_n307));
  nano23aa1d15x5               g212(.a(new_n239), .b(new_n307), .c(new_n291), .d(new_n263), .out0(new_n308));
  aoai13aa1n06x5               g213(.a(new_n308), .b(new_n213), .c(new_n128), .d(new_n200), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n307), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[26] ), .b(\b[25] ), .c(new_n299), .carry(new_n311));
  inv000aa1d42x5               g216(.a(new_n311), .o1(new_n312));
  aoi012aa1n12x5               g217(.a(new_n312), .b(new_n294), .c(new_n310), .o1(new_n313));
  xorc02aa1n12x5               g218(.a(\a[27] ), .b(\b[26] ), .out0(new_n314));
  xnbna2aa1n03x5               g219(.a(new_n314), .b(new_n313), .c(new_n309), .out0(\s[27] ));
  norp02aa1n02x5               g220(.a(\b[26] ), .b(\a[27] ), .o1(new_n316));
  inv040aa1n03x5               g221(.a(new_n316), .o1(new_n317));
  aoai13aa1n04x5               g222(.a(new_n291), .b(new_n270), .c(new_n266), .d(new_n268), .o1(new_n318));
  aoai13aa1n06x5               g223(.a(new_n311), .b(new_n307), .c(new_n318), .d(new_n293), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n314), .b(new_n319), .c(new_n229), .d(new_n308), .o1(new_n320));
  xnrc02aa1n02x5               g225(.a(\b[27] ), .b(\a[28] ), .out0(new_n321));
  tech160nm_fiaoi012aa1n02p5x5 g226(.a(new_n321), .b(new_n320), .c(new_n317), .o1(new_n322));
  aobi12aa1n02x7               g227(.a(new_n314), .b(new_n313), .c(new_n309), .out0(new_n323));
  nano22aa1n03x5               g228(.a(new_n323), .b(new_n317), .c(new_n321), .out0(new_n324));
  norp02aa1n03x5               g229(.a(new_n322), .b(new_n324), .o1(\s[28] ));
  norb02aa1n02x5               g230(.a(new_n314), .b(new_n321), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n319), .c(new_n229), .d(new_n308), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[28] ), .b(\b[27] ), .c(new_n317), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[28] ), .b(\a[29] ), .out0(new_n329));
  tech160nm_fiaoi012aa1n02p5x5 g234(.a(new_n329), .b(new_n327), .c(new_n328), .o1(new_n330));
  aobi12aa1n02x7               g235(.a(new_n326), .b(new_n313), .c(new_n309), .out0(new_n331));
  nano22aa1n03x5               g236(.a(new_n331), .b(new_n328), .c(new_n329), .out0(new_n332));
  norp02aa1n03x5               g237(.a(new_n330), .b(new_n332), .o1(\s[29] ));
  xorb03aa1n02x5               g238(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g239(.a(new_n314), .b(new_n329), .c(new_n321), .out0(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n319), .c(new_n229), .d(new_n308), .o1(new_n336));
  oao003aa1n02x5               g241(.a(\a[29] ), .b(\b[28] ), .c(new_n328), .carry(new_n337));
  xnrc02aa1n02x5               g242(.a(\b[29] ), .b(\a[30] ), .out0(new_n338));
  tech160nm_fiaoi012aa1n02p5x5 g243(.a(new_n338), .b(new_n336), .c(new_n337), .o1(new_n339));
  aobi12aa1n02x7               g244(.a(new_n335), .b(new_n313), .c(new_n309), .out0(new_n340));
  nano22aa1n03x5               g245(.a(new_n340), .b(new_n337), .c(new_n338), .out0(new_n341));
  norp02aa1n03x5               g246(.a(new_n339), .b(new_n341), .o1(\s[30] ));
  xnrc02aa1n02x5               g247(.a(\b[30] ), .b(\a[31] ), .out0(new_n343));
  nona32aa1n02x4               g248(.a(new_n314), .b(new_n338), .c(new_n329), .d(new_n321), .out0(new_n344));
  aoi012aa1n02x7               g249(.a(new_n344), .b(new_n313), .c(new_n309), .o1(new_n345));
  oao003aa1n02x5               g250(.a(\a[30] ), .b(\b[29] ), .c(new_n337), .carry(new_n346));
  nano22aa1n03x5               g251(.a(new_n345), .b(new_n343), .c(new_n346), .out0(new_n347));
  inv000aa1n02x5               g252(.a(new_n344), .o1(new_n348));
  aoai13aa1n03x5               g253(.a(new_n348), .b(new_n319), .c(new_n229), .d(new_n308), .o1(new_n349));
  tech160nm_fiaoi012aa1n02p5x5 g254(.a(new_n343), .b(new_n349), .c(new_n346), .o1(new_n350));
  norp02aa1n03x5               g255(.a(new_n350), .b(new_n347), .o1(\s[31] ));
  xnbna2aa1n03x5               g256(.a(new_n134), .b(new_n121), .c(new_n140), .out0(\s[3] ));
  aoai13aa1n02x5               g257(.a(new_n122), .b(new_n112), .c(new_n115), .d(new_n114), .o1(new_n353));
  aoi022aa1n02x5               g258(.a(new_n136), .b(new_n117), .c(new_n138), .d(new_n139), .o1(new_n354));
  aoi022aa1n02x5               g259(.a(new_n142), .b(new_n136), .c(new_n354), .d(new_n353), .o1(\s[4] ));
  xorb03aa1n02x5               g260(.a(new_n142), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n02x5               g261(.a(new_n108), .b(new_n110), .c(new_n123), .d(new_n124), .o1(new_n357));
  xorb03aa1n02x5               g262(.a(new_n357), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  orn002aa1n02x5               g263(.a(new_n105), .b(new_n110), .o(new_n359));
  aoai13aa1n02x5               g264(.a(new_n143), .b(new_n359), .c(new_n123), .d(new_n124), .o1(new_n360));
  xorb03aa1n02x5               g265(.a(new_n360), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g266(.a(new_n101), .b(new_n360), .c(new_n100), .o1(new_n362));
  xnrb03aa1n02x5               g267(.a(new_n362), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g268(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


