// Benchmark "adder" written by ABC on Wed Jul 17 15:57:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n347, new_n349, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n357, new_n358, new_n360, new_n362, new_n363, new_n364;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n08x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n10x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n03x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  norp02aa1n24x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv040aa1d32x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nand22aa1n12x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nand22aa1n12x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  aob012aa1n12x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .out0(new_n107));
  nor042aa1n06x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand22aa1n09x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  norb02aa1n06x5               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  nor042aa1n06x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nand22aa1n03x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  norb02aa1n09x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nanp03aa1d12x5               g018(.a(new_n107), .b(new_n110), .c(new_n113), .o1(new_n114));
  aoi012aa1n12x5               g019(.a(new_n108), .b(new_n111), .c(new_n109), .o1(new_n115));
  nor042aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand22aa1n03x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand22aa1n12x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nor002aa1d32x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano23aa1n03x7               g024(.a(new_n119), .b(new_n116), .c(new_n117), .d(new_n118), .out0(new_n120));
  nor042aa1n06x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nand22aa1n12x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  nand22aa1n12x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nor042aa1d18x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nano23aa1n09x5               g029(.a(new_n124), .b(new_n121), .c(new_n122), .d(new_n123), .out0(new_n125));
  nand02aa1d04x5               g030(.a(new_n125), .b(new_n120), .o1(new_n126));
  inv040aa1n06x5               g031(.a(new_n119), .o1(new_n127));
  oaoi03aa1n12x5               g032(.a(\a[6] ), .b(\b[5] ), .c(new_n127), .o1(new_n128));
  tech160nm_fiaoi012aa1n03p5x5 g033(.a(new_n121), .b(new_n124), .c(new_n122), .o1(new_n129));
  aobi12aa1n12x5               g034(.a(new_n129), .b(new_n125), .c(new_n128), .out0(new_n130));
  aoai13aa1n12x5               g035(.a(new_n130), .b(new_n126), .c(new_n114), .d(new_n115), .o1(new_n131));
  tech160nm_fixorc02aa1n03p5x5 g036(.a(\a[9] ), .b(\b[8] ), .out0(new_n132));
  nand22aa1n03x5               g037(.a(new_n131), .b(new_n132), .o1(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n99), .b(new_n133), .c(new_n101), .out0(\s[10] ));
  nor022aa1n16x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand42aa1n20x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  inv000aa1d42x5               g042(.a(\a[10] ), .o1(new_n138));
  aoai13aa1n03x5               g043(.a(new_n98), .b(new_n100), .c(new_n131), .d(new_n132), .o1(new_n139));
  oaib12aa1n03x5               g044(.a(new_n139), .b(\b[9] ), .c(new_n138), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n133), .b(new_n101), .o1(new_n141));
  oai012aa1n02x5               g046(.a(new_n98), .b(new_n141), .c(new_n97), .o1(new_n142));
  mtn022aa1n02x5               g047(.a(new_n140), .b(new_n142), .sa(new_n137), .o1(\s[11] ));
  nor002aa1d32x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n08x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nanb02aa1n02x5               g050(.a(new_n144), .b(new_n145), .out0(new_n146));
  aoai13aa1n02x5               g051(.a(new_n146), .b(new_n135), .c(new_n140), .d(new_n136), .o1(new_n147));
  aoai13aa1n04x5               g052(.a(new_n137), .b(new_n97), .c(new_n141), .d(new_n98), .o1(new_n148));
  nona22aa1n02x4               g053(.a(new_n148), .b(new_n146), .c(new_n135), .out0(new_n149));
  nanp02aa1n03x5               g054(.a(new_n147), .b(new_n149), .o1(\s[12] ));
  nano32aa1n03x7               g055(.a(new_n146), .b(new_n132), .c(new_n137), .d(new_n99), .out0(new_n151));
  nanp02aa1n06x5               g056(.a(new_n131), .b(new_n151), .o1(new_n152));
  nano22aa1n03x7               g057(.a(new_n144), .b(new_n136), .c(new_n145), .out0(new_n153));
  aoi012aa1n02x7               g058(.a(new_n135), .b(\a[10] ), .c(\b[9] ), .o1(new_n154));
  oai112aa1n06x5               g059(.a(new_n153), .b(new_n154), .c(new_n100), .d(new_n97), .o1(new_n155));
  aoi012aa1n06x5               g060(.a(new_n144), .b(new_n135), .c(new_n145), .o1(new_n156));
  nanp02aa1n09x5               g061(.a(new_n155), .b(new_n156), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nanp02aa1n06x5               g063(.a(new_n152), .b(new_n158), .o1(new_n159));
  nor002aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand42aa1n16x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  nano22aa1n02x4               g067(.a(new_n162), .b(new_n155), .c(new_n156), .out0(new_n163));
  aoi022aa1n02x5               g068(.a(new_n159), .b(new_n162), .c(new_n152), .d(new_n163), .o1(\s[13] ));
  tech160nm_fiaoi012aa1n05x5   g069(.a(new_n160), .b(new_n159), .c(new_n161), .o1(new_n165));
  xnrb03aa1n03x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n03x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand02aa1n12x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nano23aa1d15x5               g073(.a(new_n160), .b(new_n167), .c(new_n168), .d(new_n161), .out0(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n157), .c(new_n131), .d(new_n151), .o1(new_n170));
  oa0012aa1n02x5               g075(.a(new_n168), .b(new_n167), .c(new_n160), .o(new_n171));
  nanb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  nor042aa1n03x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n06x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  oai022aa1d18x5               g080(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n176));
  aboi22aa1n03x5               g081(.a(new_n173), .b(new_n174), .c(new_n176), .d(new_n168), .out0(new_n177));
  aoi022aa1n02x5               g082(.a(new_n172), .b(new_n175), .c(new_n170), .d(new_n177), .o1(\s[15] ));
  xorc02aa1n12x5               g083(.a(\a[16] ), .b(\b[15] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  aoai13aa1n02x7               g085(.a(new_n180), .b(new_n173), .c(new_n172), .d(new_n174), .o1(new_n181));
  aoai13aa1n04x5               g086(.a(new_n175), .b(new_n171), .c(new_n159), .d(new_n169), .o1(new_n182));
  nona22aa1n02x4               g087(.a(new_n182), .b(new_n180), .c(new_n173), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n181), .b(new_n183), .o1(\s[16] ));
  nano23aa1n02x4               g089(.a(new_n135), .b(new_n144), .c(new_n145), .d(new_n136), .out0(new_n185));
  nand23aa1n09x5               g090(.a(new_n169), .b(new_n175), .c(new_n179), .o1(new_n186));
  nano32aa1n03x7               g091(.a(new_n186), .b(new_n185), .c(new_n132), .d(new_n99), .out0(new_n187));
  nand02aa1n06x5               g092(.a(new_n131), .b(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\a[16] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[15] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n190), .b(new_n189), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(\b[15] ), .b(\a[16] ), .o1(new_n192));
  nanp03aa1n02x5               g097(.a(new_n191), .b(new_n174), .c(new_n192), .o1(new_n193));
  oai112aa1n02x5               g098(.a(new_n176), .b(new_n168), .c(\b[14] ), .d(\a[15] ), .o1(new_n194));
  nor042aa1n02x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  tech160nm_fioaoi03aa1n03p5x5 g100(.a(new_n189), .b(new_n190), .c(new_n173), .o1(new_n196));
  norb02aa1n03x5               g101(.a(new_n196), .b(new_n195), .out0(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n186), .c(new_n155), .d(new_n156), .o1(new_n198));
  inv040aa1n03x5               g103(.a(new_n198), .o1(new_n199));
  nanp02aa1n06x5               g104(.a(new_n188), .b(new_n199), .o1(new_n200));
  xorc02aa1n02x5               g105(.a(\a[17] ), .b(\b[16] ), .out0(new_n201));
  nona22aa1n02x4               g106(.a(new_n196), .b(new_n195), .c(new_n201), .out0(new_n202));
  aoib12aa1n02x5               g107(.a(new_n202), .b(new_n157), .c(new_n186), .out0(new_n203));
  aoi022aa1n02x5               g108(.a(new_n200), .b(new_n201), .c(new_n188), .d(new_n203), .o1(\s[17] ));
  inv040aa1d32x5               g109(.a(\a[18] ), .o1(new_n205));
  nor042aa1n06x5               g110(.a(\b[16] ), .b(\a[17] ), .o1(new_n206));
  tech160nm_fiaoi012aa1n05x5   g111(.a(new_n206), .b(new_n200), .c(new_n201), .o1(new_n207));
  xorb03aa1n02x5               g112(.a(new_n207), .b(\b[17] ), .c(new_n205), .out0(\s[18] ));
  inv000aa1d42x5               g113(.a(\a[17] ), .o1(new_n209));
  xroi22aa1d06x4               g114(.a(new_n209), .b(\b[16] ), .c(new_n205), .d(\b[17] ), .out0(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n198), .c(new_n131), .d(new_n187), .o1(new_n211));
  nand02aa1n06x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nor042aa1n06x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  nor002aa1n03x5               g118(.a(new_n213), .b(new_n206), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n212), .b(new_n214), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  nor042aa1n04x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nand02aa1d08x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  norb02aa1n06x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n211), .c(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g125(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n06x5               g126(.a(new_n211), .b(new_n216), .o1(new_n222));
  nor042aa1n09x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nand02aa1d24x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  nanb02aa1n03x5               g129(.a(new_n223), .b(new_n224), .out0(new_n225));
  aoai13aa1n02x5               g130(.a(new_n225), .b(new_n217), .c(new_n222), .d(new_n218), .o1(new_n226));
  nanp02aa1n02x5               g131(.a(new_n222), .b(new_n219), .o1(new_n227));
  nona22aa1n02x4               g132(.a(new_n227), .b(new_n225), .c(new_n217), .out0(new_n228));
  nanp02aa1n02x5               g133(.a(new_n228), .b(new_n226), .o1(\s[20] ));
  nanb03aa1d18x5               g134(.a(new_n225), .b(new_n210), .c(new_n219), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n198), .c(new_n131), .d(new_n187), .o1(new_n232));
  nanb03aa1n02x5               g137(.a(new_n223), .b(new_n224), .c(new_n218), .out0(new_n233));
  orn002aa1n02x5               g138(.a(\a[19] ), .b(\b[18] ), .o(new_n234));
  oai112aa1n02x5               g139(.a(new_n234), .b(new_n212), .c(new_n213), .d(new_n206), .o1(new_n235));
  aoi012aa1n09x5               g140(.a(new_n223), .b(new_n217), .c(new_n224), .o1(new_n236));
  oai012aa1n04x7               g141(.a(new_n236), .b(new_n235), .c(new_n233), .o1(new_n237));
  nanb02aa1n02x5               g142(.a(new_n237), .b(new_n232), .out0(new_n238));
  xorc02aa1n12x5               g143(.a(\a[21] ), .b(\b[20] ), .out0(new_n239));
  nano22aa1n12x5               g144(.a(new_n223), .b(new_n218), .c(new_n224), .out0(new_n240));
  oai012aa1n06x5               g145(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .o1(new_n241));
  oab012aa1n02x4               g146(.a(new_n241), .b(new_n206), .c(new_n213), .out0(new_n242));
  inv000aa1n03x5               g147(.a(new_n236), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(new_n243), .b(new_n239), .c(new_n242), .d(new_n240), .o1(new_n244));
  aoi022aa1n02x5               g149(.a(new_n238), .b(new_n239), .c(new_n232), .d(new_n244), .o1(\s[21] ));
  nor042aa1d18x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[21] ), .b(\a[22] ), .out0(new_n247));
  aoai13aa1n03x5               g152(.a(new_n247), .b(new_n246), .c(new_n238), .d(new_n239), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n239), .b(new_n237), .c(new_n200), .d(new_n231), .o1(new_n249));
  nona22aa1n03x5               g154(.a(new_n249), .b(new_n247), .c(new_n246), .out0(new_n250));
  nanp02aa1n03x5               g155(.a(new_n248), .b(new_n250), .o1(\s[22] ));
  xnrc02aa1n02x5               g156(.a(\b[20] ), .b(\a[21] ), .out0(new_n252));
  nona32aa1n02x4               g157(.a(new_n200), .b(new_n247), .c(new_n252), .d(new_n230), .out0(new_n253));
  nor002aa1n04x5               g158(.a(new_n247), .b(new_n252), .o1(new_n254));
  nanb02aa1n03x5               g159(.a(new_n230), .b(new_n254), .out0(new_n255));
  nona22aa1n09x5               g160(.a(new_n240), .b(new_n214), .c(new_n241), .out0(new_n256));
  nanb02aa1n12x5               g161(.a(new_n247), .b(new_n239), .out0(new_n257));
  inv000aa1d42x5               g162(.a(\a[22] ), .o1(new_n258));
  inv040aa1d32x5               g163(.a(\b[21] ), .o1(new_n259));
  oao003aa1n03x5               g164(.a(new_n258), .b(new_n259), .c(new_n246), .carry(new_n260));
  inv040aa1n03x5               g165(.a(new_n260), .o1(new_n261));
  aoai13aa1n12x5               g166(.a(new_n261), .b(new_n257), .c(new_n256), .d(new_n236), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n04x5               g168(.a(new_n263), .b(new_n255), .c(new_n188), .d(new_n199), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[23] ), .b(\b[22] ), .out0(new_n265));
  aoi112aa1n02x5               g170(.a(new_n265), .b(new_n260), .c(new_n237), .d(new_n254), .o1(new_n266));
  aoi022aa1n02x5               g171(.a(new_n266), .b(new_n253), .c(new_n264), .d(new_n265), .o1(\s[23] ));
  nor002aa1n03x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  xnrc02aa1n12x5               g173(.a(\b[23] ), .b(\a[24] ), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n268), .c(new_n264), .d(new_n265), .o1(new_n270));
  nand42aa1n02x5               g175(.a(new_n264), .b(new_n265), .o1(new_n271));
  nona22aa1n03x5               g176(.a(new_n271), .b(new_n269), .c(new_n268), .out0(new_n272));
  nanp02aa1n03x5               g177(.a(new_n272), .b(new_n270), .o1(\s[24] ));
  norb02aa1n06x5               g178(.a(new_n265), .b(new_n269), .out0(new_n274));
  nano22aa1n03x7               g179(.a(new_n230), .b(new_n254), .c(new_n274), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n198), .c(new_n131), .d(new_n187), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n254), .b(new_n243), .c(new_n242), .d(new_n240), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n274), .o1(new_n278));
  inv000aa1d42x5               g183(.a(\a[24] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(\b[23] ), .o1(new_n280));
  tech160nm_fioaoi03aa1n03p5x5 g185(.a(new_n279), .b(new_n280), .c(new_n268), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n281), .b(new_n278), .c(new_n277), .d(new_n261), .o1(new_n282));
  nanb02aa1n06x5               g187(.a(new_n282), .b(new_n276), .out0(new_n283));
  xorc02aa1n12x5               g188(.a(\a[25] ), .b(\b[24] ), .out0(new_n284));
  inv000aa1d42x5               g189(.a(new_n281), .o1(new_n285));
  aoi112aa1n02x5               g190(.a(new_n284), .b(new_n285), .c(new_n262), .d(new_n274), .o1(new_n286));
  aoi022aa1n02x5               g191(.a(new_n283), .b(new_n284), .c(new_n276), .d(new_n286), .o1(\s[25] ));
  norp02aa1n02x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  tech160nm_fixnrc02aa1n04x5   g193(.a(\b[25] ), .b(\a[26] ), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n288), .c(new_n283), .d(new_n284), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n284), .b(new_n282), .c(new_n200), .d(new_n275), .o1(new_n291));
  nona22aa1n03x5               g196(.a(new_n291), .b(new_n289), .c(new_n288), .out0(new_n292));
  nanp02aa1n03x5               g197(.a(new_n290), .b(new_n292), .o1(\s[26] ));
  norb02aa1n06x5               g198(.a(new_n284), .b(new_n289), .out0(new_n294));
  nano32aa1d12x5               g199(.a(new_n230), .b(new_n294), .c(new_n254), .d(new_n274), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n198), .c(new_n131), .d(new_n187), .o1(new_n296));
  aoi112aa1n02x5               g201(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n297));
  oab012aa1n02x4               g202(.a(new_n297), .b(\a[26] ), .c(\b[25] ), .out0(new_n298));
  aobi12aa1n06x5               g203(.a(new_n298), .b(new_n282), .c(new_n294), .out0(new_n299));
  tech160nm_fixorc02aa1n05x5   g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  xnbna2aa1n03x5               g205(.a(new_n300), .b(new_n299), .c(new_n296), .out0(\s[27] ));
  aoai13aa1n02x7               g206(.a(new_n294), .b(new_n285), .c(new_n262), .d(new_n274), .o1(new_n302));
  nand43aa1n03x5               g207(.a(new_n296), .b(new_n302), .c(new_n298), .o1(new_n303));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  norp02aa1n02x5               g209(.a(\b[27] ), .b(\a[28] ), .o1(new_n305));
  nanp02aa1n02x5               g210(.a(\b[27] ), .b(\a[28] ), .o1(new_n306));
  nanb02aa1n09x5               g211(.a(new_n305), .b(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n304), .c(new_n303), .d(new_n300), .o1(new_n308));
  aoai13aa1n02x5               g213(.a(new_n274), .b(new_n260), .c(new_n237), .d(new_n254), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n294), .o1(new_n310));
  aoai13aa1n02x7               g215(.a(new_n298), .b(new_n310), .c(new_n309), .d(new_n281), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n300), .b(new_n311), .c(new_n200), .d(new_n295), .o1(new_n312));
  nona22aa1n02x4               g217(.a(new_n312), .b(new_n307), .c(new_n304), .out0(new_n313));
  nanp02aa1n03x5               g218(.a(new_n308), .b(new_n313), .o1(\s[28] ));
  norb02aa1n06x5               g219(.a(new_n300), .b(new_n307), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n200), .d(new_n295), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  oai012aa1n02x5               g222(.a(new_n306), .b(new_n305), .c(new_n304), .o1(new_n318));
  norb02aa1n02x5               g223(.a(new_n318), .b(new_n317), .out0(new_n319));
  inv000aa1n02x5               g224(.a(new_n315), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n318), .b(new_n320), .c(new_n299), .d(new_n296), .o1(new_n321));
  aoi022aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n316), .d(new_n319), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g228(.a(new_n307), .b(new_n317), .c(new_n300), .out0(new_n324));
  nanb02aa1n03x5               g229(.a(new_n324), .b(new_n303), .out0(new_n325));
  inv000aa1d42x5               g230(.a(\b[28] ), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\a[29] ), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n318), .b(\b[28] ), .c(new_n327), .out0(new_n328));
  oaib12aa1n02x5               g233(.a(new_n328), .b(new_n326), .c(\a[29] ), .out0(new_n329));
  aoai13aa1n02x7               g234(.a(new_n329), .b(new_n324), .c(new_n299), .d(new_n296), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .out0(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n331), .b(new_n328), .c(new_n327), .d(new_n326), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n325), .d(new_n332), .o1(\s[30] ));
  nano22aa1n06x5               g238(.a(new_n320), .b(new_n317), .c(new_n331), .out0(new_n334));
  aoai13aa1n03x5               g239(.a(new_n334), .b(new_n311), .c(new_n200), .d(new_n295), .o1(new_n335));
  aoi022aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n336));
  norb02aa1n02x5               g241(.a(\a[31] ), .b(\b[30] ), .out0(new_n337));
  obai22aa1n02x7               g242(.a(\b[30] ), .b(\a[31] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n338));
  aoi112aa1n02x5               g243(.a(new_n338), .b(new_n337), .c(new_n328), .d(new_n336), .o1(new_n339));
  inv000aa1d42x5               g244(.a(new_n334), .o1(new_n340));
  norp02aa1n02x5               g245(.a(\b[29] ), .b(\a[30] ), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n341), .b(new_n328), .c(new_n336), .o1(new_n342));
  aoai13aa1n02x7               g247(.a(new_n342), .b(new_n340), .c(new_n299), .d(new_n296), .o1(new_n343));
  xorc02aa1n02x5               g248(.a(\a[31] ), .b(\b[30] ), .out0(new_n344));
  aoi022aa1n02x7               g249(.a(new_n343), .b(new_n344), .c(new_n339), .d(new_n335), .o1(\s[31] ));
  xorb03aa1n02x5               g250(.a(new_n107), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oai012aa1n02x5               g251(.a(new_n112), .b(new_n107), .c(new_n111), .o1(new_n347));
  xnrc02aa1n02x5               g252(.a(new_n347), .b(new_n110), .out0(\s[4] ));
  norb02aa1n02x5               g253(.a(new_n118), .b(new_n119), .out0(new_n349));
  xnbna2aa1n03x5               g254(.a(new_n349), .b(new_n114), .c(new_n115), .out0(\s[5] ));
  norb02aa1n02x5               g255(.a(new_n117), .b(new_n116), .out0(new_n351));
  oaoi03aa1n02x5               g256(.a(new_n102), .b(new_n103), .c(new_n105), .o1(new_n352));
  nona23aa1n02x4               g257(.a(new_n112), .b(new_n109), .c(new_n108), .d(new_n111), .out0(new_n353));
  oai012aa1n02x5               g258(.a(new_n115), .b(new_n353), .c(new_n352), .o1(new_n354));
  nanp02aa1n02x5               g259(.a(new_n354), .b(new_n349), .o1(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n351), .b(new_n355), .c(new_n127), .out0(\s[6] ));
  aobi12aa1n02x5               g261(.a(new_n351), .b(new_n355), .c(new_n127), .out0(new_n357));
  norp02aa1n02x5               g262(.a(new_n357), .b(new_n116), .o1(new_n358));
  xnrb03aa1n02x5               g263(.a(new_n358), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oai013aa1n02x4               g264(.a(new_n123), .b(new_n357), .c(new_n124), .d(new_n116), .o1(new_n360));
  xnrb03aa1n02x5               g265(.a(new_n360), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  nanb02aa1n02x5               g266(.a(new_n126), .b(new_n354), .out0(new_n362));
  tech160nm_fiao0012aa1n02p5x5 g267(.a(new_n121), .b(new_n124), .c(new_n122), .o(new_n363));
  aoi112aa1n02x5               g268(.a(new_n132), .b(new_n363), .c(new_n125), .d(new_n128), .o1(new_n364));
  aoi022aa1n02x5               g269(.a(new_n131), .b(new_n132), .c(new_n362), .d(new_n364), .o1(\s[9] ));
endmodule


