// Benchmark "adder" written by ABC on Thu Jul 18 10:21:13 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n315, new_n317,
    new_n318, new_n321, new_n322, new_n324, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n06x5               g001(.a(\a[10] ), .b(\b[9] ), .o(new_n97));
  nand42aa1n03x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n02x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  xnrc02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .out0(new_n103));
  xnrc02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .out0(new_n104));
  orn002aa1n02x5               g009(.a(\a[4] ), .b(\b[3] ), .o(new_n105));
  aoi112aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n106));
  norb02aa1n03x5               g011(.a(new_n105), .b(new_n106), .out0(new_n107));
  oai013aa1n02x4               g012(.a(new_n107), .b(new_n102), .c(new_n103), .d(new_n104), .o1(new_n108));
  xorc02aa1n02x5               g013(.a(\a[6] ), .b(\b[5] ), .out0(new_n109));
  tech160nm_fixorc02aa1n02p5x5 g014(.a(\a[5] ), .b(\b[4] ), .out0(new_n110));
  xorc02aa1n12x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  nor042aa1n06x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanb02aa1n02x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  nano32aa1n02x4               g019(.a(new_n114), .b(new_n111), .c(new_n110), .d(new_n109), .out0(new_n115));
  nanp02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nano22aa1n09x5               g021(.a(new_n112), .b(new_n116), .c(new_n113), .out0(new_n117));
  oai022aa1n06x5               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(new_n112), .o1(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  aoi013aa1n09x5               g025(.a(new_n120), .b(new_n117), .c(new_n111), .d(new_n118), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n121), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  aoai13aa1n03x5               g028(.a(new_n123), .b(new_n122), .c(new_n115), .d(new_n108), .o1(new_n124));
  oa0012aa1n02x5               g029(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .o(new_n125));
  oai112aa1n06x5               g030(.a(new_n97), .b(new_n98), .c(\b[8] ), .d(\a[9] ), .o1(new_n126));
  nanb02aa1n06x5               g031(.a(new_n126), .b(new_n124), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n97), .d(new_n98), .o1(\s[10] ));
  nand42aa1n03x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  norp02aa1n04x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanb03aa1n02x5               g035(.a(new_n130), .b(new_n98), .c(new_n129), .out0(new_n131));
  nanb02aa1n02x5               g036(.a(new_n130), .b(new_n129), .out0(new_n132));
  oao003aa1n02x5               g037(.a(new_n99), .b(new_n100), .c(new_n101), .carry(new_n133));
  xorc02aa1n02x5               g038(.a(\a[4] ), .b(\b[3] ), .out0(new_n134));
  xorc02aa1n02x5               g039(.a(\a[3] ), .b(\b[2] ), .out0(new_n135));
  nanp03aa1n02x5               g040(.a(new_n133), .b(new_n134), .c(new_n135), .o1(new_n136));
  xnrc02aa1n02x5               g041(.a(\b[5] ), .b(\a[6] ), .out0(new_n137));
  nona23aa1n09x5               g042(.a(new_n110), .b(new_n111), .c(new_n137), .d(new_n114), .out0(new_n138));
  aoai13aa1n12x5               g043(.a(new_n121), .b(new_n138), .c(new_n136), .d(new_n107), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n98), .b(new_n126), .c(new_n139), .d(new_n123), .o1(new_n140));
  aboi22aa1n03x5               g045(.a(new_n131), .b(new_n127), .c(new_n140), .d(new_n132), .out0(\s[11] ));
  nor002aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n03x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  aoi113aa1n02x5               g049(.a(new_n144), .b(new_n130), .c(new_n127), .d(new_n129), .e(new_n98), .o1(new_n145));
  aoib12aa1n02x5               g050(.a(new_n130), .b(new_n127), .c(new_n131), .out0(new_n146));
  aoib12aa1n02x5               g051(.a(new_n145), .b(new_n144), .c(new_n146), .out0(\s[12] ));
  nanp02aa1n02x5               g052(.a(new_n97), .b(new_n98), .o1(new_n148));
  nona23aa1d18x5               g053(.a(new_n144), .b(new_n123), .c(new_n148), .d(new_n132), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  tech160nm_fiaoi012aa1n04x5   g055(.a(new_n130), .b(\a[10] ), .c(\b[9] ), .o1(new_n151));
  nano22aa1n03x7               g056(.a(new_n142), .b(new_n129), .c(new_n143), .out0(new_n152));
  tech160nm_fiao0012aa1n02p5x5 g057(.a(new_n142), .b(new_n130), .c(new_n143), .o(new_n153));
  aoi013aa1n09x5               g058(.a(new_n153), .b(new_n152), .c(new_n126), .d(new_n151), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  xorc02aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .out0(new_n156));
  aoai13aa1n02x5               g061(.a(new_n156), .b(new_n155), .c(new_n139), .d(new_n150), .o1(new_n157));
  aoi112aa1n02x5               g062(.a(new_n156), .b(new_n155), .c(new_n139), .d(new_n150), .o1(new_n158));
  norb02aa1n02x5               g063(.a(new_n157), .b(new_n158), .out0(\s[13] ));
  inv000aa1d42x5               g064(.a(\a[13] ), .o1(new_n160));
  nanb02aa1n12x5               g065(.a(\b[12] ), .b(new_n160), .out0(new_n161));
  xorc02aa1n02x5               g066(.a(\a[14] ), .b(\b[13] ), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n157), .c(new_n161), .out0(\s[14] ));
  inv000aa1d42x5               g068(.a(\a[14] ), .o1(new_n164));
  xroi22aa1d04x5               g069(.a(new_n160), .b(\b[12] ), .c(new_n164), .d(\b[13] ), .out0(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n155), .c(new_n139), .d(new_n150), .o1(new_n166));
  tech160nm_fioaoi03aa1n05x5   g071(.a(\a[14] ), .b(\b[13] ), .c(new_n161), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  xorc02aa1n12x5               g073(.a(\a[15] ), .b(\b[14] ), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n166), .c(new_n168), .out0(\s[15] ));
  aob012aa1n02x5               g075(.a(new_n169), .b(new_n166), .c(new_n168), .out0(new_n171));
  xorc02aa1n02x5               g076(.a(\a[16] ), .b(\b[15] ), .out0(new_n172));
  norp02aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norp02aa1n02x5               g078(.a(new_n172), .b(new_n173), .o1(new_n174));
  inv000aa1n03x5               g079(.a(new_n173), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n169), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n175), .b(new_n176), .c(new_n166), .d(new_n168), .o1(new_n177));
  aoi022aa1n02x5               g082(.a(new_n177), .b(new_n172), .c(new_n171), .d(new_n174), .o1(\s[16] ));
  nanp02aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  xnrc02aa1n02x5               g084(.a(\b[15] ), .b(\a[16] ), .out0(new_n180));
  nano22aa1n02x4               g085(.a(new_n180), .b(new_n175), .c(new_n179), .out0(new_n181));
  nano22aa1d15x5               g086(.a(new_n149), .b(new_n165), .c(new_n181), .out0(new_n182));
  aoai13aa1n03x5               g087(.a(new_n182), .b(new_n122), .c(new_n115), .d(new_n108), .o1(new_n183));
  nanp02aa1n02x5               g088(.a(new_n165), .b(new_n181), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(\a[16] ), .b(\b[15] ), .c(new_n175), .o1(new_n185));
  aoi013aa1n06x4               g090(.a(new_n185), .b(new_n167), .c(new_n169), .d(new_n172), .o1(new_n186));
  oai012aa1n18x5               g091(.a(new_n186), .b(new_n154), .c(new_n184), .o1(new_n187));
  nanb02aa1n06x5               g092(.a(new_n187), .b(new_n183), .out0(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  nanb02aa1n02x5               g095(.a(\b[16] ), .b(new_n190), .out0(new_n191));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  aoai13aa1n02x5               g097(.a(new_n192), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n193));
  xorc02aa1n02x5               g098(.a(\a[18] ), .b(\b[17] ), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n193), .c(new_n191), .out0(\s[18] ));
  inv000aa1d42x5               g100(.a(\a[18] ), .o1(new_n196));
  xroi22aa1d04x5               g101(.a(new_n190), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n197));
  aoai13aa1n02x5               g102(.a(new_n197), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n198));
  oai022aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n199));
  oaib12aa1n02x5               g104(.a(new_n199), .b(new_n196), .c(\b[17] ), .out0(new_n200));
  nor042aa1n06x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nanb02aa1n02x5               g107(.a(new_n201), .b(new_n202), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n198), .c(new_n200), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n02x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n191), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n204), .b(new_n207), .c(new_n188), .d(new_n197), .o1(new_n208));
  nor042aa1n02x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanp02aa1n02x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  aoib12aa1n02x5               g116(.a(new_n201), .b(new_n210), .c(new_n209), .out0(new_n212));
  inv000aa1n02x5               g117(.a(new_n201), .o1(new_n213));
  aoai13aa1n02x5               g118(.a(new_n213), .b(new_n203), .c(new_n198), .d(new_n200), .o1(new_n214));
  aoi022aa1n02x5               g119(.a(new_n214), .b(new_n211), .c(new_n208), .d(new_n212), .o1(\s[20] ));
  nano23aa1n06x5               g120(.a(new_n201), .b(new_n209), .c(new_n210), .d(new_n202), .out0(new_n216));
  nand23aa1n04x5               g121(.a(new_n216), .b(new_n192), .c(new_n194), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n02x5               g123(.a(new_n218), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n219));
  nona23aa1n09x5               g124(.a(new_n210), .b(new_n202), .c(new_n201), .d(new_n209), .out0(new_n220));
  oaoi03aa1n02x5               g125(.a(\a[20] ), .b(\b[19] ), .c(new_n213), .o1(new_n221));
  oabi12aa1n12x5               g126(.a(new_n221), .b(new_n220), .c(new_n200), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  xnrc02aa1n12x5               g128(.a(\b[20] ), .b(\a[21] ), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n219), .c(new_n223), .out0(\s[21] ));
  aoai13aa1n02x5               g131(.a(new_n225), .b(new_n222), .c(new_n188), .d(new_n218), .o1(new_n227));
  xnrc02aa1n02x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  nor042aa1n06x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n228), .b(new_n229), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n229), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n231), .b(new_n224), .c(new_n219), .d(new_n223), .o1(new_n232));
  aboi22aa1n03x5               g137(.a(new_n228), .b(new_n232), .c(new_n227), .d(new_n230), .out0(\s[22] ));
  nor042aa1n04x5               g138(.a(new_n228), .b(new_n224), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n217), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n236));
  oao003aa1n12x5               g141(.a(\a[22] ), .b(\b[21] ), .c(new_n231), .carry(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(new_n222), .c(new_n234), .o1(new_n239));
  xorc02aa1n12x5               g144(.a(\a[23] ), .b(\b[22] ), .out0(new_n240));
  aob012aa1n03x5               g145(.a(new_n240), .b(new_n236), .c(new_n239), .out0(new_n241));
  aoi112aa1n02x5               g146(.a(new_n240), .b(new_n238), .c(new_n222), .d(new_n234), .o1(new_n242));
  aobi12aa1n02x7               g147(.a(new_n241), .b(new_n242), .c(new_n236), .out0(\s[23] ));
  xorc02aa1n02x5               g148(.a(\a[24] ), .b(\b[23] ), .out0(new_n244));
  nor042aa1n03x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  norp02aa1n02x5               g150(.a(new_n244), .b(new_n245), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n245), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n240), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n247), .b(new_n248), .c(new_n236), .d(new_n239), .o1(new_n249));
  aoi022aa1n02x5               g154(.a(new_n249), .b(new_n244), .c(new_n241), .d(new_n246), .o1(\s[24] ));
  nano32aa1n03x7               g155(.a(new_n217), .b(new_n244), .c(new_n234), .d(new_n240), .out0(new_n251));
  aoai13aa1n02x5               g156(.a(new_n251), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n234), .b(new_n221), .c(new_n216), .d(new_n207), .o1(new_n253));
  and002aa1n02x5               g158(.a(new_n244), .b(new_n240), .o(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  oao003aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n247), .carry(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n255), .c(new_n253), .d(new_n237), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[25] ), .b(\b[24] ), .out0(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n252), .c(new_n258), .out0(\s[25] ));
  aoai13aa1n03x5               g165(.a(new_n259), .b(new_n257), .c(new_n188), .d(new_n251), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .out0(new_n262));
  nor042aa1n03x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  norp02aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n263), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n259), .o1(new_n266));
  aoai13aa1n02x5               g171(.a(new_n265), .b(new_n266), .c(new_n252), .d(new_n258), .o1(new_n267));
  aoi022aa1n02x5               g172(.a(new_n267), .b(new_n262), .c(new_n261), .d(new_n264), .o1(\s[26] ));
  and002aa1n06x5               g173(.a(new_n262), .b(new_n259), .o(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  nano23aa1d12x5               g175(.a(new_n270), .b(new_n217), .c(new_n254), .d(new_n234), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n187), .c(new_n139), .d(new_n182), .o1(new_n272));
  oao003aa1n02x5               g177(.a(\a[26] ), .b(\b[25] ), .c(new_n265), .carry(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  aoi012aa1n12x5               g179(.a(new_n274), .b(new_n257), .c(new_n269), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n272), .out0(\s[27] ));
  aoai13aa1n04x5               g182(.a(new_n254), .b(new_n238), .c(new_n222), .d(new_n234), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n273), .b(new_n270), .c(new_n278), .d(new_n256), .o1(new_n279));
  aoai13aa1n02x5               g184(.a(new_n276), .b(new_n279), .c(new_n188), .d(new_n271), .o1(new_n280));
  xorc02aa1n02x5               g185(.a(\a[28] ), .b(\b[27] ), .out0(new_n281));
  norp02aa1n02x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  norp02aa1n02x5               g187(.a(new_n281), .b(new_n282), .o1(new_n283));
  inv000aa1n03x5               g188(.a(new_n282), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n276), .o1(new_n285));
  aoai13aa1n02x5               g190(.a(new_n284), .b(new_n285), .c(new_n275), .d(new_n272), .o1(new_n286));
  aoi022aa1n02x5               g191(.a(new_n286), .b(new_n281), .c(new_n280), .d(new_n283), .o1(\s[28] ));
  and002aa1n02x5               g192(.a(new_n281), .b(new_n276), .o(new_n288));
  aoai13aa1n02x5               g193(.a(new_n288), .b(new_n279), .c(new_n188), .d(new_n271), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n288), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n284), .carry(new_n291));
  aoai13aa1n02x5               g196(.a(new_n291), .b(new_n290), .c(new_n275), .d(new_n272), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .out0(new_n293));
  norb02aa1n02x5               g198(.a(new_n291), .b(new_n293), .out0(new_n294));
  aoi022aa1n03x5               g199(.a(new_n292), .b(new_n293), .c(new_n289), .d(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d33x5               g201(.a(new_n285), .b(new_n281), .c(new_n293), .out0(new_n297));
  aoai13aa1n02x5               g202(.a(new_n297), .b(new_n279), .c(new_n188), .d(new_n271), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n297), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n300));
  aoai13aa1n02x5               g205(.a(new_n300), .b(new_n299), .c(new_n275), .d(new_n272), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[30] ), .b(\b[29] ), .out0(new_n302));
  norb02aa1n02x5               g207(.a(new_n300), .b(new_n302), .out0(new_n303));
  aoi022aa1n02x5               g208(.a(new_n301), .b(new_n302), .c(new_n298), .d(new_n303), .o1(\s[30] ));
  nano32aa1d15x5               g209(.a(new_n285), .b(new_n302), .c(new_n281), .d(new_n293), .out0(new_n305));
  aoai13aa1n02x5               g210(.a(new_n305), .b(new_n279), .c(new_n188), .d(new_n271), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[31] ), .b(\b[30] ), .out0(new_n307));
  and002aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .o(new_n308));
  oabi12aa1n02x5               g213(.a(new_n307), .b(\a[30] ), .c(\b[29] ), .out0(new_n309));
  oab012aa1n02x4               g214(.a(new_n309), .b(new_n300), .c(new_n308), .out0(new_n310));
  inv000aa1d42x5               g215(.a(new_n305), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n312));
  aoai13aa1n02x5               g217(.a(new_n312), .b(new_n311), .c(new_n275), .d(new_n272), .o1(new_n313));
  aoi022aa1n02x5               g218(.a(new_n313), .b(new_n307), .c(new_n306), .d(new_n310), .o1(\s[31] ));
  inv000aa1d42x5               g219(.a(\a[3] ), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n102), .b(\b[2] ), .c(new_n315), .out0(\s[3] ));
  nanp02aa1n02x5               g221(.a(new_n133), .b(new_n135), .o1(new_n317));
  aoib12aa1n02x5               g222(.a(new_n134), .b(new_n315), .c(\b[2] ), .out0(new_n318));
  aoi022aa1n02x5               g223(.a(new_n108), .b(new_n105), .c(new_n318), .d(new_n317), .o1(\s[4] ));
  xnbna2aa1n03x5               g224(.a(new_n110), .b(new_n136), .c(new_n107), .out0(\s[5] ));
  norp02aa1n02x5               g225(.a(\b[4] ), .b(\a[5] ), .o1(new_n321));
  aoi012aa1n02x5               g226(.a(new_n321), .b(new_n108), .c(new_n110), .o1(new_n322));
  xnrc02aa1n02x5               g227(.a(new_n322), .b(new_n109), .out0(\s[6] ));
  nanp02aa1n02x5               g228(.a(new_n322), .b(new_n109), .o1(new_n324));
  xnbna2aa1n03x5               g229(.a(new_n114), .b(new_n324), .c(new_n116), .out0(\s[7] ));
  nanp02aa1n02x5               g230(.a(new_n324), .b(new_n117), .o1(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n111), .b(new_n326), .c(new_n119), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n139), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


