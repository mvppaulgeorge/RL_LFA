// Benchmark "adder" written by ABC on Thu Jul 18 10:49:57 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n319, new_n322, new_n323, new_n325, new_n326, new_n327,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oao003aa1n02x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n101));
  nor002aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor042aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano23aa1n02x4               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  oa0012aa1n02x5               g011(.a(new_n103), .b(new_n104), .c(new_n102), .o(new_n107));
  nand42aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb03aa1n06x5               g015(.a(new_n109), .b(new_n110), .c(new_n108), .out0(new_n111));
  norp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanb02aa1n02x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  inv000aa1d42x5               g019(.a(\a[5] ), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\b[4] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(new_n116), .b(new_n115), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  oai112aa1n02x5               g023(.a(new_n117), .b(new_n118), .c(\b[5] ), .d(\a[6] ), .o1(new_n119));
  nor043aa1n03x5               g024(.a(new_n119), .b(new_n111), .c(new_n114), .o1(new_n120));
  aoai13aa1n02x5               g025(.a(new_n120), .b(new_n107), .c(new_n101), .d(new_n106), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n113), .o1(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  aoi013aa1n02x4               g028(.a(new_n109), .b(new_n123), .c(new_n110), .d(new_n108), .o1(new_n124));
  oab012aa1n02x4               g029(.a(new_n112), .b(new_n124), .c(new_n122), .out0(new_n125));
  nanp02aa1n02x5               g030(.a(new_n125), .b(new_n121), .o1(new_n126));
  nand42aa1n03x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  aoi012aa1n02x5               g032(.a(new_n97), .b(new_n126), .c(new_n127), .o1(new_n128));
  xnrb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nanp02aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norp02aa1n02x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nano23aa1n03x5               g036(.a(new_n97), .b(new_n131), .c(new_n130), .d(new_n127), .out0(new_n132));
  oaih22aa1n04x5               g037(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  ao0022aa1n03x5               g038(.a(new_n126), .b(new_n132), .c(new_n133), .d(new_n130), .o(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  aoi022aa1n02x5               g040(.a(new_n126), .b(new_n132), .c(new_n130), .d(new_n133), .o1(new_n136));
  oaoi03aa1n02x5               g041(.a(\a[11] ), .b(\b[10] ), .c(new_n136), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1n03x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norp02aa1n02x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanp02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nano23aa1n02x4               g047(.a(new_n139), .b(new_n141), .c(new_n142), .d(new_n140), .out0(new_n143));
  nanp02aa1n02x5               g048(.a(new_n143), .b(new_n132), .o1(new_n144));
  nanb03aa1n06x5               g049(.a(new_n139), .b(new_n140), .c(new_n130), .out0(new_n145));
  inv000aa1d42x5               g050(.a(\b[11] ), .o1(new_n146));
  nanb02aa1n02x5               g051(.a(\a[12] ), .b(new_n146), .out0(new_n147));
  nand23aa1n03x5               g052(.a(new_n133), .b(new_n147), .c(new_n142), .o1(new_n148));
  tech160nm_fioai012aa1n03p5x5 g053(.a(new_n142), .b(new_n141), .c(new_n139), .o1(new_n149));
  oai012aa1n18x5               g054(.a(new_n149), .b(new_n148), .c(new_n145), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n144), .c(new_n125), .d(new_n121), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand42aa1n03x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n154), .b(new_n152), .c(new_n155), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  oaoi03aa1n02x5               g062(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n158));
  nona23aa1n02x4               g063(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n159));
  oabi12aa1n06x5               g064(.a(new_n107), .b(new_n158), .c(new_n159), .out0(new_n160));
  oaoi03aa1n02x5               g065(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n161), .b(new_n160), .c(new_n120), .o1(new_n162));
  norp02aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand42aa1n03x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nona23aa1n02x4               g069(.a(new_n164), .b(new_n155), .c(new_n154), .d(new_n163), .out0(new_n165));
  nano23aa1n03x5               g070(.a(new_n154), .b(new_n163), .c(new_n164), .d(new_n155), .out0(new_n166));
  oa0012aa1n02x5               g071(.a(new_n164), .b(new_n163), .c(new_n154), .o(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n150), .c(new_n166), .o1(new_n168));
  oai013aa1n02x5               g073(.a(new_n168), .b(new_n162), .c(new_n144), .d(new_n165), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  xnrb03aa1n03x5               g078(.a(new_n173), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  norp02aa1n02x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nano23aa1n03x7               g081(.a(new_n171), .b(new_n175), .c(new_n176), .d(new_n172), .out0(new_n177));
  nano22aa1n03x7               g082(.a(new_n144), .b(new_n166), .c(new_n177), .out0(new_n178));
  aoai13aa1n03x5               g083(.a(new_n178), .b(new_n161), .c(new_n160), .d(new_n120), .o1(new_n179));
  aoai13aa1n09x5               g084(.a(new_n177), .b(new_n167), .c(new_n150), .d(new_n166), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n176), .b(new_n175), .c(new_n171), .o1(new_n181));
  nand23aa1n06x5               g086(.a(new_n179), .b(new_n180), .c(new_n181), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nona23aa1n02x4               g088(.a(new_n130), .b(new_n127), .c(new_n97), .d(new_n131), .out0(new_n184));
  nona23aa1n02x4               g089(.a(new_n177), .b(new_n143), .c(new_n184), .d(new_n165), .out0(new_n185));
  aoi012aa1n02x7               g090(.a(new_n185), .b(new_n125), .c(new_n121), .o1(new_n186));
  nano22aa1n03x7               g091(.a(new_n186), .b(new_n180), .c(new_n181), .out0(new_n187));
  oaoi03aa1n02x5               g092(.a(\a[17] ), .b(\b[16] ), .c(new_n187), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv040aa1d32x5               g095(.a(\a[18] ), .o1(new_n191));
  xroi22aa1d06x4               g096(.a(new_n190), .b(\b[16] ), .c(new_n191), .d(\b[17] ), .out0(new_n192));
  inv000aa1d42x5               g097(.a(\b[17] ), .o1(new_n193));
  norp02aa1n02x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  oao003aa1n02x5               g099(.a(new_n191), .b(new_n193), .c(new_n194), .carry(new_n195));
  tech160nm_fiaoi012aa1n05x5   g100(.a(new_n195), .b(new_n182), .c(new_n192), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\a[19] ), .o1(new_n197));
  nanb02aa1d24x5               g102(.a(\b[18] ), .b(new_n197), .out0(new_n198));
  nand42aa1d28x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n196), .b(new_n199), .c(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g106(.a(new_n192), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n195), .o1(new_n203));
  oaih12aa1n02x5               g108(.a(new_n203), .b(new_n187), .c(new_n202), .o1(new_n204));
  nor042aa1n04x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  tech160nm_fixorc02aa1n05x5   g110(.a(\a[20] ), .b(\b[19] ), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n207), .b(new_n205), .c(new_n204), .d(new_n199), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n199), .o1(new_n209));
  oai112aa1n03x5               g114(.a(new_n206), .b(new_n198), .c(new_n196), .d(new_n209), .o1(new_n210));
  nanp02aa1n03x5               g115(.a(new_n208), .b(new_n210), .o1(\s[20] ));
  nona23aa1d16x5               g116(.a(new_n192), .b(new_n206), .c(new_n209), .d(new_n205), .out0(new_n212));
  oai112aa1n06x5               g117(.a(new_n198), .b(new_n199), .c(new_n193), .d(new_n191), .o1(new_n213));
  oai022aa1n04x5               g118(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n214));
  inv030aa1d32x5               g119(.a(\a[20] ), .o1(new_n215));
  inv000aa1d42x5               g120(.a(\b[19] ), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(new_n216), .b(new_n215), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand23aa1n06x5               g123(.a(new_n214), .b(new_n217), .c(new_n218), .o1(new_n219));
  tech160nm_fioaoi03aa1n03p5x5 g124(.a(new_n215), .b(new_n216), .c(new_n205), .o1(new_n220));
  oai012aa1d24x5               g125(.a(new_n220), .b(new_n219), .c(new_n213), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oai012aa1n04x7               g127(.a(new_n222), .b(new_n187), .c(new_n212), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xorc02aa1n02x5               g130(.a(\a[21] ), .b(\b[20] ), .out0(new_n226));
  xorc02aa1n02x5               g131(.a(\a[22] ), .b(\b[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n226), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n212), .o1(new_n230));
  aoai13aa1n02x5               g135(.a(new_n226), .b(new_n221), .c(new_n182), .d(new_n230), .o1(new_n231));
  nona22aa1n02x4               g136(.a(new_n231), .b(new_n228), .c(new_n225), .out0(new_n232));
  nanp02aa1n03x5               g137(.a(new_n229), .b(new_n232), .o1(\s[22] ));
  inv000aa1d42x5               g138(.a(\a[21] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(\a[22] ), .o1(new_n235));
  xroi22aa1d04x5               g140(.a(new_n234), .b(\b[20] ), .c(new_n235), .d(\b[21] ), .out0(new_n236));
  norb02aa1n03x5               g141(.a(new_n236), .b(new_n212), .out0(new_n237));
  inv020aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  nanb02aa1n02x5               g143(.a(\b[20] ), .b(new_n234), .out0(new_n239));
  oaoi03aa1n02x5               g144(.a(\a[22] ), .b(\b[21] ), .c(new_n239), .o1(new_n240));
  tech160nm_fiaoi012aa1n03p5x5 g145(.a(new_n240), .b(new_n221), .c(new_n236), .o1(new_n241));
  tech160nm_fioai012aa1n05x5   g146(.a(new_n241), .b(new_n187), .c(new_n238), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  xorc02aa1n02x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  xorc02aa1n12x5               g150(.a(\a[24] ), .b(\b[23] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aoai13aa1n03x5               g152(.a(new_n247), .b(new_n244), .c(new_n242), .d(new_n245), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n241), .o1(new_n249));
  aoai13aa1n02x5               g154(.a(new_n245), .b(new_n249), .c(new_n182), .d(new_n237), .o1(new_n250));
  nona22aa1n02x5               g155(.a(new_n250), .b(new_n247), .c(new_n244), .out0(new_n251));
  nanp02aa1n03x5               g156(.a(new_n248), .b(new_n251), .o1(\s[24] ));
  and002aa1n02x5               g157(.a(new_n246), .b(new_n245), .o(new_n253));
  nano22aa1n03x7               g158(.a(new_n212), .b(new_n253), .c(new_n236), .out0(new_n254));
  inv020aa1n03x5               g159(.a(new_n254), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n253), .b(new_n240), .c(new_n221), .d(new_n236), .o1(new_n256));
  oai022aa1n02x5               g161(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n257));
  aob012aa1n02x5               g162(.a(new_n257), .b(\b[23] ), .c(\a[24] ), .out0(new_n258));
  nand02aa1d04x5               g163(.a(new_n256), .b(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  oai012aa1n04x7               g165(.a(new_n260), .b(new_n187), .c(new_n255), .o1(new_n261));
  xorb03aa1n02x5               g166(.a(new_n261), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  xnrc02aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n263), .c(new_n261), .d(new_n264), .o1(new_n266));
  aoai13aa1n02x5               g171(.a(new_n264), .b(new_n259), .c(new_n182), .d(new_n254), .o1(new_n267));
  nona22aa1n02x5               g172(.a(new_n267), .b(new_n265), .c(new_n263), .out0(new_n268));
  nanp02aa1n03x5               g173(.a(new_n266), .b(new_n268), .o1(\s[26] ));
  norb02aa1n03x5               g174(.a(new_n264), .b(new_n265), .out0(new_n270));
  nano32aa1d12x5               g175(.a(new_n212), .b(new_n270), .c(new_n236), .d(new_n253), .out0(new_n271));
  inv020aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .o1(new_n273));
  oai022aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n274));
  aoi022aa1n02x7               g179(.a(new_n259), .b(new_n270), .c(new_n273), .d(new_n274), .o1(new_n275));
  tech160nm_fioai012aa1n03p5x5 g180(.a(new_n275), .b(new_n187), .c(new_n272), .o1(new_n276));
  xorb03aa1n02x5               g181(.a(new_n276), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n06x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  xorc02aa1n02x5               g184(.a(\a[28] ), .b(\b[27] ), .out0(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n278), .c(new_n276), .d(new_n279), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n270), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n274), .b(new_n273), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n283), .c(new_n256), .d(new_n258), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n279), .b(new_n285), .c(new_n182), .d(new_n271), .o1(new_n286));
  nona22aa1n02x5               g191(.a(new_n286), .b(new_n281), .c(new_n278), .out0(new_n287));
  nanp02aa1n03x5               g192(.a(new_n282), .b(new_n287), .o1(\s[28] ));
  and002aa1n02x5               g193(.a(new_n280), .b(new_n279), .o(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n285), .c(new_n182), .d(new_n271), .o1(new_n290));
  inv000aa1d42x5               g195(.a(\a[28] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\b[27] ), .o1(new_n292));
  oaoi03aa1n12x5               g197(.a(new_n291), .b(new_n292), .c(new_n278), .o1(new_n293));
  xorc02aa1n02x5               g198(.a(\a[29] ), .b(\b[28] ), .out0(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  tech160nm_fiaoi012aa1n03p5x5 g200(.a(new_n295), .b(new_n290), .c(new_n293), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n293), .o1(new_n297));
  nona22aa1n02x5               g202(.a(new_n290), .b(new_n297), .c(new_n294), .out0(new_n298));
  norb02aa1n03x4               g203(.a(new_n298), .b(new_n296), .out0(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g205(.a(new_n295), .b(new_n279), .c(new_n280), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n285), .c(new_n182), .d(new_n271), .o1(new_n302));
  tech160nm_fioaoi03aa1n03p5x5 g207(.a(\a[29] ), .b(\b[28] ), .c(new_n293), .o1(new_n303));
  inv000aa1n03x5               g208(.a(new_n303), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .out0(new_n305));
  aobi12aa1n06x5               g210(.a(new_n305), .b(new_n302), .c(new_n304), .out0(new_n306));
  nona22aa1n02x5               g211(.a(new_n302), .b(new_n303), .c(new_n305), .out0(new_n307));
  norb02aa1n03x4               g212(.a(new_n307), .b(new_n306), .out0(\s[30] ));
  nano32aa1n02x4               g213(.a(new_n295), .b(new_n305), .c(new_n279), .d(new_n280), .out0(new_n309));
  aoai13aa1n06x5               g214(.a(new_n309), .b(new_n285), .c(new_n182), .d(new_n271), .o1(new_n310));
  tech160nm_fioaoi03aa1n05x5   g215(.a(\a[30] ), .b(\b[29] ), .c(new_n304), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n311), .o1(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[30] ), .b(\a[31] ), .out0(new_n313));
  tech160nm_fiaoi012aa1n03p5x5 g218(.a(new_n313), .b(new_n310), .c(new_n312), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  nona22aa1n02x5               g220(.a(new_n310), .b(new_n311), .c(new_n315), .out0(new_n316));
  norb02aa1n03x4               g221(.a(new_n316), .b(new_n314), .out0(\s[31] ));
  xnrb03aa1n02x5               g222(.a(new_n158), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g223(.a(\a[3] ), .b(\b[2] ), .c(new_n158), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g225(.a(new_n160), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  orn002aa1n02x5               g226(.a(\a[6] ), .b(\b[5] ), .o(new_n322));
  oaoi03aa1n02x5               g227(.a(new_n115), .b(new_n116), .c(new_n160), .o1(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n323), .b(new_n108), .c(new_n322), .out0(\s[6] ));
  nano22aa1n02x4               g229(.a(new_n323), .b(new_n108), .c(new_n322), .out0(new_n325));
  aoi013aa1n02x4               g230(.a(new_n123), .b(new_n160), .c(new_n117), .d(new_n118), .o1(new_n326));
  oaib12aa1n02x5               g231(.a(new_n322), .b(new_n109), .c(new_n110), .out0(new_n327));
  oa0022aa1n02x5               g232(.a(new_n325), .b(new_n327), .c(new_n111), .d(new_n326), .o(\s[7] ));
  oai022aa1n02x5               g233(.a(new_n326), .b(new_n111), .c(\b[6] ), .d(\a[7] ), .o1(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g235(.a(new_n162), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


