// Benchmark "adder" written by ABC on Wed Jul 17 13:52:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n332, new_n333, new_n334, new_n336, new_n337, new_n338, new_n339,
    new_n341, new_n342, new_n343, new_n345, new_n346, new_n348, new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  orn002aa1n03x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nanp02aa1n06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n12x5               g005(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(new_n101));
  inv040aa1d32x5               g006(.a(\a[3] ), .o1(new_n102));
  inv040aa1d30x5               g007(.a(\b[2] ), .o1(new_n103));
  nand02aa1n04x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand22aa1n03x5               g010(.a(new_n104), .b(new_n105), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\a[4] ), .o1(new_n107));
  aboi22aa1n03x5               g012(.a(\b[3] ), .b(new_n107), .c(new_n102), .d(new_n103), .out0(new_n108));
  aoai13aa1n06x5               g013(.a(new_n108), .b(new_n106), .c(new_n101), .d(new_n99), .o1(new_n109));
  and002aa1n02x5               g014(.a(\b[4] ), .b(\a[5] ), .o(new_n110));
  oai022aa1n09x5               g015(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n111));
  norp02aa1n02x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[3] ), .o1(new_n113));
  oai022aa1n02x5               g018(.a(new_n107), .b(new_n113), .c(\b[7] ), .d(\a[8] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  oai012aa1n02x5               g020(.a(new_n115), .b(\b[6] ), .c(\a[7] ), .o1(new_n116));
  aoi022aa1n02x7               g021(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n117));
  norb03aa1n03x5               g022(.a(new_n117), .b(new_n114), .c(new_n116), .out0(new_n118));
  nanp03aa1n09x5               g023(.a(new_n109), .b(new_n112), .c(new_n118), .o1(new_n119));
  nor042aa1d18x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  and002aa1n02x7               g025(.a(\b[6] ), .b(\a[7] ), .o(new_n121));
  aoi112aa1n03x5               g026(.a(new_n121), .b(new_n120), .c(\a[6] ), .d(\b[5] ), .o1(new_n122));
  tech160nm_fixorc02aa1n05x5   g027(.a(\a[8] ), .b(\b[7] ), .out0(new_n123));
  inv000aa1d42x5               g028(.a(new_n120), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n122), .c(new_n123), .d(new_n111), .o1(new_n126));
  nanp02aa1n06x5               g031(.a(new_n119), .b(new_n126), .o1(new_n127));
  xnrc02aa1n12x5               g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(new_n127), .b(new_n129), .o1(new_n130));
  xnrc02aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  aoai13aa1n06x5               g038(.a(new_n132), .b(new_n97), .c(new_n127), .d(new_n129), .o1(new_n134));
  nand02aa1n04x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  oai022aa1d18x5               g040(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  norp02aa1n24x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand02aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n06x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n134), .c(new_n137), .out0(\s[11] ));
  aob012aa1n03x5               g046(.a(new_n140), .b(new_n134), .c(new_n137), .out0(new_n142));
  nor002aa1n20x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand22aa1n09x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  norp02aa1n02x5               g050(.a(new_n145), .b(new_n138), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n138), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n140), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n147), .b(new_n148), .c(new_n134), .d(new_n137), .o1(new_n149));
  aoi022aa1n03x5               g054(.a(new_n149), .b(new_n145), .c(new_n142), .d(new_n146), .o1(\s[12] ));
  nona23aa1n09x5               g055(.a(new_n144), .b(new_n139), .c(new_n138), .d(new_n143), .out0(new_n151));
  nona32aa1n02x4               g056(.a(new_n127), .b(new_n151), .c(new_n131), .d(new_n128), .out0(new_n152));
  nona23aa1n02x4               g057(.a(new_n140), .b(new_n145), .c(new_n131), .d(new_n128), .out0(new_n153));
  nanb03aa1n12x5               g058(.a(new_n143), .b(new_n144), .c(new_n139), .out0(new_n154));
  oai112aa1n06x5               g059(.a(new_n136), .b(new_n135), .c(\b[10] ), .d(\a[11] ), .o1(new_n155));
  aoi012aa1n12x5               g060(.a(new_n143), .b(new_n138), .c(new_n144), .o1(new_n156));
  oai012aa1d24x5               g061(.a(new_n156), .b(new_n155), .c(new_n154), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n153), .c(new_n119), .d(new_n126), .o1(new_n159));
  nor042aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand22aa1n04x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  oaib12aa1n02x5               g067(.a(new_n156), .b(new_n160), .c(new_n161), .out0(new_n163));
  oab012aa1n02x4               g068(.a(new_n163), .b(new_n155), .c(new_n154), .out0(new_n164));
  aoi022aa1n02x5               g069(.a(new_n164), .b(new_n152), .c(new_n159), .d(new_n162), .o1(\s[13] ));
  norp02aa1n12x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanp02aa1n04x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoi112aa1n02x5               g073(.a(new_n160), .b(new_n168), .c(new_n159), .d(new_n162), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n168), .b(new_n160), .c(new_n159), .d(new_n161), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(\s[14] ));
  nano23aa1n02x4               g076(.a(new_n160), .b(new_n166), .c(new_n167), .d(new_n161), .out0(new_n172));
  oa0012aa1n02x5               g077(.a(new_n167), .b(new_n166), .c(new_n160), .o(new_n173));
  norp02aa1n09x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nand42aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  aoai13aa1n03x5               g081(.a(new_n176), .b(new_n173), .c(new_n159), .d(new_n172), .o1(new_n177));
  aoi112aa1n02x5               g082(.a(new_n176), .b(new_n173), .c(new_n159), .d(new_n172), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(\s[15] ));
  norp02aa1n12x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nand22aa1n03x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n181), .b(new_n180), .out0(new_n182));
  norp02aa1n02x5               g087(.a(new_n182), .b(new_n174), .o1(new_n183));
  oai012aa1n02x7               g088(.a(new_n177), .b(\b[14] ), .c(\a[15] ), .o1(new_n184));
  aoi022aa1n02x5               g089(.a(new_n184), .b(new_n182), .c(new_n177), .d(new_n183), .o1(\s[16] ));
  nona23aa1n09x5               g090(.a(new_n167), .b(new_n161), .c(new_n160), .d(new_n166), .out0(new_n186));
  nona23aa1n06x5               g091(.a(new_n181), .b(new_n175), .c(new_n174), .d(new_n180), .out0(new_n187));
  nor042aa1n06x5               g092(.a(new_n187), .b(new_n186), .o1(new_n188));
  nona32aa1d24x5               g093(.a(new_n188), .b(new_n151), .c(new_n131), .d(new_n128), .out0(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n127), .b(new_n190), .o1(new_n191));
  nanb03aa1n02x5               g096(.a(new_n180), .b(new_n181), .c(new_n175), .out0(new_n192));
  oai122aa1n02x7               g097(.a(new_n167), .b(new_n166), .c(new_n160), .d(\b[14] ), .e(\a[15] ), .o1(new_n193));
  aoi012aa1n02x5               g098(.a(new_n180), .b(new_n174), .c(new_n181), .o1(new_n194));
  oai012aa1n03x5               g099(.a(new_n194), .b(new_n193), .c(new_n192), .o1(new_n195));
  aoi012aa1n09x5               g100(.a(new_n195), .b(new_n157), .c(new_n188), .o1(new_n196));
  aoai13aa1n12x5               g101(.a(new_n196), .b(new_n189), .c(new_n119), .d(new_n126), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  norp02aa1n02x5               g103(.a(new_n193), .b(new_n192), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n194), .out0(new_n200));
  aoi112aa1n02x5               g105(.a(new_n200), .b(new_n199), .c(new_n157), .d(new_n188), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n197), .b(new_n198), .c(new_n191), .d(new_n201), .o1(\s[17] ));
  nor022aa1n04x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  tech160nm_fixorc02aa1n05x5   g108(.a(\a[18] ), .b(\b[17] ), .out0(new_n204));
  aoi112aa1n02x5               g109(.a(new_n203), .b(new_n204), .c(new_n197), .d(new_n198), .o1(new_n205));
  aoai13aa1n02x5               g110(.a(new_n204), .b(new_n203), .c(new_n197), .d(new_n198), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(\s[18] ));
  and002aa1n06x5               g112(.a(new_n204), .b(new_n198), .o(new_n208));
  nanp02aa1n02x5               g113(.a(new_n197), .b(new_n208), .o1(new_n209));
  inv000aa1d42x5               g114(.a(\a[18] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(\b[17] ), .o1(new_n211));
  oaoi03aa1n02x5               g116(.a(new_n210), .b(new_n211), .c(new_n203), .o1(new_n212));
  tech160nm_fixorc02aa1n04x5   g117(.a(\a[19] ), .b(\b[18] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g120(.a(new_n213), .b(new_n209), .c(new_n212), .out0(new_n216));
  norp02aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  and002aa1n12x5               g122(.a(\b[19] ), .b(\a[20] ), .o(new_n218));
  nor002aa1n02x5               g123(.a(new_n218), .b(new_n217), .o1(new_n219));
  norp02aa1n02x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  oab012aa1n02x4               g125(.a(new_n220), .b(new_n218), .c(new_n217), .out0(new_n221));
  aobi12aa1n02x5               g126(.a(new_n212), .b(new_n197), .c(new_n208), .out0(new_n222));
  oaoi03aa1n02x5               g127(.a(\a[19] ), .b(\b[18] ), .c(new_n222), .o1(new_n223));
  aoi022aa1n02x5               g128(.a(new_n223), .b(new_n219), .c(new_n216), .d(new_n221), .o1(\s[20] ));
  nand23aa1n04x5               g129(.a(new_n208), .b(new_n213), .c(new_n219), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoi012aa1n02x5               g131(.a(new_n203), .b(new_n210), .c(new_n211), .o1(new_n227));
  aoi112aa1n03x5               g132(.a(new_n218), .b(new_n217), .c(\a[19] ), .d(\b[18] ), .o1(new_n228));
  oai022aa1n02x5               g133(.a(new_n210), .b(new_n211), .c(\b[18] ), .d(\a[19] ), .o1(new_n229));
  nona22aa1n09x5               g134(.a(new_n228), .b(new_n229), .c(new_n227), .out0(new_n230));
  aoib12aa1n06x5               g135(.a(new_n217), .b(new_n220), .c(new_n218), .out0(new_n231));
  nanp02aa1n02x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  xorc02aa1n12x5               g137(.a(\a[21] ), .b(\b[20] ), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n232), .c(new_n197), .d(new_n226), .o1(new_n234));
  nano22aa1n02x4               g139(.a(new_n233), .b(new_n230), .c(new_n231), .out0(new_n235));
  aobi12aa1n02x5               g140(.a(new_n235), .b(new_n197), .c(new_n226), .out0(new_n236));
  norb02aa1n02x5               g141(.a(new_n234), .b(new_n236), .out0(\s[21] ));
  xorc02aa1n12x5               g142(.a(\a[22] ), .b(\b[21] ), .out0(new_n238));
  nor042aa1n03x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  norp02aa1n02x5               g144(.a(new_n238), .b(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(\a[21] ), .o1(new_n241));
  oaib12aa1n06x5               g146(.a(new_n234), .b(\b[20] ), .c(new_n241), .out0(new_n242));
  aoi022aa1n02x7               g147(.a(new_n242), .b(new_n238), .c(new_n234), .d(new_n240), .o1(\s[22] ));
  nand02aa1d06x5               g148(.a(new_n238), .b(new_n233), .o1(new_n244));
  nano32aa1n02x4               g149(.a(new_n244), .b(new_n208), .c(new_n213), .d(new_n219), .out0(new_n245));
  inv000aa1d42x5               g150(.a(new_n239), .o1(new_n246));
  oao003aa1n02x5               g151(.a(\a[22] ), .b(\b[21] ), .c(new_n246), .carry(new_n247));
  aoai13aa1n04x5               g152(.a(new_n247), .b(new_n244), .c(new_n230), .d(new_n231), .o1(new_n248));
  xorc02aa1n02x5               g153(.a(\a[23] ), .b(\b[22] ), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n248), .c(new_n197), .d(new_n245), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n244), .o1(new_n251));
  nanb02aa1n02x5               g156(.a(new_n249), .b(new_n247), .out0(new_n252));
  aoi012aa1n02x5               g157(.a(new_n252), .b(new_n232), .c(new_n251), .o1(new_n253));
  aobi12aa1n02x5               g158(.a(new_n253), .b(new_n197), .c(new_n245), .out0(new_n254));
  norb02aa1n02x5               g159(.a(new_n250), .b(new_n254), .out0(\s[23] ));
  xorc02aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  norp02aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  norp02aa1n02x5               g162(.a(new_n256), .b(new_n257), .o1(new_n258));
  tech160nm_fioai012aa1n03p5x5 g163(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .o1(new_n259));
  aoi022aa1n02x5               g164(.a(new_n259), .b(new_n256), .c(new_n250), .d(new_n258), .o1(\s[24] ));
  and002aa1n02x5               g165(.a(new_n256), .b(new_n249), .o(new_n261));
  nano22aa1n03x7               g166(.a(new_n225), .b(new_n261), .c(new_n251), .out0(new_n262));
  inv000aa1d42x5               g167(.a(\a[24] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(\b[23] ), .o1(new_n264));
  tech160nm_fioaoi03aa1n02p5x5 g169(.a(new_n263), .b(new_n264), .c(new_n257), .o1(new_n265));
  aob012aa1n02x5               g170(.a(new_n265), .b(new_n248), .c(new_n261), .out0(new_n266));
  xorc02aa1n02x5               g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n266), .c(new_n197), .d(new_n262), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n265), .o1(new_n269));
  aoi112aa1n02x5               g174(.a(new_n267), .b(new_n269), .c(new_n248), .d(new_n261), .o1(new_n270));
  aobi12aa1n02x5               g175(.a(new_n270), .b(new_n262), .c(new_n197), .out0(new_n271));
  norb02aa1n03x4               g176(.a(new_n268), .b(new_n271), .out0(\s[25] ));
  xorc02aa1n02x5               g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  norp02aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  norp02aa1n02x5               g179(.a(new_n273), .b(new_n274), .o1(new_n275));
  inv000aa1d42x5               g180(.a(\a[25] ), .o1(new_n276));
  oaib12aa1n06x5               g181(.a(new_n268), .b(\b[24] ), .c(new_n276), .out0(new_n277));
  aoi022aa1n02x7               g182(.a(new_n277), .b(new_n273), .c(new_n268), .d(new_n275), .o1(\s[26] ));
  inv000aa1d42x5               g183(.a(\a[26] ), .o1(new_n279));
  xroi22aa1d04x5               g184(.a(new_n276), .b(\b[24] ), .c(new_n279), .d(\b[25] ), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n269), .c(new_n248), .d(new_n261), .o1(new_n281));
  nano32aa1n03x7               g186(.a(new_n225), .b(new_n280), .c(new_n251), .d(new_n261), .out0(new_n282));
  nand22aa1n03x5               g187(.a(new_n197), .b(new_n282), .o1(new_n283));
  inv000aa1d42x5               g188(.a(\b[25] ), .o1(new_n284));
  oaoi03aa1n02x5               g189(.a(new_n279), .b(new_n284), .c(new_n274), .o1(new_n285));
  nand23aa1n04x5               g190(.a(new_n283), .b(new_n281), .c(new_n285), .o1(new_n286));
  xorc02aa1n02x5               g191(.a(\a[27] ), .b(\b[26] ), .out0(new_n287));
  inv000aa1n02x5               g192(.a(new_n285), .o1(new_n288));
  aoi112aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n197), .d(new_n282), .o1(new_n289));
  aoi022aa1n02x5               g194(.a(new_n286), .b(new_n287), .c(new_n289), .d(new_n281), .o1(\s[27] ));
  nanp02aa1n03x5               g195(.a(new_n286), .b(new_n287), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[28] ), .b(\b[27] ), .out0(new_n292));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  norp02aa1n02x5               g198(.a(new_n292), .b(new_n293), .o1(new_n294));
  tech160nm_fiaoi012aa1n05x5   g199(.a(new_n288), .b(new_n197), .c(new_n282), .o1(new_n295));
  inv000aa1n03x5               g200(.a(new_n293), .o1(new_n296));
  inv030aa1n02x5               g201(.a(new_n287), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n296), .b(new_n297), .c(new_n295), .d(new_n281), .o1(new_n298));
  aoi022aa1n03x5               g203(.a(new_n298), .b(new_n292), .c(new_n291), .d(new_n294), .o1(\s[28] ));
  and002aa1n02x5               g204(.a(new_n292), .b(new_n287), .o(new_n300));
  nanp02aa1n03x5               g205(.a(new_n286), .b(new_n300), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[29] ), .b(\b[28] ), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n296), .carry(new_n303));
  norb02aa1n02x5               g208(.a(new_n303), .b(new_n302), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n300), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n303), .b(new_n305), .c(new_n295), .d(new_n281), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g213(.a(new_n292), .b(new_n287), .c(new_n302), .o1(new_n309));
  nanb02aa1n06x5               g214(.a(new_n309), .b(new_n286), .out0(new_n310));
  xorc02aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .out0(new_n311));
  inv000aa1d42x5               g216(.a(\a[29] ), .o1(new_n312));
  inv000aa1d42x5               g217(.a(\b[28] ), .o1(new_n313));
  oaib12aa1n02x5               g218(.a(new_n303), .b(\b[28] ), .c(new_n312), .out0(new_n314));
  oaoi13aa1n04x5               g219(.a(new_n311), .b(new_n314), .c(new_n312), .d(new_n313), .o1(new_n315));
  oaib12aa1n02x5               g220(.a(new_n314), .b(new_n313), .c(\a[29] ), .out0(new_n316));
  aoai13aa1n02x7               g221(.a(new_n316), .b(new_n309), .c(new_n295), .d(new_n281), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n311), .c(new_n310), .d(new_n315), .o1(\s[30] ));
  nano32aa1n02x4               g223(.a(new_n297), .b(new_n311), .c(new_n292), .d(new_n302), .out0(new_n319));
  nanp02aa1n03x5               g224(.a(new_n286), .b(new_n319), .o1(new_n320));
  aoi022aa1n02x5               g225(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n321));
  norb02aa1n02x5               g226(.a(\b[30] ), .b(\a[31] ), .out0(new_n322));
  obai22aa1n02x7               g227(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n323));
  aoi112aa1n02x5               g228(.a(new_n323), .b(new_n322), .c(new_n314), .d(new_n321), .o1(new_n324));
  inv000aa1n02x5               g229(.a(new_n319), .o1(new_n325));
  norp02aa1n02x5               g230(.a(\b[29] ), .b(\a[30] ), .o1(new_n326));
  aoi012aa1n02x5               g231(.a(new_n326), .b(new_n314), .c(new_n321), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n325), .c(new_n295), .d(new_n281), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n328), .b(new_n329), .c(new_n324), .d(new_n320), .o1(\s[31] ));
  xobna2aa1n03x5               g235(.a(new_n106), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  nanp02aa1n02x5               g236(.a(new_n101), .b(new_n99), .o1(new_n332));
  nanp03aa1n02x5               g237(.a(new_n332), .b(new_n104), .c(new_n105), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[4] ), .b(\b[3] ), .out0(new_n334));
  xnbna2aa1n03x5               g239(.a(new_n334), .b(new_n333), .c(new_n104), .out0(\s[4] ));
  norp02aa1n02x5               g240(.a(\b[4] ), .b(\a[5] ), .o1(new_n336));
  aoi112aa1n02x5               g241(.a(new_n110), .b(new_n336), .c(\a[4] ), .d(\b[3] ), .o1(new_n337));
  oaib12aa1n02x5               g242(.a(new_n109), .b(new_n113), .c(\a[4] ), .out0(new_n338));
  xnrc02aa1n02x5               g243(.a(\b[4] ), .b(\a[5] ), .out0(new_n339));
  aoi022aa1n02x5               g244(.a(new_n338), .b(new_n339), .c(new_n337), .d(new_n109), .o1(\s[5] ));
  xorc02aa1n02x5               g245(.a(\a[6] ), .b(\b[5] ), .out0(new_n341));
  aoai13aa1n02x5               g246(.a(new_n341), .b(new_n336), .c(new_n109), .d(new_n337), .o1(new_n342));
  aoi112aa1n02x5               g247(.a(new_n336), .b(new_n341), .c(new_n109), .d(new_n337), .o1(new_n343));
  norb02aa1n02x5               g248(.a(new_n342), .b(new_n343), .out0(\s[6] ));
  orn002aa1n02x5               g249(.a(\a[6] ), .b(\b[5] ), .o(new_n345));
  norp02aa1n02x5               g250(.a(new_n121), .b(new_n120), .o1(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n342), .c(new_n345), .out0(\s[7] ));
  aob012aa1n02x5               g252(.a(new_n346), .b(new_n342), .c(new_n345), .out0(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n123), .b(new_n348), .c(new_n124), .out0(\s[8] ));
  aoi113aa1n02x5               g254(.a(new_n129), .b(new_n125), .c(new_n122), .d(new_n123), .e(new_n111), .o1(new_n350));
  aoi022aa1n02x5               g255(.a(new_n127), .b(new_n129), .c(new_n119), .d(new_n350), .o1(\s[9] ));
endmodule


