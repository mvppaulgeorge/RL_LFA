// Benchmark "adder" written by ABC on Thu Jul 18 02:33:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n330, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor042aa1d18x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  tech160nm_fixnrc02aa1n03p5x5 g006(.a(\b[7] ), .b(\a[8] ), .out0(new_n102));
  nor002aa1d24x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nanb02aa1n03x5               g009(.a(new_n103), .b(new_n104), .out0(new_n105));
  nanp02aa1n02x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor022aa1n04x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nor042aa1n04x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  oaih12aa1n02x5               g013(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n109));
  inv000aa1d42x5               g014(.a(new_n103), .o1(new_n110));
  oao003aa1n02x5               g015(.a(\a[8] ), .b(\b[7] ), .c(new_n110), .carry(new_n111));
  oai013aa1n03x5               g016(.a(new_n111), .b(new_n102), .c(new_n109), .d(new_n105), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  nor042aa1n04x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  nand02aa1n03x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  tech160nm_fiaoi012aa1n03p5x5 g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  nand22aa1n03x5               g022(.a(\b[0] ), .b(\a[1] ), .o1(new_n118));
  nor042aa1n03x5               g023(.a(\b[1] ), .b(\a[2] ), .o1(new_n119));
  tech160nm_fioai012aa1n03p5x5 g024(.a(new_n117), .b(new_n119), .c(new_n118), .o1(new_n120));
  nanp02aa1n03x5               g025(.a(\b[2] ), .b(\a[3] ), .o1(new_n121));
  nona23aa1n09x5               g026(.a(new_n115), .b(new_n121), .c(new_n114), .d(new_n113), .out0(new_n122));
  oai012aa1n09x5               g027(.a(new_n116), .b(new_n122), .c(new_n120), .o1(new_n123));
  nanb02aa1n02x5               g028(.a(new_n107), .b(new_n106), .out0(new_n124));
  nanp02aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  nona23aa1n02x5               g030(.a(new_n125), .b(new_n104), .c(new_n103), .d(new_n108), .out0(new_n126));
  nor043aa1n03x5               g031(.a(new_n126), .b(new_n124), .c(new_n102), .o1(new_n127));
  nand42aa1n16x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n03x5               g034(.a(new_n129), .b(new_n112), .c(new_n123), .d(new_n127), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  inv040aa1d32x5               g036(.a(\a[11] ), .o1(new_n132));
  inv040aa1n20x5               g037(.a(\b[10] ), .o1(new_n133));
  nand22aa1n04x5               g038(.a(new_n133), .b(new_n132), .o1(new_n134));
  nand22aa1n09x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand22aa1n02x5               g040(.a(new_n134), .b(new_n135), .o1(new_n136));
  nona22aa1n02x4               g041(.a(new_n130), .b(new_n100), .c(new_n97), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n136), .b(new_n137), .c(new_n98), .out0(\s[11] ));
  inv040aa1d32x5               g043(.a(\a[12] ), .o1(new_n139));
  inv040aa1d28x5               g044(.a(\b[11] ), .o1(new_n140));
  nanp02aa1n06x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  nand42aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norp02aa1n04x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  aoi013aa1n03x5               g048(.a(new_n143), .b(new_n137), .c(new_n135), .d(new_n98), .o1(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n141), .c(new_n142), .out0(\s[12] ));
  tech160nm_fiaoi012aa1n05x5   g050(.a(new_n112), .b(new_n123), .c(new_n127), .o1(new_n146));
  nand02aa1n03x5               g051(.a(new_n141), .b(new_n142), .o1(new_n147));
  nano23aa1d15x5               g052(.a(new_n97), .b(new_n100), .c(new_n128), .d(new_n98), .out0(new_n148));
  nona22aa1d24x5               g053(.a(new_n148), .b(new_n147), .c(new_n136), .out0(new_n149));
  nanb03aa1n03x5               g054(.a(new_n143), .b(new_n135), .c(new_n98), .out0(new_n150));
  oai112aa1n06x5               g055(.a(new_n141), .b(new_n142), .c(new_n100), .d(new_n97), .o1(new_n151));
  oaoi03aa1n02x5               g056(.a(new_n139), .b(new_n140), .c(new_n143), .o1(new_n152));
  oaih12aa1n02x5               g057(.a(new_n152), .b(new_n151), .c(new_n150), .o1(new_n153));
  oabi12aa1n02x5               g058(.a(new_n153), .b(new_n146), .c(new_n149), .out0(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1n06x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n156), .b(new_n154), .c(new_n157), .o1(new_n158));
  xnrb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n03x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nano23aa1n06x5               g066(.a(new_n156), .b(new_n160), .c(new_n161), .d(new_n157), .out0(new_n162));
  oa0012aa1n02x5               g067(.a(new_n161), .b(new_n160), .c(new_n156), .o(new_n163));
  aoi012aa1n02x5               g068(.a(new_n163), .b(new_n153), .c(new_n162), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n149), .o1(new_n165));
  nano22aa1n03x7               g070(.a(new_n146), .b(new_n165), .c(new_n162), .out0(new_n166));
  nor042aa1n09x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n02x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  oaib12aa1n06x5               g074(.a(new_n169), .b(new_n166), .c(new_n164), .out0(new_n170));
  norb03aa1n02x5               g075(.a(new_n164), .b(new_n166), .c(new_n169), .out0(new_n171));
  norb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(\s[15] ));
  inv000aa1d42x5               g077(.a(new_n167), .o1(new_n173));
  nor042aa1n03x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1n06x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n170), .c(new_n173), .out0(\s[16] ));
  nano23aa1n06x5               g082(.a(new_n167), .b(new_n174), .c(new_n175), .d(new_n168), .out0(new_n178));
  nano22aa1n03x7               g083(.a(new_n149), .b(new_n162), .c(new_n178), .out0(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n112), .c(new_n123), .d(new_n127), .o1(new_n180));
  aoai13aa1n06x5               g085(.a(new_n178), .b(new_n163), .c(new_n153), .d(new_n162), .o1(new_n181));
  aoi012aa1d18x5               g086(.a(new_n174), .b(new_n167), .c(new_n175), .o1(new_n182));
  nand23aa1n06x5               g087(.a(new_n180), .b(new_n181), .c(new_n182), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[18] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[17] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[16] ), .o1(new_n187));
  oaoi03aa1n03x5               g092(.a(new_n186), .b(new_n187), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  nona23aa1n02x4               g094(.a(new_n161), .b(new_n157), .c(new_n156), .d(new_n160), .out0(new_n190));
  oaoi13aa1n06x5               g095(.a(new_n190), .b(new_n152), .c(new_n151), .d(new_n150), .o1(new_n191));
  inv000aa1n02x5               g096(.a(new_n182), .o1(new_n192));
  oaoi13aa1n04x5               g097(.a(new_n192), .b(new_n178), .c(new_n191), .d(new_n163), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n186), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n194));
  inv030aa1n03x5               g099(.a(new_n194), .o1(new_n195));
  inv000aa1d42x5               g100(.a(\b[17] ), .o1(new_n196));
  oai022aa1d24x5               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oa0012aa1n02x5               g102(.a(new_n197), .b(new_n196), .c(new_n185), .o(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  aoai13aa1n02x7               g104(.a(new_n199), .b(new_n195), .c(new_n193), .d(new_n180), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g106(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g107(.a(\a[19] ), .o1(new_n203));
  inv040aa1d28x5               g108(.a(\b[18] ), .o1(new_n204));
  nand22aa1n09x5               g109(.a(new_n204), .b(new_n203), .o1(new_n205));
  tech160nm_fixorc02aa1n03p5x5 g110(.a(\a[19] ), .b(\b[18] ), .out0(new_n206));
  aoai13aa1n03x5               g111(.a(new_n206), .b(new_n198), .c(new_n183), .d(new_n194), .o1(new_n207));
  xorc02aa1n12x5               g112(.a(\a[20] ), .b(\b[19] ), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  tech160nm_fiaoi012aa1n02p5x5 g114(.a(new_n209), .b(new_n207), .c(new_n205), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n205), .o1(new_n211));
  aoi112aa1n02x5               g116(.a(new_n211), .b(new_n208), .c(new_n200), .d(new_n206), .o1(new_n212));
  nor002aa1n02x5               g117(.a(new_n210), .b(new_n212), .o1(\s[20] ));
  nano22aa1n12x5               g118(.a(new_n195), .b(new_n206), .c(new_n208), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  and002aa1n02x5               g120(.a(\b[19] ), .b(\a[20] ), .o(new_n216));
  oai122aa1n06x5               g121(.a(new_n197), .b(new_n203), .c(new_n204), .d(new_n185), .e(new_n196), .o1(new_n217));
  oai112aa1n06x5               g122(.a(new_n217), .b(new_n205), .c(\b[19] ), .d(\a[20] ), .o1(new_n218));
  norb02aa1n15x5               g123(.a(new_n218), .b(new_n216), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n02x7               g125(.a(new_n220), .b(new_n215), .c(new_n193), .d(new_n180), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  nand42aa1n03x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  norb02aa1n02x5               g130(.a(new_n225), .b(new_n223), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n219), .c(new_n183), .d(new_n214), .o1(new_n227));
  nor042aa1n06x5               g132(.a(\b[21] ), .b(\a[22] ), .o1(new_n228));
  nand42aa1n08x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  nanb02aa1d36x5               g134(.a(new_n228), .b(new_n229), .out0(new_n230));
  aoi012aa1n02x7               g135(.a(new_n230), .b(new_n227), .c(new_n224), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n230), .o1(new_n232));
  aoi112aa1n02x5               g137(.a(new_n223), .b(new_n232), .c(new_n221), .d(new_n225), .o1(new_n233));
  nor002aa1n02x5               g138(.a(new_n231), .b(new_n233), .o1(\s[22] ));
  xorc02aa1n02x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  nano23aa1n09x5               g140(.a(new_n223), .b(new_n228), .c(new_n229), .d(new_n225), .out0(new_n236));
  nand23aa1n04x5               g141(.a(new_n183), .b(new_n214), .c(new_n236), .o1(new_n237));
  tech160nm_fioai012aa1n05x5   g142(.a(new_n229), .b(new_n228), .c(new_n223), .o1(new_n238));
  aob012aa1n02x5               g143(.a(new_n238), .b(new_n219), .c(new_n236), .out0(new_n239));
  norb02aa1n03x5               g144(.a(new_n235), .b(new_n239), .out0(new_n240));
  tech160nm_finand02aa1n03p5x5 g145(.a(new_n237), .b(new_n240), .o1(new_n241));
  aoi013aa1n02x4               g146(.a(new_n239), .b(new_n183), .c(new_n214), .d(new_n236), .o1(new_n242));
  oai012aa1n02x5               g147(.a(new_n241), .b(new_n242), .c(new_n235), .o1(\s[23] ));
  and002aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o(new_n244));
  xorc02aa1n02x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoai13aa1n02x7               g150(.a(new_n245), .b(new_n244), .c(new_n237), .d(new_n240), .o1(new_n246));
  nona22aa1n03x5               g151(.a(new_n241), .b(new_n245), .c(new_n244), .out0(new_n247));
  nanp02aa1n03x5               g152(.a(new_n247), .b(new_n246), .o1(\s[24] ));
  inv000aa1d42x5               g153(.a(\a[23] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\b[22] ), .o1(new_n250));
  nand42aa1n02x5               g155(.a(new_n250), .b(new_n249), .o1(new_n251));
  nand42aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  orn002aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .o(new_n253));
  oai112aa1n06x5               g158(.a(new_n253), .b(new_n252), .c(new_n250), .d(new_n249), .o1(new_n254));
  nano22aa1n06x5               g159(.a(new_n254), .b(new_n236), .c(new_n251), .out0(new_n255));
  inv000aa1n06x5               g160(.a(new_n255), .o1(new_n256));
  nano32aa1n03x7               g161(.a(new_n256), .b(new_n194), .c(new_n206), .d(new_n208), .out0(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  aoi112aa1n03x5               g163(.a(new_n254), .b(new_n238), .c(new_n249), .d(new_n250), .o1(new_n259));
  oaoi03aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .o1(new_n260));
  nor042aa1n04x5               g165(.a(new_n259), .b(new_n260), .o1(new_n261));
  nano32aa1n03x7               g166(.a(new_n230), .b(new_n224), .c(new_n251), .d(new_n225), .out0(new_n262));
  nona23aa1d18x5               g167(.a(new_n218), .b(new_n262), .c(new_n254), .d(new_n216), .out0(new_n263));
  nand22aa1n12x5               g168(.a(new_n263), .b(new_n261), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  aoai13aa1n02x7               g170(.a(new_n265), .b(new_n258), .c(new_n193), .d(new_n180), .o1(new_n266));
  xorb03aa1n02x5               g171(.a(new_n266), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g172(.a(\b[24] ), .b(\a[25] ), .o1(new_n268));
  inv000aa1n03x5               g173(.a(new_n268), .o1(new_n269));
  xorc02aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n264), .c(new_n183), .d(new_n257), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[26] ), .b(\b[25] ), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  tech160nm_fiaoi012aa1n02p5x5 g178(.a(new_n273), .b(new_n271), .c(new_n269), .o1(new_n274));
  aoi112aa1n02x5               g179(.a(new_n268), .b(new_n272), .c(new_n266), .d(new_n270), .o1(new_n275));
  nor002aa1n02x5               g180(.a(new_n274), .b(new_n275), .o1(\s[26] ));
  and002aa1n12x5               g181(.a(new_n272), .b(new_n270), .o(new_n277));
  nand23aa1n03x5               g182(.a(new_n214), .b(new_n255), .c(new_n277), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .c(new_n269), .carry(new_n279));
  inv000aa1n02x5               g184(.a(new_n279), .o1(new_n280));
  tech160nm_fiaoi012aa1n05x5   g185(.a(new_n280), .b(new_n264), .c(new_n277), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n281), .b(new_n278), .c(new_n193), .d(new_n180), .o1(new_n282));
  xorb03aa1n02x5               g187(.a(new_n282), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[28] ), .b(\b[27] ), .out0(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n278), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n277), .o1(new_n290));
  aoai13aa1n12x5               g195(.a(new_n279), .b(new_n290), .c(new_n263), .d(new_n261), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n288), .b(new_n291), .c(new_n183), .d(new_n289), .o1(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n287), .b(new_n292), .c(new_n285), .o1(new_n293));
  aoi112aa1n03x4               g198(.a(new_n286), .b(new_n284), .c(new_n282), .d(new_n288), .o1(new_n294));
  nor002aa1n02x5               g199(.a(new_n293), .b(new_n294), .o1(\s[28] ));
  nano22aa1n02x4               g200(.a(new_n287), .b(new_n285), .c(new_n288), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n291), .c(new_n183), .d(new_n289), .o1(new_n297));
  oao003aa1n09x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n298));
  xorc02aa1n12x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n297), .c(new_n298), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n298), .o1(new_n302));
  aoi112aa1n03x4               g207(.a(new_n299), .b(new_n302), .c(new_n282), .d(new_n296), .o1(new_n303));
  nor002aa1n02x5               g208(.a(new_n301), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n118), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g210(.a(new_n300), .b(new_n286), .c(new_n288), .d(new_n285), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n291), .c(new_n183), .d(new_n289), .o1(new_n307));
  oao003aa1n09x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n308));
  xorc02aa1n12x5               g213(.a(\a[30] ), .b(\b[29] ), .out0(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n310), .b(new_n307), .c(new_n308), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n308), .o1(new_n312));
  aoi112aa1n03x4               g217(.a(new_n309), .b(new_n312), .c(new_n282), .d(new_n306), .o1(new_n313));
  nor002aa1n02x5               g218(.a(new_n311), .b(new_n313), .o1(\s[30] ));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  and003aa1n02x5               g220(.a(new_n296), .b(new_n309), .c(new_n299), .o(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n291), .c(new_n183), .d(new_n289), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n318));
  aoi012aa1n03x5               g223(.a(new_n315), .b(new_n317), .c(new_n318), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n315), .o1(new_n320));
  inv000aa1n02x5               g225(.a(new_n318), .o1(new_n321));
  aoi112aa1n02x5               g226(.a(new_n320), .b(new_n321), .c(new_n282), .d(new_n316), .o1(new_n322));
  nor002aa1n02x5               g227(.a(new_n319), .b(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n120), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g229(.a(\a[3] ), .b(\b[2] ), .c(new_n120), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n123), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g232(.a(new_n125), .b(new_n123), .c(new_n108), .o1(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oab012aa1n02x4               g234(.a(new_n107), .b(new_n328), .c(new_n124), .out0(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n330), .b(new_n110), .c(new_n104), .out0(\s[7] ));
  oaoi03aa1n02x5               g236(.a(\a[7] ), .b(\b[6] ), .c(new_n330), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g238(.a(new_n146), .b(new_n128), .c(new_n101), .out0(\s[9] ));
endmodule


