// Benchmark "adder" written by ABC on Thu Jul 18 00:27:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n312, new_n315, new_n317, new_n319;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[3] ), .b(\a[4] ), .out0(new_n97));
  tech160nm_fixnrc02aa1n05x5   g002(.a(\b[2] ), .b(\a[3] ), .out0(new_n98));
  nanp02aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1d12x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai012aa1n12x5               g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\a[3] ), .o1(new_n103));
  nanb02aa1n03x5               g008(.a(\b[2] ), .b(new_n103), .out0(new_n104));
  oao003aa1n03x5               g009(.a(\a[4] ), .b(\b[3] ), .c(new_n104), .carry(new_n105));
  oai013aa1d12x5               g010(.a(new_n105), .b(new_n98), .c(new_n97), .d(new_n102), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nanp02aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor022aa1n16x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nona23aa1d18x5               g015(.a(new_n110), .b(new_n108), .c(new_n107), .d(new_n109), .out0(new_n111));
  xnrc02aa1n02x5               g016(.a(\b[5] ), .b(\a[6] ), .out0(new_n112));
  nor042aa1d18x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanb02aa1n02x5               g019(.a(new_n113), .b(new_n114), .out0(new_n115));
  nor043aa1n06x5               g020(.a(new_n111), .b(new_n112), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[6] ), .o1(new_n117));
  aob012aa1n03x5               g022(.a(new_n113), .b(\b[5] ), .c(\a[6] ), .out0(new_n118));
  oaib12aa1n03x5               g023(.a(new_n118), .b(\b[5] ), .c(new_n117), .out0(new_n119));
  tech160nm_fioai012aa1n02p5x5 g024(.a(new_n108), .b(new_n109), .c(new_n107), .o1(new_n120));
  oaib12aa1n09x5               g025(.a(new_n120), .b(new_n111), .c(new_n119), .out0(new_n121));
  aoi012aa1n03x5               g026(.a(new_n121), .b(new_n106), .c(new_n116), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[9] ), .b(\b[8] ), .c(new_n122), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n04x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nand42aa1d28x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nor042aa1n06x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nand42aa1n04x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nano23aa1d18x5               g033(.a(new_n125), .b(new_n127), .c(new_n128), .d(new_n126), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n121), .c(new_n106), .d(new_n116), .o1(new_n130));
  tech160nm_fiaoi012aa1n05x5   g035(.a(new_n125), .b(new_n127), .c(new_n126), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(new_n130), .b(new_n131), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand02aa1d24x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n134), .b(new_n132), .c(new_n135), .o1(new_n136));
  xnrb03aa1n02x5               g041(.a(new_n136), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv000aa1d42x5               g042(.a(\a[13] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n106), .b(new_n116), .o1(new_n139));
  inv000aa1n02x5               g044(.a(new_n121), .o1(new_n140));
  nanp02aa1n03x5               g045(.a(new_n139), .b(new_n140), .o1(new_n141));
  nor002aa1d32x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d16x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nano23aa1d15x5               g048(.a(new_n134), .b(new_n142), .c(new_n143), .d(new_n135), .out0(new_n144));
  nona23aa1n03x5               g049(.a(new_n143), .b(new_n135), .c(new_n134), .d(new_n142), .out0(new_n145));
  oa0012aa1n03x5               g050(.a(new_n143), .b(new_n142), .c(new_n134), .o(new_n146));
  oabi12aa1n03x5               g051(.a(new_n146), .b(new_n131), .c(new_n145), .out0(new_n147));
  aoi013aa1n03x5               g052(.a(new_n147), .b(new_n141), .c(new_n129), .d(new_n144), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[12] ), .c(new_n138), .out0(\s[13] ));
  nanb02aa1d24x5               g054(.a(\b[12] ), .b(new_n138), .out0(new_n150));
  xnrc02aa1n12x5               g055(.a(\b[12] ), .b(\a[13] ), .out0(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[13] ), .b(\a[14] ), .out0(new_n152));
  oai112aa1n02x5               g057(.a(new_n152), .b(new_n150), .c(new_n148), .d(new_n151), .o1(new_n153));
  oaoi13aa1n02x7               g058(.a(new_n152), .b(new_n150), .c(new_n148), .d(new_n151), .o1(new_n154));
  norb02aa1n03x4               g059(.a(new_n153), .b(new_n154), .out0(\s[14] ));
  xorc02aa1n02x5               g060(.a(\a[15] ), .b(\b[14] ), .out0(new_n156));
  nor042aa1n09x5               g061(.a(new_n152), .b(new_n151), .o1(new_n157));
  nano32aa1n03x7               g062(.a(new_n122), .b(new_n157), .c(new_n129), .d(new_n144), .out0(new_n158));
  inv020aa1n03x5               g063(.a(new_n131), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n157), .b(new_n146), .c(new_n144), .d(new_n159), .o1(new_n160));
  oaoi03aa1n02x5               g065(.a(\a[14] ), .b(\b[13] ), .c(new_n150), .o1(new_n161));
  inv000aa1n02x5               g066(.a(new_n161), .o1(new_n162));
  nand22aa1n03x5               g067(.a(new_n160), .b(new_n162), .o1(new_n163));
  tech160nm_fioai012aa1n05x5   g068(.a(new_n156), .b(new_n158), .c(new_n163), .o1(new_n164));
  norp03aa1n02x5               g069(.a(new_n158), .b(new_n163), .c(new_n156), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(\s[15] ));
  inv040aa1d30x5               g071(.a(\a[15] ), .o1(new_n167));
  inv040aa1d28x5               g072(.a(\b[14] ), .o1(new_n168));
  nand02aa1d24x5               g073(.a(new_n168), .b(new_n167), .o1(new_n169));
  nor002aa1d32x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand02aa1d16x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nanb02aa1d36x5               g076(.a(new_n170), .b(new_n171), .out0(new_n172));
  xobna2aa1n03x5               g077(.a(new_n172), .b(new_n164), .c(new_n169), .out0(\s[16] ));
  nand02aa1d28x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nano22aa1d33x5               g079(.a(new_n172), .b(new_n169), .c(new_n174), .out0(new_n175));
  aoai13aa1n04x5               g080(.a(new_n175), .b(new_n161), .c(new_n147), .d(new_n157), .o1(new_n176));
  aoai13aa1n06x5               g081(.a(new_n171), .b(new_n170), .c(new_n167), .d(new_n168), .o1(new_n177));
  nand22aa1n12x5               g082(.a(new_n175), .b(new_n129), .o1(new_n178));
  nano22aa1d15x5               g083(.a(new_n178), .b(new_n157), .c(new_n144), .out0(new_n179));
  aoai13aa1n12x5               g084(.a(new_n179), .b(new_n121), .c(new_n106), .d(new_n116), .o1(new_n180));
  nand23aa1d12x5               g085(.a(new_n180), .b(new_n176), .c(new_n177), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  nand42aa1d28x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  tech160nm_fioai012aa1n05x5   g089(.a(new_n184), .b(new_n181), .c(new_n183), .o1(new_n185));
  xnrb03aa1n03x5               g090(.a(new_n185), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  aobi12aa1n12x5               g091(.a(new_n177), .b(new_n163), .c(new_n175), .out0(new_n187));
  nor022aa1n16x5               g092(.a(\b[17] ), .b(\a[18] ), .o1(new_n188));
  nand42aa1d28x5               g093(.a(\b[17] ), .b(\a[18] ), .o1(new_n189));
  nano23aa1d15x5               g094(.a(new_n183), .b(new_n188), .c(new_n189), .d(new_n184), .out0(new_n190));
  inv000aa1d42x5               g095(.a(new_n190), .o1(new_n191));
  aoi012aa1d18x5               g096(.a(new_n188), .b(new_n183), .c(new_n189), .o1(new_n192));
  aoai13aa1n04x5               g097(.a(new_n192), .b(new_n191), .c(new_n187), .d(new_n180), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nand02aa1d08x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  nor002aa1d32x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1n08x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1n02x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  aoi112aa1n03x4               g106(.a(new_n196), .b(new_n201), .c(new_n193), .d(new_n198), .o1(new_n202));
  inv040aa1n08x5               g107(.a(new_n196), .o1(new_n203));
  inv020aa1n04x5               g108(.a(new_n192), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n198), .b(new_n204), .c(new_n181), .d(new_n190), .o1(new_n205));
  aobi12aa1n06x5               g110(.a(new_n201), .b(new_n205), .c(new_n203), .out0(new_n206));
  nor002aa1n02x5               g111(.a(new_n206), .b(new_n202), .o1(\s[20] ));
  nano23aa1n09x5               g112(.a(new_n196), .b(new_n199), .c(new_n200), .d(new_n197), .out0(new_n208));
  nand22aa1n09x5               g113(.a(new_n208), .b(new_n190), .o1(new_n209));
  nona23aa1d18x5               g114(.a(new_n200), .b(new_n197), .c(new_n196), .d(new_n199), .out0(new_n210));
  oaoi03aa1n09x5               g115(.a(\a[20] ), .b(\b[19] ), .c(new_n203), .o1(new_n211));
  inv040aa1n03x5               g116(.a(new_n211), .o1(new_n212));
  oai012aa1d24x5               g117(.a(new_n212), .b(new_n210), .c(new_n192), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  aoai13aa1n04x5               g119(.a(new_n214), .b(new_n209), .c(new_n187), .d(new_n180), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xorc02aa1n02x5               g123(.a(\a[22] ), .b(\b[21] ), .out0(new_n219));
  aoi112aa1n02x5               g124(.a(new_n217), .b(new_n219), .c(new_n215), .d(new_n218), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n217), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n209), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n218), .b(new_n213), .c(new_n181), .d(new_n222), .o1(new_n223));
  aobi12aa1n06x5               g128(.a(new_n219), .b(new_n223), .c(new_n221), .out0(new_n224));
  nor002aa1n02x5               g129(.a(new_n224), .b(new_n220), .o1(\s[22] ));
  inv040aa1d30x5               g130(.a(\a[21] ), .o1(new_n226));
  inv040aa1n08x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  oao003aa1n12x5               g133(.a(\a[22] ), .b(\b[21] ), .c(new_n221), .carry(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoi012aa1d18x5               g135(.a(new_n230), .b(new_n213), .c(new_n228), .o1(new_n231));
  nano22aa1n02x5               g136(.a(new_n209), .b(new_n218), .c(new_n219), .out0(new_n232));
  inv000aa1n02x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n04x5               g138(.a(new_n231), .b(new_n233), .c(new_n187), .d(new_n180), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  xorc02aa1n12x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  xorc02aa1n12x5               g142(.a(\a[24] ), .b(\b[23] ), .out0(new_n238));
  aoi112aa1n03x4               g143(.a(new_n236), .b(new_n238), .c(new_n234), .d(new_n237), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n236), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n231), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n237), .b(new_n241), .c(new_n181), .d(new_n232), .o1(new_n242));
  aobi12aa1n06x5               g147(.a(new_n238), .b(new_n242), .c(new_n240), .out0(new_n243));
  nor042aa1n03x5               g148(.a(new_n243), .b(new_n239), .o1(\s[24] ));
  and002aa1n03x5               g149(.a(new_n238), .b(new_n237), .o(new_n245));
  inv030aa1n03x5               g150(.a(new_n245), .o1(new_n246));
  nano32aa1n02x4               g151(.a(new_n246), .b(new_n228), .c(new_n208), .d(new_n190), .out0(new_n247));
  inv000aa1n02x5               g152(.a(new_n247), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n228), .b(new_n211), .c(new_n208), .d(new_n204), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  oai022aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(new_n251), .b(new_n250), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n252), .b(new_n246), .c(new_n249), .d(new_n229), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  aoai13aa1n04x5               g159(.a(new_n254), .b(new_n248), .c(new_n187), .d(new_n180), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  xorc02aa1n12x5               g163(.a(\a[26] ), .b(\b[25] ), .out0(new_n259));
  aoi112aa1n03x4               g164(.a(new_n257), .b(new_n259), .c(new_n255), .d(new_n258), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n257), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n258), .b(new_n253), .c(new_n181), .d(new_n247), .o1(new_n262));
  aobi12aa1n06x5               g167(.a(new_n259), .b(new_n262), .c(new_n261), .out0(new_n263));
  nor002aa1n02x5               g168(.a(new_n263), .b(new_n260), .o1(\s[26] ));
  inv000aa1d42x5               g169(.a(new_n175), .o1(new_n265));
  aoai13aa1n02x7               g170(.a(new_n177), .b(new_n265), .c(new_n160), .d(new_n162), .o1(new_n266));
  and002aa1n18x5               g171(.a(new_n259), .b(new_n258), .o(new_n267));
  nano23aa1n06x5               g172(.a(new_n209), .b(new_n246), .c(new_n267), .d(new_n228), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n266), .c(new_n141), .d(new_n179), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .c(new_n261), .carry(new_n270));
  aobi12aa1n06x5               g175(.a(new_n270), .b(new_n253), .c(new_n267), .out0(new_n271));
  nor042aa1n04x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  norb02aa1n02x5               g178(.a(new_n273), .b(new_n272), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n269), .c(new_n271), .out0(\s[27] ));
  xorc02aa1n02x5               g180(.a(\a[28] ), .b(\b[27] ), .out0(new_n276));
  aoai13aa1n04x5               g181(.a(new_n245), .b(new_n230), .c(new_n213), .d(new_n228), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n267), .o1(new_n278));
  aoai13aa1n12x5               g183(.a(new_n270), .b(new_n278), .c(new_n277), .d(new_n252), .o1(new_n279));
  aoi112aa1n03x4               g184(.a(new_n279), .b(new_n272), .c(new_n181), .d(new_n268), .o1(new_n280));
  nano22aa1n03x7               g185(.a(new_n280), .b(new_n273), .c(new_n276), .out0(new_n281));
  inv000aa1d42x5               g186(.a(new_n272), .o1(new_n282));
  nanp03aa1n03x5               g187(.a(new_n269), .b(new_n271), .c(new_n282), .o1(new_n283));
  aoi012aa1n03x5               g188(.a(new_n276), .b(new_n283), .c(new_n273), .o1(new_n284));
  nor002aa1n02x5               g189(.a(new_n284), .b(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g190(.a(new_n276), .b(new_n274), .o(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n279), .c(new_n181), .d(new_n268), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .carry(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[28] ), .b(\a[29] ), .out0(new_n289));
  tech160nm_fiaoi012aa1n02p5x5 g194(.a(new_n289), .b(new_n287), .c(new_n288), .o1(new_n290));
  aobi12aa1n02x7               g195(.a(new_n286), .b(new_n269), .c(new_n271), .out0(new_n291));
  nano22aa1n02x4               g196(.a(new_n291), .b(new_n288), .c(new_n289), .out0(new_n292));
  norp02aa1n03x5               g197(.a(new_n290), .b(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g199(.a(new_n289), .b(new_n276), .c(new_n274), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n279), .c(new_n181), .d(new_n268), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[29] ), .b(\b[28] ), .c(new_n288), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[29] ), .b(\a[30] ), .out0(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n298), .b(new_n296), .c(new_n297), .o1(new_n299));
  aobi12aa1n02x7               g204(.a(new_n295), .b(new_n269), .c(new_n271), .out0(new_n300));
  nano22aa1n02x4               g205(.a(new_n300), .b(new_n297), .c(new_n298), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[30] ));
  nano23aa1n02x4               g207(.a(new_n298), .b(new_n289), .c(new_n276), .d(new_n274), .out0(new_n303));
  aobi12aa1n02x7               g208(.a(new_n303), .b(new_n269), .c(new_n271), .out0(new_n304));
  oao003aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .c(new_n297), .carry(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  nano22aa1n02x4               g211(.a(new_n304), .b(new_n305), .c(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n303), .b(new_n279), .c(new_n181), .d(new_n268), .o1(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n306), .b(new_n308), .c(new_n305), .o1(new_n309));
  norp02aa1n03x5               g214(.a(new_n309), .b(new_n307), .o1(\s[31] ));
  xorb03aa1n02x5               g215(.a(new_n102), .b(\b[2] ), .c(new_n103), .out0(\s[3] ));
  oaoi03aa1n02x5               g216(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g218(.a(new_n106), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioai012aa1n05x5   g219(.a(new_n114), .b(new_n106), .c(new_n113), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[5] ), .c(new_n117), .out0(\s[6] ));
  oaoi03aa1n02x5               g221(.a(\a[6] ), .b(\b[5] ), .c(new_n315), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g223(.a(new_n109), .b(new_n317), .c(new_n110), .o1(new_n319));
  xnrb03aa1n03x5               g224(.a(new_n319), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g225(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


