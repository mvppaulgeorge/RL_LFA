// Benchmark "adder" written by ABC on Thu Jul 18 14:53:55 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n327,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n353, new_n355, new_n356, new_n358, new_n359, new_n361,
    new_n362, new_n363, new_n365, new_n366, new_n367;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n20x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  oai112aa1n06x5               g004(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n100));
  orn002aa1n24x5               g005(.a(\a[3] ), .b(\b[2] ), .o(new_n101));
  nand22aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nor042aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanb03aa1n03x5               g009(.a(new_n103), .b(new_n104), .c(new_n102), .out0(new_n105));
  nano32aa1n03x7               g010(.a(new_n105), .b(new_n100), .c(new_n101), .d(new_n99), .out0(new_n106));
  oaoi03aa1n09x5               g011(.a(\a[4] ), .b(\b[3] ), .c(new_n101), .o1(new_n107));
  nor002aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nand02aa1n06x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nor002aa1n16x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n06x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n03x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  nor042aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nand42aa1n03x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  norb02aa1n03x4               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  norp02aa1n02x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand42aa1n04x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  norb02aa1n06x4               g022(.a(new_n117), .b(new_n116), .out0(new_n118));
  nano22aa1n03x7               g023(.a(new_n112), .b(new_n115), .c(new_n118), .out0(new_n119));
  oai012aa1n12x5               g024(.a(new_n119), .b(new_n106), .c(new_n107), .o1(new_n120));
  oai022aa1n02x7               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  nano22aa1n03x7               g026(.a(new_n110), .b(new_n109), .c(new_n111), .out0(new_n122));
  oai022aa1n02x5               g027(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n117), .b(new_n123), .c(new_n122), .d(new_n121), .o1(new_n124));
  nand02aa1d06x5               g029(.a(new_n120), .b(new_n124), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  nand22aa1n03x5               g031(.a(new_n125), .b(new_n126), .o1(new_n127));
  nor042aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanp02aa1n09x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n06x4               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  nona22aa1n02x4               g036(.a(new_n127), .b(new_n128), .c(new_n97), .out0(new_n132));
  nor042aa1d18x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1d04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1n02x5               g039(.a(new_n134), .b(new_n129), .o1(new_n135));
  nona22aa1n03x5               g040(.a(new_n132), .b(new_n133), .c(new_n135), .out0(new_n136));
  inv000aa1d42x5               g041(.a(new_n133), .o1(new_n137));
  aoi022aa1n02x5               g042(.a(new_n132), .b(new_n129), .c(new_n134), .d(new_n137), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n136), .b(new_n138), .out0(\s[11] ));
  aoi022aa1n06x5               g044(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n140));
  aob012aa1n03x5               g045(.a(new_n137), .b(new_n132), .c(new_n140), .out0(new_n141));
  nor042aa1n06x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand22aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  inv000aa1d42x5               g049(.a(\b[11] ), .o1(new_n145));
  nanb02aa1n02x5               g050(.a(\a[12] ), .b(new_n145), .out0(new_n146));
  aoi012aa1n02x5               g051(.a(new_n133), .b(new_n146), .c(new_n143), .o1(new_n147));
  aoi022aa1n02x5               g052(.a(new_n141), .b(new_n144), .c(new_n136), .d(new_n147), .o1(\s[12] ));
  nona23aa1n09x5               g053(.a(new_n143), .b(new_n134), .c(new_n133), .d(new_n142), .out0(new_n149));
  nano22aa1n03x7               g054(.a(new_n149), .b(new_n126), .c(new_n130), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n125), .b(new_n150), .o1(new_n151));
  nanb03aa1n03x5               g056(.a(new_n149), .b(new_n126), .c(new_n130), .out0(new_n152));
  oai112aa1n04x5               g057(.a(new_n146), .b(new_n143), .c(\b[10] ), .d(\a[11] ), .o1(new_n153));
  tech160nm_fioai012aa1n04x5   g058(.a(new_n140), .b(new_n128), .c(new_n97), .o1(new_n154));
  aoi012aa1n09x5               g059(.a(new_n142), .b(new_n133), .c(new_n143), .o1(new_n155));
  oai012aa1n02x5               g060(.a(new_n155), .b(new_n153), .c(new_n154), .o1(new_n156));
  inv020aa1n02x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n152), .c(new_n120), .d(new_n124), .o1(new_n158));
  nor042aa1d18x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand02aa1d04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  norb03aa1n03x5               g067(.a(new_n143), .b(new_n133), .c(new_n142), .out0(new_n163));
  oab012aa1n06x5               g068(.a(new_n135), .b(new_n97), .c(new_n128), .out0(new_n164));
  inv000aa1n02x5               g069(.a(new_n155), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n162), .c(new_n164), .d(new_n163), .o1(new_n166));
  aoi022aa1n02x5               g071(.a(new_n158), .b(new_n162), .c(new_n151), .d(new_n166), .o1(\s[13] ));
  inv000aa1d42x5               g072(.a(new_n159), .o1(new_n168));
  nanp02aa1n02x5               g073(.a(new_n158), .b(new_n162), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand02aa1d04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(new_n172));
  xobna2aa1n03x5               g077(.a(new_n172), .b(new_n169), .c(new_n168), .out0(\s[14] ));
  nona23aa1d18x5               g078(.a(new_n171), .b(new_n160), .c(new_n159), .d(new_n170), .out0(new_n174));
  inv040aa1n06x5               g079(.a(new_n174), .o1(new_n175));
  oaoi03aa1n12x5               g080(.a(\a[14] ), .b(\b[13] ), .c(new_n168), .o1(new_n176));
  xorc02aa1n12x5               g081(.a(\a[15] ), .b(\b[14] ), .out0(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n176), .c(new_n158), .d(new_n175), .o1(new_n178));
  aoi112aa1n02x5               g083(.a(new_n177), .b(new_n176), .c(new_n158), .d(new_n175), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(\s[15] ));
  inv000aa1d42x5               g085(.a(\a[15] ), .o1(new_n181));
  oaib12aa1n02x5               g086(.a(new_n178), .b(\b[14] ), .c(new_n181), .out0(new_n182));
  tech160nm_fixorc02aa1n02p5x5 g087(.a(\a[16] ), .b(\b[15] ), .out0(new_n183));
  nor042aa1n03x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norp02aa1n02x5               g089(.a(new_n183), .b(new_n184), .o1(new_n185));
  aoi022aa1n02x5               g090(.a(new_n182), .b(new_n183), .c(new_n178), .d(new_n185), .o1(\s[16] ));
  inv000aa1d42x5               g091(.a(\a[16] ), .o1(new_n187));
  xroi22aa1d04x5               g092(.a(new_n181), .b(\b[14] ), .c(new_n187), .d(\b[15] ), .out0(new_n188));
  nano22aa1n03x7               g093(.a(new_n152), .b(new_n175), .c(new_n188), .out0(new_n189));
  nand22aa1n12x5               g094(.a(new_n125), .b(new_n189), .o1(new_n190));
  oaoi13aa1n09x5               g095(.a(new_n174), .b(new_n155), .c(new_n153), .d(new_n154), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[15] ), .o1(new_n192));
  oaoi03aa1n12x5               g097(.a(new_n187), .b(new_n192), .c(new_n184), .o1(new_n193));
  inv000aa1n02x5               g098(.a(new_n193), .o1(new_n194));
  oaoi13aa1n12x5               g099(.a(new_n194), .b(new_n188), .c(new_n191), .d(new_n176), .o1(new_n195));
  nand22aa1n12x5               g100(.a(new_n190), .b(new_n195), .o1(new_n196));
  xorc02aa1n12x5               g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  nanb02aa1n02x5               g102(.a(new_n197), .b(new_n193), .out0(new_n198));
  oaoi13aa1n02x5               g103(.a(new_n198), .b(new_n188), .c(new_n191), .d(new_n176), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n196), .b(new_n197), .c(new_n190), .d(new_n199), .o1(\s[17] ));
  nor002aa1d32x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  nand02aa1d04x5               g107(.a(new_n183), .b(new_n177), .o1(new_n203));
  nona22aa1n03x5               g108(.a(new_n150), .b(new_n203), .c(new_n174), .out0(new_n204));
  aoi012aa1d18x5               g109(.a(new_n204), .b(new_n120), .c(new_n124), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n176), .o1(new_n206));
  aoai13aa1n12x5               g111(.a(new_n175), .b(new_n165), .c(new_n164), .d(new_n163), .o1(new_n207));
  aoai13aa1n12x5               g112(.a(new_n193), .b(new_n203), .c(new_n207), .d(new_n206), .o1(new_n208));
  oai012aa1n06x5               g113(.a(new_n197), .b(new_n208), .c(new_n205), .o1(new_n209));
  nor002aa1n10x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nand22aa1n09x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  norb02aa1n06x5               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n209), .c(new_n202), .out0(\s[18] ));
  and002aa1n02x5               g118(.a(new_n197), .b(new_n212), .o(new_n214));
  tech160nm_fioai012aa1n05x5   g119(.a(new_n214), .b(new_n208), .c(new_n205), .o1(new_n215));
  oaoi03aa1n02x5               g120(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  nor042aa1d18x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nand02aa1n08x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  norb02aa1n09x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  xnbna2aa1n03x5               g125(.a(new_n220), .b(new_n215), .c(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g127(.a(new_n220), .b(new_n216), .c(new_n196), .d(new_n214), .o1(new_n223));
  inv030aa1n03x5               g128(.a(new_n218), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n220), .o1(new_n225));
  aoai13aa1n02x7               g130(.a(new_n224), .b(new_n225), .c(new_n215), .d(new_n217), .o1(new_n226));
  nor002aa1d32x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nand02aa1d28x5               g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  norb02aa1n06x4               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  inv000aa1d42x5               g134(.a(\a[19] ), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\b[18] ), .o1(new_n231));
  aboi22aa1n03x5               g136(.a(new_n227), .b(new_n228), .c(new_n230), .d(new_n231), .out0(new_n232));
  aoi022aa1n03x5               g137(.a(new_n226), .b(new_n229), .c(new_n223), .d(new_n232), .o1(\s[20] ));
  nano32aa1n09x5               g138(.a(new_n225), .b(new_n197), .c(new_n229), .d(new_n212), .out0(new_n234));
  tech160nm_fioai012aa1n05x5   g139(.a(new_n234), .b(new_n208), .c(new_n205), .o1(new_n235));
  inv000aa1n02x5               g140(.a(new_n234), .o1(new_n236));
  nanb03aa1n09x5               g141(.a(new_n227), .b(new_n228), .c(new_n219), .out0(new_n237));
  oai112aa1n06x5               g142(.a(new_n224), .b(new_n211), .c(new_n210), .d(new_n201), .o1(new_n238));
  aoi012aa1d18x5               g143(.a(new_n227), .b(new_n218), .c(new_n228), .o1(new_n239));
  oai012aa1n18x5               g144(.a(new_n239), .b(new_n238), .c(new_n237), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n04x5               g146(.a(new_n241), .b(new_n236), .c(new_n190), .d(new_n195), .o1(new_n242));
  nor002aa1d32x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  nand42aa1d28x5               g148(.a(\b[20] ), .b(\a[21] ), .o1(new_n244));
  norb02aa1n03x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  nano22aa1n12x5               g150(.a(new_n227), .b(new_n219), .c(new_n228), .out0(new_n246));
  oai012aa1n02x5               g151(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .o1(new_n247));
  oab012aa1n03x5               g152(.a(new_n247), .b(new_n201), .c(new_n210), .out0(new_n248));
  inv000aa1n02x5               g153(.a(new_n239), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(new_n249), .b(new_n245), .c(new_n248), .d(new_n246), .o1(new_n250));
  aoi022aa1n02x5               g155(.a(new_n242), .b(new_n245), .c(new_n235), .d(new_n250), .o1(\s[21] ));
  nand22aa1n02x5               g156(.a(new_n242), .b(new_n245), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n243), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n245), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n253), .b(new_n254), .c(new_n235), .d(new_n241), .o1(new_n255));
  nor042aa1n09x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  nand42aa1d28x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  aoib12aa1n02x5               g163(.a(new_n243), .b(new_n257), .c(new_n256), .out0(new_n259));
  aoi022aa1n03x5               g164(.a(new_n255), .b(new_n258), .c(new_n252), .d(new_n259), .o1(\s[22] ));
  nano23aa1d15x5               g165(.a(new_n243), .b(new_n256), .c(new_n257), .d(new_n244), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  nano32aa1n02x4               g167(.a(new_n262), .b(new_n214), .c(new_n220), .d(new_n229), .out0(new_n263));
  oai012aa1n06x5               g168(.a(new_n263), .b(new_n208), .c(new_n205), .o1(new_n264));
  aoi012aa1d24x5               g169(.a(new_n256), .b(new_n243), .c(new_n257), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  tech160nm_fiaoi012aa1n03p5x5 g171(.a(new_n266), .b(new_n240), .c(new_n261), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  xorc02aa1n12x5               g173(.a(\a[23] ), .b(\b[22] ), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n268), .c(new_n196), .d(new_n263), .o1(new_n270));
  aoi112aa1n02x5               g175(.a(new_n269), .b(new_n266), .c(new_n240), .d(new_n261), .o1(new_n271));
  aobi12aa1n02x7               g176(.a(new_n270), .b(new_n271), .c(new_n264), .out0(\s[23] ));
  nor042aa1n09x5               g177(.a(\b[22] ), .b(\a[23] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n269), .o1(new_n275));
  aoai13aa1n03x5               g180(.a(new_n274), .b(new_n275), .c(new_n264), .d(new_n267), .o1(new_n276));
  tech160nm_fixorc02aa1n02p5x5 g181(.a(\a[24] ), .b(\b[23] ), .out0(new_n277));
  norp02aa1n02x5               g182(.a(new_n277), .b(new_n273), .o1(new_n278));
  aoi022aa1n02x7               g183(.a(new_n276), .b(new_n277), .c(new_n270), .d(new_n278), .o1(\s[24] ));
  and002aa1n12x5               g184(.a(new_n277), .b(new_n269), .o(new_n280));
  nano22aa1n02x5               g185(.a(new_n236), .b(new_n261), .c(new_n280), .out0(new_n281));
  tech160nm_fioai012aa1n05x5   g186(.a(new_n281), .b(new_n208), .c(new_n205), .o1(new_n282));
  aoai13aa1n06x5               g187(.a(new_n261), .b(new_n249), .c(new_n248), .d(new_n246), .o1(new_n283));
  inv030aa1n04x5               g188(.a(new_n280), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[24] ), .b(\b[23] ), .c(new_n274), .carry(new_n285));
  aoai13aa1n12x5               g190(.a(new_n285), .b(new_n284), .c(new_n283), .d(new_n265), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[25] ), .b(\b[24] ), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n287), .b(new_n286), .c(new_n196), .d(new_n281), .o1(new_n288));
  aoai13aa1n04x5               g193(.a(new_n280), .b(new_n266), .c(new_n240), .d(new_n261), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n287), .o1(new_n290));
  and003aa1n02x5               g195(.a(new_n289), .b(new_n290), .c(new_n285), .o(new_n291));
  aobi12aa1n03x7               g196(.a(new_n288), .b(new_n291), .c(new_n282), .out0(\s[25] ));
  inv000aa1d42x5               g197(.a(new_n286), .o1(new_n293));
  nor042aa1n06x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n290), .c(new_n282), .d(new_n293), .o1(new_n296));
  tech160nm_fixorc02aa1n03p5x5 g201(.a(\a[26] ), .b(\b[25] ), .out0(new_n297));
  norp02aa1n02x5               g202(.a(new_n297), .b(new_n294), .o1(new_n298));
  aoi022aa1n02x7               g203(.a(new_n296), .b(new_n297), .c(new_n288), .d(new_n298), .o1(\s[26] ));
  and002aa1n12x5               g204(.a(new_n297), .b(new_n287), .o(new_n300));
  nano32aa1n03x7               g205(.a(new_n236), .b(new_n300), .c(new_n261), .d(new_n280), .out0(new_n301));
  oai012aa1n18x5               g206(.a(new_n301), .b(new_n208), .c(new_n205), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n300), .o1(new_n303));
  oao003aa1n06x5               g208(.a(\a[26] ), .b(\b[25] ), .c(new_n295), .carry(new_n304));
  aoai13aa1n04x5               g209(.a(new_n304), .b(new_n303), .c(new_n289), .d(new_n285), .o1(new_n305));
  xorc02aa1n12x5               g210(.a(\a[27] ), .b(\b[26] ), .out0(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n305), .c(new_n196), .d(new_n301), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n304), .o1(new_n308));
  aoi112aa1n02x5               g213(.a(new_n306), .b(new_n308), .c(new_n286), .d(new_n300), .o1(new_n309));
  aobi12aa1n02x7               g214(.a(new_n307), .b(new_n309), .c(new_n302), .out0(\s[27] ));
  aoi012aa1d18x5               g215(.a(new_n308), .b(new_n286), .c(new_n300), .o1(new_n311));
  norp02aa1n02x5               g216(.a(\b[26] ), .b(\a[27] ), .o1(new_n312));
  inv000aa1n03x5               g217(.a(new_n312), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n306), .o1(new_n314));
  aoai13aa1n06x5               g219(.a(new_n313), .b(new_n314), .c(new_n302), .d(new_n311), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .out0(new_n316));
  norp02aa1n02x5               g221(.a(new_n316), .b(new_n312), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n315), .b(new_n316), .c(new_n307), .d(new_n317), .o1(\s[28] ));
  and002aa1n02x5               g223(.a(new_n316), .b(new_n306), .o(new_n319));
  aoai13aa1n02x5               g224(.a(new_n319), .b(new_n305), .c(new_n196), .d(new_n301), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n319), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[28] ), .b(\b[27] ), .c(new_n313), .carry(new_n322));
  aoai13aa1n06x5               g227(.a(new_n322), .b(new_n321), .c(new_n302), .d(new_n311), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[29] ), .b(\b[28] ), .out0(new_n324));
  norb02aa1n02x5               g229(.a(new_n322), .b(new_n324), .out0(new_n325));
  aoi022aa1n03x5               g230(.a(new_n323), .b(new_n324), .c(new_n320), .d(new_n325), .o1(\s[29] ));
  nanp02aa1n02x5               g231(.a(\b[0] ), .b(\a[1] ), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g233(.a(new_n314), .b(new_n316), .c(new_n324), .out0(new_n329));
  aoai13aa1n02x5               g234(.a(new_n329), .b(new_n305), .c(new_n196), .d(new_n301), .o1(new_n330));
  inv000aa1n02x5               g235(.a(new_n329), .o1(new_n331));
  inv000aa1d42x5               g236(.a(\b[28] ), .o1(new_n332));
  inv000aa1d42x5               g237(.a(\a[29] ), .o1(new_n333));
  oaib12aa1n02x5               g238(.a(new_n322), .b(\b[28] ), .c(new_n333), .out0(new_n334));
  oaib12aa1n02x5               g239(.a(new_n334), .b(new_n332), .c(\a[29] ), .out0(new_n335));
  aoai13aa1n06x5               g240(.a(new_n335), .b(new_n331), .c(new_n302), .d(new_n311), .o1(new_n336));
  xorc02aa1n02x5               g241(.a(\a[30] ), .b(\b[29] ), .out0(new_n337));
  oaoi13aa1n02x5               g242(.a(new_n337), .b(new_n334), .c(new_n333), .d(new_n332), .o1(new_n338));
  aoi022aa1n03x5               g243(.a(new_n336), .b(new_n337), .c(new_n330), .d(new_n338), .o1(\s[30] ));
  nanb02aa1n02x5               g244(.a(\a[31] ), .b(\b[30] ), .out0(new_n340));
  nanb02aa1n02x5               g245(.a(\b[30] ), .b(\a[31] ), .out0(new_n341));
  nanp02aa1n02x5               g246(.a(new_n341), .b(new_n340), .o1(new_n342));
  nano32aa1n03x7               g247(.a(new_n314), .b(new_n337), .c(new_n316), .d(new_n324), .out0(new_n343));
  aoai13aa1n02x5               g248(.a(new_n343), .b(new_n305), .c(new_n196), .d(new_n301), .o1(new_n344));
  inv000aa1d42x5               g249(.a(new_n343), .o1(new_n345));
  norp02aa1n02x5               g250(.a(\b[29] ), .b(\a[30] ), .o1(new_n346));
  aoi022aa1n02x5               g251(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n347));
  aoi012aa1n02x5               g252(.a(new_n346), .b(new_n334), .c(new_n347), .o1(new_n348));
  aoai13aa1n06x5               g253(.a(new_n348), .b(new_n345), .c(new_n302), .d(new_n311), .o1(new_n349));
  oai112aa1n02x5               g254(.a(new_n340), .b(new_n341), .c(\b[29] ), .d(\a[30] ), .o1(new_n350));
  aoi012aa1n02x5               g255(.a(new_n350), .b(new_n334), .c(new_n347), .o1(new_n351));
  aoi022aa1n03x5               g256(.a(new_n349), .b(new_n342), .c(new_n344), .d(new_n351), .o1(\s[31] ));
  xorc02aa1n02x5               g257(.a(\a[3] ), .b(\b[2] ), .out0(new_n353));
  xobna2aa1n03x5               g258(.a(new_n353), .b(new_n100), .c(new_n99), .out0(\s[3] ));
  nanb02aa1n02x5               g259(.a(new_n103), .b(new_n104), .out0(new_n355));
  aob012aa1n02x5               g260(.a(new_n353), .b(new_n100), .c(new_n99), .out0(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n355), .b(new_n356), .c(new_n102), .out0(\s[4] ));
  oai012aa1n03x5               g262(.a(new_n115), .b(new_n106), .c(new_n107), .o1(new_n358));
  norp03aa1n02x5               g263(.a(new_n106), .b(new_n107), .c(new_n115), .o1(new_n359));
  norb02aa1n02x5               g264(.a(new_n358), .b(new_n359), .out0(\s[5] ));
  nanb02aa1n02x5               g265(.a(new_n108), .b(new_n109), .out0(new_n361));
  oaoi13aa1n02x5               g266(.a(new_n113), .b(new_n114), .c(new_n106), .d(new_n107), .o1(new_n362));
  nona23aa1n02x4               g267(.a(new_n358), .b(new_n109), .c(new_n108), .d(new_n113), .out0(new_n363));
  oaib12aa1n02x5               g268(.a(new_n363), .b(new_n362), .c(new_n361), .out0(\s[6] ));
  inv000aa1d42x5               g269(.a(new_n110), .o1(new_n365));
  aoi022aa1n02x5               g270(.a(new_n363), .b(new_n109), .c(new_n365), .d(new_n111), .o1(new_n366));
  nanp02aa1n03x5               g271(.a(new_n363), .b(new_n122), .o1(new_n367));
  norb02aa1n02x5               g272(.a(new_n367), .b(new_n366), .out0(\s[7] ));
  xnbna2aa1n03x5               g273(.a(new_n118), .b(new_n367), .c(new_n365), .out0(\s[8] ));
  xnbna2aa1n03x5               g274(.a(new_n126), .b(new_n120), .c(new_n124), .out0(\s[9] ));
endmodule


