// Benchmark "adder" written by ABC on Thu Jul 18 05:04:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n130, new_n131, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n177, new_n178, new_n179, new_n180, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n193, new_n194, new_n195, new_n196, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n209, new_n210, new_n211, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n304, new_n305, new_n306, new_n309, new_n311, new_n313;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv020aa1d32x5               g001(.a(\b[2] ), .o1(new_n97));
  nanb02aa1d24x5               g002(.a(\a[3] ), .b(new_n97), .out0(new_n98));
  nand02aa1d16x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nand42aa1n16x5               g004(.a(new_n98), .b(new_n99), .o1(new_n100));
  nanp02aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor042aa1n09x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand02aa1d24x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  oai012aa1d24x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  oa0022aa1n06x5               g009(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n105));
  oai012aa1d24x5               g010(.a(new_n105), .b(new_n104), .c(new_n100), .o1(new_n106));
  nand42aa1n08x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  inv040aa1d32x5               g012(.a(\a[6] ), .o1(new_n108));
  inv040aa1n16x5               g013(.a(\b[5] ), .o1(new_n109));
  nanp02aa1n12x5               g014(.a(new_n109), .b(new_n108), .o1(new_n110));
  nand42aa1n08x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand02aa1n06x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nanb02aa1n12x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  nano32aa1n09x5               g019(.a(new_n114), .b(new_n110), .c(new_n111), .d(new_n107), .out0(new_n115));
  nand42aa1d28x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nor002aa1n12x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor002aa1d32x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand42aa1d28x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n118), .b(new_n117), .c(new_n119), .d(new_n116), .out0(new_n120));
  nona23aa1n09x5               g025(.a(new_n116), .b(new_n119), .c(new_n118), .d(new_n117), .out0(new_n121));
  tech160nm_fioaoi03aa1n02p5x5 g026(.a(new_n108), .b(new_n109), .c(new_n112), .o1(new_n122));
  oaih12aa1n02x5               g027(.a(new_n116), .b(new_n118), .c(new_n117), .o1(new_n123));
  oai012aa1n06x5               g028(.a(new_n123), .b(new_n121), .c(new_n122), .o1(new_n124));
  aoi013aa1n09x5               g029(.a(new_n124), .b(new_n106), .c(new_n115), .d(new_n120), .o1(new_n125));
  oao003aa1n03x5               g030(.a(\a[9] ), .b(\b[8] ), .c(new_n125), .carry(new_n126));
  xnrb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  oaoi03aa1n09x5               g032(.a(\a[10] ), .b(\b[9] ), .c(new_n126), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nand42aa1n16x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor002aa1n20x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  xnrc02aa1n12x5               g036(.a(\b[11] ), .b(\a[12] ), .out0(new_n132));
  aoai13aa1n03x5               g037(.a(new_n132), .b(new_n131), .c(new_n128), .d(new_n130), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n130), .b(new_n131), .out0(new_n134));
  nand42aa1n02x5               g039(.a(new_n128), .b(new_n134), .o1(new_n135));
  nona22aa1n03x5               g040(.a(new_n135), .b(new_n132), .c(new_n131), .out0(new_n136));
  nanp02aa1n03x5               g041(.a(new_n136), .b(new_n133), .o1(\s[12] ));
  nor022aa1n16x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  nand02aa1n08x5               g043(.a(\b[9] ), .b(\a[10] ), .o1(new_n139));
  nona23aa1n09x5               g044(.a(new_n130), .b(new_n139), .c(new_n131), .d(new_n138), .out0(new_n140));
  xnrc02aa1n03x5               g045(.a(\b[8] ), .b(\a[9] ), .out0(new_n141));
  orn003aa1n02x5               g046(.a(new_n140), .b(new_n132), .c(new_n141), .o(new_n142));
  oai022aa1d18x5               g047(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n143));
  nand03aa1n06x5               g048(.a(new_n143), .b(new_n139), .c(new_n130), .o1(new_n144));
  oai122aa1n12x5               g049(.a(new_n144), .b(\a[12] ), .c(\b[11] ), .d(\a[11] ), .e(\b[10] ), .o1(new_n145));
  aob012aa1n02x5               g050(.a(new_n145), .b(\b[11] ), .c(\a[12] ), .out0(new_n146));
  tech160nm_fioai012aa1n05x5   g051(.a(new_n146), .b(new_n125), .c(new_n142), .o1(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n12x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nand42aa1n08x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  aoi012aa1n02x5               g055(.a(new_n149), .b(new_n147), .c(new_n150), .o1(new_n151));
  xnrb03aa1n02x5               g056(.a(new_n151), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nand02aa1n16x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nor022aa1n16x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nano23aa1n03x7               g059(.a(new_n149), .b(new_n154), .c(new_n153), .d(new_n150), .out0(new_n155));
  nanp02aa1n03x5               g060(.a(new_n147), .b(new_n155), .o1(new_n156));
  oai022aa1d18x5               g061(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n157));
  aob012aa1n06x5               g062(.a(new_n156), .b(new_n157), .c(new_n153), .out0(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nand02aa1n08x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[15] ), .b(\a[16] ), .out0(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n160), .c(new_n158), .d(new_n161), .o1(new_n163));
  nanb02aa1n12x5               g068(.a(new_n160), .b(new_n161), .out0(new_n164));
  nanb02aa1n03x5               g069(.a(new_n164), .b(new_n158), .out0(new_n165));
  nona22aa1n02x4               g070(.a(new_n165), .b(new_n162), .c(new_n160), .out0(new_n166));
  nanp02aa1n03x5               g071(.a(new_n166), .b(new_n163), .o1(\s[16] ));
  nona23aa1d18x5               g072(.a(new_n153), .b(new_n150), .c(new_n149), .d(new_n154), .out0(new_n168));
  nor043aa1d12x5               g073(.a(new_n168), .b(new_n164), .c(new_n162), .o1(new_n169));
  nona32aa1n09x5               g074(.a(new_n169), .b(new_n140), .c(new_n141), .d(new_n132), .out0(new_n170));
  aoi022aa1n06x5               g075(.a(\b[15] ), .b(\a[16] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n171));
  aoai13aa1n04x5               g076(.a(new_n161), .b(new_n160), .c(new_n157), .d(new_n153), .o1(new_n172));
  oaoi03aa1n12x5               g077(.a(\a[16] ), .b(\b[15] ), .c(new_n172), .o1(new_n173));
  aoi013aa1n06x4               g078(.a(new_n173), .b(new_n169), .c(new_n145), .d(new_n171), .o1(new_n174));
  oai012aa1d24x5               g079(.a(new_n174), .b(new_n125), .c(new_n170), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g081(.a(\a[18] ), .o1(new_n177));
  inv040aa1d30x5               g082(.a(\a[17] ), .o1(new_n178));
  inv000aa1d42x5               g083(.a(\b[16] ), .o1(new_n179));
  oaoi03aa1n03x5               g084(.a(new_n178), .b(new_n179), .c(new_n175), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[17] ), .c(new_n177), .out0(\s[18] ));
  xroi22aa1d06x4               g086(.a(new_n178), .b(\b[16] ), .c(new_n177), .d(\b[17] ), .out0(new_n182));
  nand22aa1n06x5               g087(.a(\b[17] ), .b(\a[18] ), .o1(new_n183));
  nona22aa1n03x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(new_n184));
  oaib12aa1n09x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n177), .out0(new_n185));
  nor002aa1d32x5               g090(.a(\b[18] ), .b(\a[19] ), .o1(new_n186));
  nand22aa1n12x5               g091(.a(\b[18] ), .b(\a[19] ), .o1(new_n187));
  norb02aa1n02x5               g092(.a(new_n187), .b(new_n186), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n185), .c(new_n175), .d(new_n182), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(new_n188), .b(new_n185), .c(new_n175), .d(new_n182), .o1(new_n190));
  norb02aa1n02x7               g095(.a(new_n189), .b(new_n190), .out0(\s[19] ));
  xnrc02aa1n02x5               g096(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g097(.a(new_n186), .o1(new_n193));
  nor002aa1d32x5               g098(.a(\b[19] ), .b(\a[20] ), .o1(new_n194));
  nand02aa1n08x5               g099(.a(\b[19] ), .b(\a[20] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n189), .c(new_n193), .out0(\s[20] ));
  nona23aa1n09x5               g102(.a(new_n195), .b(new_n187), .c(new_n186), .d(new_n194), .out0(new_n198));
  norb02aa1n03x5               g103(.a(new_n182), .b(new_n198), .out0(new_n199));
  norp02aa1n02x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  aoi013aa1n02x4               g105(.a(new_n200), .b(new_n183), .c(new_n178), .d(new_n179), .o1(new_n201));
  oaoi03aa1n09x5               g106(.a(\a[20] ), .b(\b[19] ), .c(new_n193), .o1(new_n202));
  inv040aa1n03x5               g107(.a(new_n202), .o1(new_n203));
  oai012aa1n06x5               g108(.a(new_n203), .b(new_n198), .c(new_n201), .o1(new_n204));
  xorc02aa1n02x5               g109(.a(\a[21] ), .b(\b[20] ), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n204), .c(new_n175), .d(new_n199), .o1(new_n206));
  aoi112aa1n02x5               g111(.a(new_n205), .b(new_n204), .c(new_n175), .d(new_n199), .o1(new_n207));
  norb02aa1n02x7               g112(.a(new_n206), .b(new_n207), .out0(\s[21] ));
  nor042aa1n03x5               g113(.a(\b[20] ), .b(\a[21] ), .o1(new_n209));
  inv000aa1n03x5               g114(.a(new_n209), .o1(new_n210));
  xorc02aa1n02x5               g115(.a(\a[22] ), .b(\b[21] ), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n206), .c(new_n210), .out0(\s[22] ));
  nano23aa1d15x5               g117(.a(new_n186), .b(new_n194), .c(new_n195), .d(new_n187), .out0(new_n213));
  inv000aa1d42x5               g118(.a(\a[21] ), .o1(new_n214));
  inv040aa1n09x5               g119(.a(\a[22] ), .o1(new_n215));
  xroi22aa1d06x4               g120(.a(new_n214), .b(\b[20] ), .c(new_n215), .d(\b[21] ), .out0(new_n216));
  nand03aa1n02x5               g121(.a(new_n216), .b(new_n182), .c(new_n213), .o1(new_n217));
  inv000aa1n02x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n216), .b(new_n202), .c(new_n213), .d(new_n185), .o1(new_n219));
  oaoi03aa1n02x5               g124(.a(\a[22] ), .b(\b[21] ), .c(new_n210), .o1(new_n220));
  inv000aa1n02x5               g125(.a(new_n220), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(new_n219), .b(new_n221), .o1(new_n222));
  xorc02aa1n12x5               g127(.a(\a[23] ), .b(\b[22] ), .out0(new_n223));
  aoai13aa1n06x5               g128(.a(new_n223), .b(new_n222), .c(new_n175), .d(new_n218), .o1(new_n224));
  aoi112aa1n02x5               g129(.a(new_n223), .b(new_n222), .c(new_n175), .d(new_n218), .o1(new_n225));
  norb02aa1n02x7               g130(.a(new_n224), .b(new_n225), .out0(\s[23] ));
  nor042aa1n06x5               g131(.a(\b[22] ), .b(\a[23] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  xnrc02aa1n12x5               g133(.a(\b[23] ), .b(\a[24] ), .out0(new_n229));
  xobna2aa1n03x5               g134(.a(new_n229), .b(new_n224), .c(new_n228), .out0(\s[24] ));
  nanp03aa1n02x5               g135(.a(new_n106), .b(new_n115), .c(new_n120), .o1(new_n231));
  nanb02aa1n02x5               g136(.a(new_n124), .b(new_n231), .out0(new_n232));
  inv040aa1n03x5               g137(.a(new_n170), .o1(new_n233));
  nona23aa1n03x5               g138(.a(new_n155), .b(new_n171), .c(new_n162), .d(new_n164), .out0(new_n234));
  inv000aa1n02x5               g139(.a(new_n173), .o1(new_n235));
  oaib12aa1n06x5               g140(.a(new_n235), .b(new_n234), .c(new_n145), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n199), .b(new_n236), .c(new_n232), .d(new_n233), .o1(new_n237));
  norb02aa1n03x4               g142(.a(new_n223), .b(new_n229), .out0(new_n238));
  inv030aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  oao003aa1n02x5               g144(.a(\a[24] ), .b(\b[23] ), .c(new_n228), .carry(new_n240));
  aoai13aa1n04x5               g145(.a(new_n240), .b(new_n239), .c(new_n219), .d(new_n221), .o1(new_n241));
  nanp02aa1n02x5               g146(.a(new_n238), .b(new_n216), .o1(new_n242));
  oabi12aa1n06x5               g147(.a(new_n241), .b(new_n237), .c(new_n242), .out0(new_n243));
  xorb03aa1n02x5               g148(.a(new_n243), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g149(.a(\b[24] ), .b(\a[25] ), .o1(new_n245));
  xorc02aa1n12x5               g150(.a(\a[25] ), .b(\b[24] ), .out0(new_n246));
  nor002aa1n02x5               g151(.a(\b[25] ), .b(\a[26] ), .o1(new_n247));
  nand42aa1n03x5               g152(.a(\b[25] ), .b(\a[26] ), .o1(new_n248));
  nanb02aa1n06x5               g153(.a(new_n247), .b(new_n248), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n245), .c(new_n243), .d(new_n246), .o1(new_n250));
  aoi012aa1n06x5               g155(.a(new_n236), .b(new_n232), .c(new_n233), .o1(new_n251));
  nano32aa1n03x7               g156(.a(new_n251), .b(new_n238), .c(new_n199), .d(new_n216), .out0(new_n252));
  oai012aa1n02x5               g157(.a(new_n246), .b(new_n252), .c(new_n241), .o1(new_n253));
  nona22aa1n02x5               g158(.a(new_n253), .b(new_n249), .c(new_n245), .out0(new_n254));
  nanp02aa1n03x5               g159(.a(new_n250), .b(new_n254), .o1(\s[26] ));
  norb02aa1n06x4               g160(.a(new_n246), .b(new_n249), .out0(new_n256));
  oai012aa1n02x5               g161(.a(new_n248), .b(new_n247), .c(new_n245), .o1(new_n257));
  aobi12aa1n09x5               g162(.a(new_n257), .b(new_n241), .c(new_n256), .out0(new_n258));
  inv000aa1n02x5               g163(.a(new_n256), .o1(new_n259));
  nona32aa1n09x5               g164(.a(new_n175), .b(new_n259), .c(new_n239), .d(new_n217), .out0(new_n260));
  xorc02aa1n02x5               g165(.a(\a[27] ), .b(\b[26] ), .out0(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n258), .c(new_n260), .out0(\s[27] ));
  nand42aa1n06x5               g167(.a(new_n258), .b(new_n260), .o1(new_n263));
  norp02aa1n02x5               g168(.a(\b[26] ), .b(\a[27] ), .o1(new_n264));
  norp02aa1n02x5               g169(.a(\b[27] ), .b(\a[28] ), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(\b[27] ), .b(\a[28] ), .o1(new_n266));
  norb02aa1n09x5               g171(.a(new_n266), .b(new_n265), .out0(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n264), .c(new_n263), .d(new_n261), .o1(new_n269));
  oaoi13aa1n04x5               g174(.a(new_n217), .b(new_n174), .c(new_n125), .d(new_n170), .o1(new_n270));
  aoai13aa1n02x7               g175(.a(new_n238), .b(new_n220), .c(new_n204), .d(new_n216), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n257), .b(new_n259), .c(new_n271), .d(new_n240), .o1(new_n272));
  nano23aa1n02x4               g177(.a(new_n249), .b(new_n229), .c(new_n223), .d(new_n246), .out0(new_n273));
  aoai13aa1n03x5               g178(.a(new_n261), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n274));
  nona22aa1n02x5               g179(.a(new_n274), .b(new_n268), .c(new_n264), .out0(new_n275));
  nanp02aa1n03x5               g180(.a(new_n269), .b(new_n275), .o1(\s[28] ));
  tech160nm_fixorc02aa1n03p5x5 g181(.a(\a[29] ), .b(\b[28] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n261), .b(new_n268), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n280));
  aoi012aa1n02x5               g185(.a(new_n265), .b(new_n264), .c(new_n266), .o1(new_n281));
  tech160nm_fiaoi012aa1n02p5x5 g186(.a(new_n278), .b(new_n280), .c(new_n281), .o1(new_n282));
  aobi12aa1n06x5               g187(.a(new_n279), .b(new_n258), .c(new_n260), .out0(new_n283));
  nano22aa1n03x5               g188(.a(new_n283), .b(new_n278), .c(new_n281), .out0(new_n284));
  norp02aa1n03x5               g189(.a(new_n282), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g190(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g191(.a(new_n278), .b(new_n261), .c(new_n267), .out0(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n288));
  xorc02aa1n02x5               g193(.a(\a[30] ), .b(\b[29] ), .out0(new_n289));
  norp02aa1n02x5               g194(.a(\b[28] ), .b(\a[29] ), .o1(new_n290));
  aoi012aa1n02x5               g195(.a(new_n281), .b(\a[29] ), .c(\b[28] ), .o1(new_n291));
  norp03aa1n02x5               g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .c(new_n281), .carry(new_n293));
  nand42aa1n02x5               g198(.a(new_n288), .b(new_n293), .o1(new_n294));
  aoi022aa1n02x7               g199(.a(new_n294), .b(new_n289), .c(new_n288), .d(new_n292), .o1(\s[30] ));
  nand23aa1n03x5               g200(.a(new_n279), .b(new_n277), .c(new_n289), .o1(new_n296));
  nanb02aa1n03x5               g201(.a(new_n296), .b(new_n263), .out0(new_n297));
  xorc02aa1n02x5               g202(.a(\a[31] ), .b(\b[30] ), .out0(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n299));
  norb02aa1n02x5               g204(.a(new_n299), .b(new_n298), .out0(new_n300));
  aoai13aa1n02x7               g205(.a(new_n299), .b(new_n296), .c(new_n258), .d(new_n260), .o1(new_n301));
  aoi022aa1n03x5               g206(.a(new_n297), .b(new_n300), .c(new_n301), .d(new_n298), .o1(\s[31] ));
  xnbna2aa1n03x5               g207(.a(new_n104), .b(new_n98), .c(new_n99), .out0(\s[3] ));
  orn002aa1n02x5               g208(.a(\a[4] ), .b(\b[3] ), .o(new_n304));
  aob012aa1n02x5               g209(.a(new_n98), .b(new_n304), .c(new_n111), .out0(new_n305));
  oab012aa1n02x4               g210(.a(new_n305), .b(new_n100), .c(new_n104), .out0(new_n306));
  aoi013aa1n02x4               g211(.a(new_n306), .b(new_n106), .c(new_n111), .d(new_n304), .o1(\s[4] ));
  xnbna2aa1n03x5               g212(.a(new_n114), .b(new_n106), .c(new_n111), .out0(\s[5] ));
  aoi013aa1n02x4               g213(.a(new_n112), .b(new_n106), .c(new_n111), .d(new_n113), .o1(new_n309));
  xnbna2aa1n03x5               g214(.a(new_n309), .b(new_n107), .c(new_n110), .out0(\s[6] ));
  aob012aa1n03x5               g215(.a(new_n107), .b(new_n309), .c(new_n110), .out0(new_n311));
  xnrb03aa1n02x5               g216(.a(new_n311), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g217(.a(\a[7] ), .b(\b[6] ), .c(new_n311), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g219(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


