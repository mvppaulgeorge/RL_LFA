// Benchmark "adder" written by ABC on Thu Jul 18 03:58:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n324,
    new_n327, new_n329, new_n330, new_n331, new_n332, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv020aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nor002aa1d32x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  inv040aa1n03x5               g004(.a(new_n99), .o1(new_n100));
  oaoi03aa1n09x5               g005(.a(\a[8] ), .b(\b[7] ), .c(new_n100), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nanp02aa1n06x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nona23aa1d18x5               g009(.a(new_n102), .b(new_n104), .c(new_n99), .d(new_n103), .out0(new_n105));
  inv000aa1d42x5               g010(.a(\a[6] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[5] ), .o1(new_n107));
  nor042aa1n04x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  oaoi03aa1n12x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  oabi12aa1n18x5               g014(.a(new_n101), .b(new_n105), .c(new_n109), .out0(new_n110));
  nor022aa1n04x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nand02aa1n06x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nor022aa1n12x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  nanp02aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand22aa1n09x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  nor002aa1n03x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  oai012aa1n04x7               g023(.a(new_n116), .b(new_n118), .c(new_n117), .o1(new_n119));
  tech160nm_fiaoi012aa1n03p5x5 g024(.a(new_n111), .b(new_n113), .c(new_n112), .o1(new_n120));
  oai012aa1n18x5               g025(.a(new_n120), .b(new_n115), .c(new_n119), .o1(new_n121));
  xnrc02aa1n02x5               g026(.a(\b[5] ), .b(\a[6] ), .out0(new_n122));
  tech160nm_fixnrc02aa1n04x5   g027(.a(\b[4] ), .b(\a[5] ), .out0(new_n123));
  nor043aa1n06x5               g028(.a(new_n105), .b(new_n122), .c(new_n123), .o1(new_n124));
  nand42aa1n03x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n97), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n110), .c(new_n121), .d(new_n124), .o1(new_n127));
  nor042aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanp02aa1n04x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  nor042aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n08x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n06x4               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  tech160nm_fioai012aa1n04x5   g039(.a(new_n129), .b(new_n128), .c(new_n97), .o1(new_n135));
  nano23aa1n06x5               g040(.a(new_n97), .b(new_n128), .c(new_n129), .d(new_n125), .out0(new_n136));
  aoai13aa1n02x5               g041(.a(new_n136), .b(new_n110), .c(new_n121), .d(new_n124), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n134), .b(new_n137), .c(new_n135), .out0(\s[11] ));
  inv000aa1d42x5               g043(.a(new_n110), .o1(new_n139));
  nand42aa1n02x5               g044(.a(new_n121), .b(new_n124), .o1(new_n140));
  nand22aa1n03x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  oaoi03aa1n06x5               g046(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n142));
  aoai13aa1n02x5               g047(.a(new_n134), .b(new_n142), .c(new_n141), .d(new_n136), .o1(new_n143));
  oai012aa1n02x5               g048(.a(new_n143), .b(\b[10] ), .c(\a[11] ), .o1(new_n144));
  xorb03aa1n02x5               g049(.a(new_n144), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor022aa1n08x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n16x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanb02aa1n02x5               g052(.a(new_n146), .b(new_n147), .out0(new_n148));
  nano32aa1n03x7               g053(.a(new_n148), .b(new_n134), .c(new_n130), .d(new_n126), .out0(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n110), .c(new_n121), .d(new_n124), .o1(new_n150));
  nano23aa1n03x7               g055(.a(new_n132), .b(new_n146), .c(new_n147), .d(new_n133), .out0(new_n151));
  aoi012aa1n12x5               g056(.a(new_n146), .b(new_n132), .c(new_n147), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n153), .b(new_n151), .c(new_n142), .o1(new_n154));
  nor022aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n06x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n150), .c(new_n154), .out0(\s[13] ));
  inv000aa1d42x5               g063(.a(\a[13] ), .o1(new_n159));
  inv000aa1d42x5               g064(.a(\b[12] ), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(new_n150), .b(new_n154), .o1(new_n161));
  oaoi03aa1n02x5               g066(.a(new_n159), .b(new_n160), .c(new_n161), .o1(new_n162));
  xnrb03aa1n02x5               g067(.a(new_n162), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nand42aa1n06x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nona23aa1n02x4               g070(.a(new_n165), .b(new_n156), .c(new_n155), .d(new_n164), .out0(new_n166));
  aoai13aa1n04x5               g071(.a(new_n165), .b(new_n164), .c(new_n159), .d(new_n160), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n166), .c(new_n150), .d(new_n154), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand02aa1d06x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nor002aa1n12x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  nand02aa1n06x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  aoi122aa1n06x5               g079(.a(new_n170), .b(new_n174), .c(new_n173), .d(new_n168), .e(new_n171), .o1(new_n175));
  aoi012aa1n02x5               g080(.a(new_n170), .b(new_n168), .c(new_n171), .o1(new_n176));
  nanb02aa1n06x5               g081(.a(new_n172), .b(new_n174), .out0(new_n177));
  norp02aa1n02x5               g082(.a(new_n176), .b(new_n177), .o1(new_n178));
  norp02aa1n03x5               g083(.a(new_n178), .b(new_n175), .o1(\s[16] ));
  nano23aa1n06x5               g084(.a(new_n155), .b(new_n164), .c(new_n165), .d(new_n156), .out0(new_n180));
  nano23aa1n06x5               g085(.a(new_n170), .b(new_n172), .c(new_n174), .d(new_n171), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n181), .b(new_n180), .o1(new_n182));
  nano22aa1n03x7               g087(.a(new_n182), .b(new_n136), .c(new_n151), .out0(new_n183));
  aoai13aa1n12x5               g088(.a(new_n183), .b(new_n110), .c(new_n121), .d(new_n124), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n167), .b(new_n181), .out0(new_n185));
  aoi112aa1n03x5               g090(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  nanp02aa1n02x5               g092(.a(new_n151), .b(new_n142), .o1(new_n188));
  aoi012aa1n03x5               g093(.a(new_n182), .b(new_n188), .c(new_n152), .o1(new_n189));
  nano32aa1n09x5               g094(.a(new_n189), .b(new_n187), .c(new_n185), .d(new_n173), .out0(new_n190));
  xorc02aa1n12x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n190), .c(new_n184), .out0(\s[17] ));
  nanp02aa1n09x5               g097(.a(new_n190), .b(new_n184), .o1(new_n193));
  norp02aa1n02x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  tech160nm_fiaoi012aa1n05x5   g099(.a(new_n194), .b(new_n193), .c(new_n191), .o1(new_n195));
  xnrc02aa1n06x5               g100(.a(\b[17] ), .b(\a[18] ), .out0(new_n196));
  xorc02aa1n02x5               g101(.a(new_n195), .b(new_n196), .out0(\s[18] ));
  norb02aa1n03x5               g102(.a(new_n191), .b(new_n196), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  oaih22aa1n04x5               g104(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n200));
  aob012aa1n06x5               g105(.a(new_n200), .b(\b[17] ), .c(\a[18] ), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n199), .c(new_n190), .d(new_n184), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  xnrc02aa1n12x5               g110(.a(\b[18] ), .b(\a[19] ), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  xnrc02aa1n12x5               g112(.a(\b[19] ), .b(\a[20] ), .out0(new_n208));
  inv020aa1n06x5               g113(.a(new_n208), .o1(new_n209));
  aoi112aa1n03x4               g114(.a(new_n205), .b(new_n209), .c(new_n202), .d(new_n207), .o1(new_n210));
  inv000aa1n02x5               g115(.a(new_n205), .o1(new_n211));
  nand02aa1n02x5               g116(.a(new_n202), .b(new_n207), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n208), .b(new_n212), .c(new_n211), .o1(new_n213));
  norp02aa1n03x5               g118(.a(new_n213), .b(new_n210), .o1(\s[20] ));
  nona23aa1n09x5               g119(.a(new_n191), .b(new_n209), .c(new_n206), .d(new_n196), .out0(new_n215));
  oao003aa1n02x5               g120(.a(\a[20] ), .b(\b[19] ), .c(new_n211), .carry(new_n216));
  oai013aa1d12x5               g121(.a(new_n216), .b(new_n201), .c(new_n206), .d(new_n208), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n215), .c(new_n190), .d(new_n184), .o1(new_n219));
  xorb03aa1n02x5               g124(.a(new_n219), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  xorc02aa1n02x5               g126(.a(\a[21] ), .b(\b[20] ), .out0(new_n222));
  xorc02aa1n12x5               g127(.a(\a[22] ), .b(\b[21] ), .out0(new_n223));
  aoi112aa1n03x4               g128(.a(new_n221), .b(new_n223), .c(new_n219), .d(new_n222), .o1(new_n224));
  inv000aa1n02x5               g129(.a(new_n221), .o1(new_n225));
  nand02aa1n02x5               g130(.a(new_n219), .b(new_n222), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n223), .o1(new_n227));
  aoi012aa1n06x5               g132(.a(new_n227), .b(new_n226), .c(new_n225), .o1(new_n228));
  nor002aa1n02x5               g133(.a(new_n228), .b(new_n224), .o1(\s[22] ));
  inv000aa1d42x5               g134(.a(\a[21] ), .o1(new_n230));
  inv040aa1d32x5               g135(.a(\a[22] ), .o1(new_n231));
  xroi22aa1d04x5               g136(.a(new_n230), .b(\b[20] ), .c(new_n231), .d(\b[21] ), .out0(new_n232));
  oaoi03aa1n02x5               g137(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .o1(new_n233));
  aoi012aa1n02x7               g138(.a(new_n233), .b(new_n217), .c(new_n232), .o1(new_n234));
  nona23aa1n02x4               g139(.a(new_n198), .b(new_n232), .c(new_n208), .d(new_n206), .out0(new_n235));
  aoai13aa1n04x5               g140(.a(new_n234), .b(new_n235), .c(new_n190), .d(new_n184), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  xorc02aa1n12x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xorc02aa1n12x5               g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  aoi112aa1n03x4               g145(.a(new_n238), .b(new_n240), .c(new_n236), .d(new_n239), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n238), .o1(new_n242));
  nanp02aa1n03x5               g147(.a(new_n236), .b(new_n239), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n240), .o1(new_n244));
  aoi012aa1n06x5               g149(.a(new_n244), .b(new_n243), .c(new_n242), .o1(new_n245));
  nor002aa1n02x5               g150(.a(new_n245), .b(new_n241), .o1(\s[24] ));
  nanp02aa1n02x5               g151(.a(new_n223), .b(new_n222), .o1(new_n247));
  nano22aa1n02x4               g152(.a(new_n247), .b(new_n239), .c(new_n240), .out0(new_n248));
  nanb02aa1n03x5               g153(.a(new_n215), .b(new_n248), .out0(new_n249));
  nona22aa1n03x5               g154(.a(new_n209), .b(new_n201), .c(new_n206), .out0(new_n250));
  inv000aa1d42x5               g155(.a(\a[23] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\a[24] ), .o1(new_n252));
  xroi22aa1d04x5               g157(.a(new_n251), .b(\b[22] ), .c(new_n252), .d(\b[23] ), .out0(new_n253));
  nand22aa1n04x5               g158(.a(new_n253), .b(new_n232), .o1(new_n254));
  oaoi03aa1n02x5               g159(.a(\a[24] ), .b(\b[23] ), .c(new_n242), .o1(new_n255));
  aoi013aa1n06x4               g160(.a(new_n255), .b(new_n233), .c(new_n239), .d(new_n240), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n254), .c(new_n250), .d(new_n216), .o1(new_n257));
  inv020aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n249), .c(new_n190), .d(new_n184), .o1(new_n259));
  xorb03aa1n02x5               g164(.a(new_n259), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xorc02aa1n12x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  aoi112aa1n03x4               g168(.a(new_n261), .b(new_n263), .c(new_n259), .d(new_n262), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n261), .o1(new_n265));
  nanp02aa1n03x5               g170(.a(new_n259), .b(new_n262), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n263), .o1(new_n267));
  tech160nm_fiaoi012aa1n05x5   g172(.a(new_n267), .b(new_n266), .c(new_n265), .o1(new_n268));
  norp02aa1n03x5               g173(.a(new_n268), .b(new_n264), .o1(\s[26] ));
  nanb02aa1n02x5               g174(.a(new_n170), .b(new_n171), .out0(new_n270));
  norp03aa1n02x5               g175(.a(new_n167), .b(new_n177), .c(new_n270), .o1(new_n271));
  norb03aa1n02x5               g176(.a(new_n134), .b(new_n135), .c(new_n148), .out0(new_n272));
  nor043aa1n03x5               g177(.a(new_n166), .b(new_n177), .c(new_n270), .o1(new_n273));
  oai012aa1n02x5               g178(.a(new_n273), .b(new_n272), .c(new_n153), .o1(new_n274));
  nona32aa1n03x5               g179(.a(new_n274), .b(new_n186), .c(new_n271), .d(new_n172), .out0(new_n275));
  and002aa1n12x5               g180(.a(new_n263), .b(new_n262), .o(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  nor043aa1n06x5               g182(.a(new_n277), .b(new_n254), .c(new_n215), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n275), .c(new_n141), .d(new_n183), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .c(new_n265), .carry(new_n280));
  aobi12aa1n06x5               g185(.a(new_n280), .b(new_n257), .c(new_n276), .out0(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n279), .c(new_n281), .out0(\s[27] ));
  nor042aa1n03x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n282), .o1(new_n286));
  tech160nm_fiaoi012aa1n02p5x5 g191(.a(new_n286), .b(new_n279), .c(new_n281), .o1(new_n287));
  xnrc02aa1n12x5               g192(.a(\b[27] ), .b(\a[28] ), .out0(new_n288));
  nano22aa1n03x5               g193(.a(new_n287), .b(new_n285), .c(new_n288), .out0(new_n289));
  nand02aa1n04x5               g194(.a(new_n217), .b(new_n248), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n280), .b(new_n277), .c(new_n290), .d(new_n256), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n282), .b(new_n291), .c(new_n193), .d(new_n278), .o1(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n288), .b(new_n292), .c(new_n285), .o1(new_n293));
  norp02aa1n03x5               g198(.a(new_n293), .b(new_n289), .o1(\s[28] ));
  norb02aa1d21x5               g199(.a(new_n282), .b(new_n288), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n291), .c(new_n193), .d(new_n278), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[28] ), .b(\a[29] ), .out0(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n298), .b(new_n296), .c(new_n297), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n295), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n279), .c(new_n281), .o1(new_n301));
  nano22aa1n03x5               g206(.a(new_n301), .b(new_n297), .c(new_n298), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n299), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n09x5               g209(.a(new_n282), .b(new_n298), .c(new_n288), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n291), .c(new_n193), .d(new_n278), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n305), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n310), .b(new_n279), .c(new_n281), .o1(new_n311));
  nano22aa1n02x4               g216(.a(new_n311), .b(new_n307), .c(new_n308), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n309), .b(new_n312), .o1(\s[30] ));
  norb02aa1n03x5               g218(.a(new_n305), .b(new_n308), .out0(new_n314));
  inv020aa1n02x5               g219(.a(new_n314), .o1(new_n315));
  tech160nm_fiaoi012aa1n02p5x5 g220(.a(new_n315), .b(new_n279), .c(new_n281), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  nano22aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n318), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n314), .b(new_n291), .c(new_n193), .d(new_n278), .o1(new_n320));
  tech160nm_fiaoi012aa1n02p5x5 g225(.a(new_n318), .b(new_n320), .c(new_n317), .o1(new_n321));
  nor002aa1n02x5               g226(.a(new_n321), .b(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g227(.a(new_n119), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g228(.a(\a[3] ), .b(\b[2] ), .c(new_n119), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoib12aa1n06x5               g231(.a(new_n108), .b(new_n121), .c(new_n123), .out0(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(new_n106), .out0(\s[6] ));
  norb02aa1n02x5               g233(.a(new_n104), .b(new_n99), .out0(new_n329));
  nanb02aa1n02x5               g234(.a(new_n122), .b(new_n327), .out0(new_n330));
  oai112aa1n03x5               g235(.a(new_n330), .b(new_n329), .c(new_n107), .d(new_n106), .o1(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n329), .b(new_n330), .c(new_n106), .d(new_n107), .o1(new_n332));
  norb02aa1n02x5               g237(.a(new_n331), .b(new_n332), .out0(\s[7] ));
  norb02aa1n02x5               g238(.a(new_n102), .b(new_n103), .out0(new_n334));
  xnbna2aa1n03x5               g239(.a(new_n334), .b(new_n331), .c(new_n100), .out0(\s[8] ));
  xnbna2aa1n03x5               g240(.a(new_n126), .b(new_n140), .c(new_n139), .out0(\s[9] ));
endmodule


