// Benchmark "adder" written by ABC on Wed Jul 17 18:48:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n343, new_n344, new_n347,
    new_n348, new_n350, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .o(new_n97));
  nanp02aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nor042aa1n06x5               g003(.a(\b[8] ), .b(\a[9] ), .o1(new_n99));
  and002aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o(new_n100));
  oaoi03aa1n02x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  nor022aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand22aa1n06x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n02x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor022aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n02x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nanp03aa1n02x5               g012(.a(new_n101), .b(new_n104), .c(new_n107), .o1(new_n108));
  aoi012aa1n02x7               g013(.a(new_n102), .b(new_n105), .c(new_n103), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nand22aa1n03x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor002aa1n03x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nano23aa1n02x4               g018(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n114));
  nor002aa1n03x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  nor042aa1n03x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand02aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nanb02aa1n03x5               g024(.a(new_n118), .b(new_n119), .out0(new_n120));
  nona22aa1n02x4               g025(.a(new_n114), .b(new_n117), .c(new_n120), .out0(new_n121));
  inv000aa1n02x5               g026(.a(new_n115), .o1(new_n122));
  aoi112aa1n06x5               g027(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n123), .o1(new_n124));
  oai022aa1n02x5               g029(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n125));
  nanb03aa1n02x5               g030(.a(new_n118), .b(new_n119), .c(new_n111), .out0(new_n126));
  nano32aa1n02x4               g031(.a(new_n126), .b(new_n125), .c(new_n122), .d(new_n116), .out0(new_n127));
  nano22aa1n03x7               g032(.a(new_n127), .b(new_n122), .c(new_n124), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n121), .c(new_n108), .d(new_n109), .o1(new_n129));
  nanp02aa1n04x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  aoi012aa1n02x5               g035(.a(new_n99), .b(new_n129), .c(new_n130), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n97), .c(new_n98), .out0(\s[10] ));
  nor042aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  inv000aa1n02x5               g038(.a(new_n98), .o1(new_n134));
  norb02aa1n15x5               g039(.a(new_n130), .b(new_n99), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nona32aa1n02x4               g041(.a(new_n129), .b(new_n136), .c(new_n134), .d(new_n133), .out0(new_n137));
  aoi012aa1n06x5               g042(.a(new_n133), .b(new_n99), .c(new_n98), .o1(new_n138));
  nor042aa1d18x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1n02x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  xobna2aa1n03x5               g046(.a(new_n141), .b(new_n137), .c(new_n138), .out0(\s[11] ));
  inv000aa1d42x5               g047(.a(new_n139), .o1(new_n143));
  aoai13aa1n03x5               g048(.a(new_n143), .b(new_n141), .c(new_n137), .d(new_n138), .o1(new_n144));
  xorb03aa1n02x5               g049(.a(new_n144), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv000aa1d42x5               g050(.a(\a[1] ), .o1(new_n146));
  inv000aa1d42x5               g051(.a(\b[0] ), .o1(new_n147));
  nor002aa1n02x5               g052(.a(\b[1] ), .b(\a[2] ), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(\b[1] ), .b(\a[2] ), .o1(new_n149));
  oaoi13aa1n04x5               g054(.a(new_n148), .b(new_n149), .c(new_n146), .d(new_n147), .o1(new_n150));
  nona23aa1n03x5               g055(.a(new_n106), .b(new_n103), .c(new_n102), .d(new_n105), .out0(new_n151));
  tech160nm_fioai012aa1n04x5   g056(.a(new_n109), .b(new_n151), .c(new_n150), .o1(new_n152));
  nona23aa1n02x4               g057(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n153));
  nor043aa1n04x5               g058(.a(new_n153), .b(new_n117), .c(new_n120), .o1(new_n154));
  norb02aa1n06x4               g059(.a(new_n116), .b(new_n115), .out0(new_n155));
  nano22aa1n03x7               g060(.a(new_n118), .b(new_n111), .c(new_n119), .out0(new_n156));
  nand03aa1n02x5               g061(.a(new_n156), .b(new_n155), .c(new_n125), .o1(new_n157));
  nona22aa1d18x5               g062(.a(new_n157), .b(new_n123), .c(new_n115), .out0(new_n158));
  nona32aa1n09x5               g063(.a(new_n135), .b(new_n134), .c(new_n139), .d(new_n133), .out0(new_n159));
  nor042aa1n06x5               g064(.a(\b[11] ), .b(\a[12] ), .o1(new_n160));
  nanp02aa1n04x5               g065(.a(\b[11] ), .b(\a[12] ), .o1(new_n161));
  nano22aa1n02x4               g066(.a(new_n160), .b(new_n140), .c(new_n161), .out0(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n159), .out0(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n158), .c(new_n152), .d(new_n154), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n160), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(new_n139), .b(new_n161), .o1(new_n166));
  nano32aa1n02x4               g071(.a(new_n138), .b(new_n161), .c(new_n143), .d(new_n140), .out0(new_n167));
  nano22aa1n06x5               g072(.a(new_n167), .b(new_n165), .c(new_n166), .out0(new_n168));
  nor002aa1n03x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  and002aa1n02x5               g074(.a(\b[12] ), .b(\a[13] ), .o(new_n170));
  norp02aa1n02x5               g075(.a(new_n170), .b(new_n169), .o1(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n164), .c(new_n168), .out0(\s[13] ));
  orn002aa1n02x5               g077(.a(\a[13] ), .b(\b[12] ), .o(new_n173));
  aoai13aa1n02x7               g078(.a(new_n161), .b(new_n133), .c(new_n99), .d(new_n98), .o1(new_n174));
  oai112aa1n03x5               g079(.a(new_n166), .b(new_n165), .c(new_n174), .d(new_n141), .o1(new_n175));
  aoai13aa1n02x5               g080(.a(new_n171), .b(new_n175), .c(new_n129), .d(new_n163), .o1(new_n176));
  norp02aa1n04x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nanp02aa1n06x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  norb02aa1n06x4               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n176), .c(new_n173), .out0(\s[14] ));
  nona22aa1n02x4               g085(.a(new_n179), .b(new_n170), .c(new_n169), .out0(new_n181));
  aoi012aa1n02x5               g086(.a(new_n177), .b(new_n169), .c(new_n178), .o1(new_n182));
  aoai13aa1n03x5               g087(.a(new_n182), .b(new_n181), .c(new_n164), .d(new_n168), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  nand02aa1n04x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  nanb02aa1n12x5               g092(.a(new_n185), .b(new_n187), .out0(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n183), .b(new_n189), .o1(new_n190));
  nor042aa1n06x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nand22aa1n02x5               g096(.a(\b[15] ), .b(\a[16] ), .o1(new_n192));
  norb02aa1n09x5               g097(.a(new_n192), .b(new_n191), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  aoi012aa1n06x5               g099(.a(new_n194), .b(new_n190), .c(new_n186), .o1(new_n195));
  aoi112aa1n02x5               g100(.a(new_n185), .b(new_n193), .c(new_n183), .d(new_n187), .o1(new_n196));
  norp02aa1n02x5               g101(.a(new_n195), .b(new_n196), .o1(\s[16] ));
  nona32aa1n02x4               g102(.a(new_n179), .b(new_n170), .c(new_n185), .d(new_n169), .out0(new_n198));
  nano22aa1n03x5               g103(.a(new_n191), .b(new_n187), .c(new_n192), .out0(new_n199));
  nano23aa1n06x5               g104(.a(new_n159), .b(new_n198), .c(new_n199), .d(new_n162), .out0(new_n200));
  aoai13aa1n12x5               g105(.a(new_n200), .b(new_n158), .c(new_n152), .d(new_n154), .o1(new_n201));
  nano32aa1n03x7               g106(.a(new_n181), .b(new_n193), .c(new_n186), .d(new_n187), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n191), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n185), .b(new_n192), .o1(new_n204));
  aoai13aa1n02x5               g109(.a(new_n192), .b(new_n177), .c(new_n169), .d(new_n178), .o1(new_n205));
  oai112aa1n04x5               g110(.a(new_n204), .b(new_n203), .c(new_n205), .d(new_n188), .o1(new_n206));
  aoi012aa1n09x5               g111(.a(new_n206), .b(new_n175), .c(new_n202), .o1(new_n207));
  nanp02aa1n09x5               g112(.a(new_n201), .b(new_n207), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g114(.a(\a[18] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(\a[17] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(\b[16] ), .o1(new_n212));
  oaoi03aa1n03x5               g117(.a(new_n211), .b(new_n212), .c(new_n208), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[17] ), .c(new_n210), .out0(\s[18] ));
  xroi22aa1d06x4               g119(.a(new_n211), .b(\b[16] ), .c(new_n210), .d(\b[17] ), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  norp02aa1n02x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  aoi013aa1n06x4               g123(.a(new_n217), .b(new_n218), .c(new_n211), .d(new_n212), .o1(new_n219));
  aoai13aa1n04x5               g124(.a(new_n219), .b(new_n216), .c(new_n201), .d(new_n207), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g127(.a(\a[19] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[18] ), .o1(new_n224));
  nand02aa1d08x5               g129(.a(new_n224), .b(new_n223), .o1(new_n225));
  nand02aa1n04x5               g130(.a(\b[18] ), .b(\a[19] ), .o1(new_n226));
  nanp02aa1n02x5               g131(.a(new_n225), .b(new_n226), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(new_n220), .b(new_n228), .o1(new_n229));
  nor042aa1n04x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nanp02aa1n02x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  norb02aa1n09x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv040aa1n02x5               g137(.a(new_n232), .o1(new_n233));
  tech160nm_fiaoi012aa1n02p5x5 g138(.a(new_n233), .b(new_n229), .c(new_n225), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n225), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n235), .b(new_n232), .c(new_n220), .d(new_n226), .o1(new_n236));
  nor002aa1n02x5               g141(.a(new_n234), .b(new_n236), .o1(\s[20] ));
  nona23aa1d18x5               g142(.a(new_n215), .b(new_n226), .c(new_n233), .d(new_n235), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n230), .o1(new_n239));
  aoi112aa1n09x5               g144(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  nano32aa1n02x4               g146(.a(new_n219), .b(new_n231), .c(new_n225), .d(new_n226), .out0(new_n242));
  nano22aa1n03x5               g147(.a(new_n242), .b(new_n239), .c(new_n241), .out0(new_n243));
  aoai13aa1n04x5               g148(.a(new_n243), .b(new_n238), .c(new_n201), .d(new_n207), .o1(new_n244));
  xorb03aa1n02x5               g149(.a(new_n244), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[21] ), .b(\b[20] ), .out0(new_n248));
  nanp02aa1n02x5               g153(.a(new_n244), .b(new_n248), .o1(new_n249));
  xnrc02aa1n02x5               g154(.a(\b[21] ), .b(\a[22] ), .out0(new_n250));
  tech160nm_fiaoi012aa1n02p5x5 g155(.a(new_n250), .b(new_n249), .c(new_n247), .o1(new_n251));
  tech160nm_fixorc02aa1n05x5   g156(.a(\a[22] ), .b(\b[21] ), .out0(new_n252));
  aoi112aa1n02x5               g157(.a(new_n246), .b(new_n252), .c(new_n244), .d(new_n248), .o1(new_n253));
  nor002aa1n02x5               g158(.a(new_n251), .b(new_n253), .o1(\s[22] ));
  nand02aa1n08x5               g159(.a(new_n252), .b(new_n248), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  nanb02aa1n03x5               g161(.a(new_n238), .b(new_n256), .out0(new_n257));
  oaoi03aa1n03x5               g162(.a(\a[22] ), .b(\b[21] ), .c(new_n247), .o1(new_n258));
  oab012aa1n02x4               g163(.a(new_n258), .b(new_n243), .c(new_n255), .out0(new_n259));
  aoai13aa1n04x5               g164(.a(new_n259), .b(new_n257), .c(new_n201), .d(new_n207), .o1(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n12x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n264), .b(new_n262), .out0(new_n265));
  nand02aa1n02x5               g170(.a(new_n260), .b(new_n265), .o1(new_n266));
  norp02aa1n02x5               g171(.a(\b[23] ), .b(\a[24] ), .o1(new_n267));
  nanp02aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .o1(new_n268));
  norb02aa1n02x5               g173(.a(new_n268), .b(new_n267), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  tech160nm_fiaoi012aa1n03p5x5 g175(.a(new_n270), .b(new_n266), .c(new_n263), .o1(new_n271));
  aoi112aa1n03x4               g176(.a(new_n262), .b(new_n269), .c(new_n260), .d(new_n264), .o1(new_n272));
  nor042aa1n03x5               g177(.a(new_n271), .b(new_n272), .o1(\s[24] ));
  nano22aa1n03x7               g178(.a(new_n267), .b(new_n264), .c(new_n268), .out0(new_n274));
  nano22aa1n03x7               g179(.a(new_n255), .b(new_n263), .c(new_n274), .out0(new_n275));
  nanb02aa1n03x5               g180(.a(new_n238), .b(new_n275), .out0(new_n276));
  nona23aa1n09x5               g181(.a(new_n274), .b(new_n248), .c(new_n250), .d(new_n262), .out0(new_n277));
  aoi112aa1n02x5               g182(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n278));
  aoi113aa1n02x5               g183(.a(new_n278), .b(new_n267), .c(new_n258), .d(new_n268), .e(new_n265), .o1(new_n279));
  oa0012aa1n02x5               g184(.a(new_n279), .b(new_n243), .c(new_n277), .o(new_n280));
  aoai13aa1n04x5               g185(.a(new_n280), .b(new_n276), .c(new_n201), .d(new_n207), .o1(new_n281));
  xorb03aa1n02x5               g186(.a(new_n281), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  nand02aa1n02x5               g190(.a(new_n281), .b(new_n285), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[26] ), .b(\b[25] ), .out0(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  tech160nm_fiaoi012aa1n03p5x5 g193(.a(new_n288), .b(new_n286), .c(new_n284), .o1(new_n289));
  aoi112aa1n03x4               g194(.a(new_n283), .b(new_n287), .c(new_n281), .d(new_n285), .o1(new_n290));
  nor002aa1n02x5               g195(.a(new_n289), .b(new_n290), .o1(\s[26] ));
  nanb02aa1n02x5               g196(.a(new_n177), .b(new_n178), .out0(new_n292));
  nona23aa1n02x4               g197(.a(new_n199), .b(new_n171), .c(new_n292), .d(new_n185), .out0(new_n293));
  oabi12aa1n02x5               g198(.a(new_n206), .b(new_n168), .c(new_n293), .out0(new_n294));
  nanp02aa1n02x5               g199(.a(new_n287), .b(new_n285), .o1(new_n295));
  nor043aa1d12x5               g200(.a(new_n238), .b(new_n277), .c(new_n295), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n294), .c(new_n129), .d(new_n200), .o1(new_n297));
  oaoi13aa1n02x7               g202(.a(new_n295), .b(new_n279), .c(new_n243), .d(new_n277), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[26] ), .b(\b[25] ), .c(new_n284), .carry(new_n299));
  norb02aa1n03x5               g204(.a(new_n299), .b(new_n298), .out0(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  xnbna2aa1n03x5               g206(.a(new_n301), .b(new_n300), .c(new_n297), .out0(\s[27] ));
  nor042aa1n03x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  oai013aa1n02x4               g209(.a(new_n275), .b(new_n242), .c(new_n230), .d(new_n240), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n299), .b(new_n295), .c(new_n305), .d(new_n279), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n301), .b(new_n306), .c(new_n208), .d(new_n296), .o1(new_n307));
  tech160nm_fixnrc02aa1n04x5   g212(.a(\b[27] ), .b(\a[28] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n307), .c(new_n304), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n301), .o1(new_n310));
  aoi012aa1n02x7               g215(.a(new_n310), .b(new_n300), .c(new_n297), .o1(new_n311));
  nano22aa1n03x5               g216(.a(new_n311), .b(new_n304), .c(new_n308), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n309), .b(new_n312), .o1(\s[28] ));
  norb02aa1d21x5               g218(.a(new_n301), .b(new_n308), .out0(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n306), .c(new_n208), .d(new_n296), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n316));
  xnrc02aa1n02x5               g221(.a(\b[28] ), .b(\a[29] ), .out0(new_n317));
  tech160nm_fiaoi012aa1n02p5x5 g222(.a(new_n317), .b(new_n315), .c(new_n316), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n314), .o1(new_n319));
  aoi012aa1n02x7               g224(.a(new_n319), .b(new_n300), .c(new_n297), .o1(new_n320));
  nano22aa1n03x5               g225(.a(new_n320), .b(new_n316), .c(new_n317), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n318), .b(new_n321), .o1(\s[29] ));
  xnrb03aa1n02x5               g227(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n06x5               g228(.a(new_n301), .b(new_n317), .c(new_n308), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n306), .c(new_n208), .d(new_n296), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .carry(new_n326));
  xnrc02aa1n02x5               g231(.a(\b[29] ), .b(\a[30] ), .out0(new_n327));
  tech160nm_fiaoi012aa1n02p5x5 g232(.a(new_n327), .b(new_n325), .c(new_n326), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n324), .o1(new_n329));
  aoi012aa1n02x7               g234(.a(new_n329), .b(new_n300), .c(new_n297), .o1(new_n330));
  nano22aa1n03x5               g235(.a(new_n330), .b(new_n326), .c(new_n327), .out0(new_n331));
  norp02aa1n03x5               g236(.a(new_n328), .b(new_n331), .o1(\s[30] ));
  norb02aa1n06x5               g237(.a(new_n324), .b(new_n327), .out0(new_n333));
  inv000aa1n02x5               g238(.a(new_n333), .o1(new_n334));
  aoi012aa1n02x7               g239(.a(new_n334), .b(new_n300), .c(new_n297), .o1(new_n335));
  oao003aa1n02x5               g240(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n336));
  xnrc02aa1n02x5               g241(.a(\b[30] ), .b(\a[31] ), .out0(new_n337));
  nano22aa1n03x5               g242(.a(new_n335), .b(new_n336), .c(new_n337), .out0(new_n338));
  aoai13aa1n03x5               g243(.a(new_n333), .b(new_n306), .c(new_n208), .d(new_n296), .o1(new_n339));
  tech160nm_fiaoi012aa1n02p5x5 g244(.a(new_n337), .b(new_n339), .c(new_n336), .o1(new_n340));
  norp02aa1n03x5               g245(.a(new_n340), .b(new_n338), .o1(\s[31] ));
  xnrc02aa1n02x5               g246(.a(new_n150), .b(new_n107), .out0(\s[3] ));
  obai22aa1n02x7               g247(.a(new_n103), .b(new_n102), .c(\a[3] ), .d(\b[2] ), .out0(new_n343));
  aoi012aa1n02x5               g248(.a(new_n343), .b(new_n101), .c(new_n107), .o1(new_n344));
  oaoi13aa1n02x5               g249(.a(new_n344), .b(new_n152), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g250(.a(new_n152), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g251(.a(\a[6] ), .o1(new_n347));
  aoi012aa1n02x5               g252(.a(new_n112), .b(new_n152), .c(new_n113), .o1(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[5] ), .c(new_n347), .out0(\s[6] ));
  oaib12aa1n02x5               g254(.a(new_n348), .b(\b[5] ), .c(new_n347), .out0(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n120), .b(new_n350), .c(new_n111), .out0(\s[7] ));
  aoi012aa1n02x5               g256(.a(new_n118), .b(new_n350), .c(new_n156), .o1(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n352), .b(new_n122), .c(new_n116), .out0(\s[8] ));
  xorb03aa1n02x5               g258(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


