// Benchmark "adder" written by ABC on Wed Jul 17 19:02:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n330, new_n332, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n04x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  inv000aa1n02x5               g003(.a(new_n98), .o1(new_n99));
  nand22aa1n03x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aob012aa1n02x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  nor002aa1n03x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n02x7               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor002aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n02x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nanp03aa1n06x5               g013(.a(new_n102), .b(new_n105), .c(new_n108), .o1(new_n109));
  tech160nm_fiaoi012aa1n03p5x5 g014(.a(new_n103), .b(new_n106), .c(new_n104), .o1(new_n110));
  norp02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor042aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nano23aa1n02x4               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  norp02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano23aa1n02x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nanp02aa1n02x5               g025(.a(new_n120), .b(new_n115), .o1(new_n121));
  norb02aa1n03x5               g026(.a(new_n114), .b(new_n113), .out0(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  aoi022aa1n02x5               g028(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n124));
  oa0012aa1n02x5               g029(.a(new_n112), .b(new_n113), .c(new_n111), .o(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n122), .c(new_n123), .d(new_n124), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n126), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n127));
  nand42aa1n03x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  aoi012aa1n02x5               g033(.a(new_n97), .b(new_n127), .c(new_n128), .o1(new_n129));
  xnrb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1n03x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  xorc02aa1n12x5               g036(.a(\a[11] ), .b(\b[10] ), .out0(new_n132));
  norb02aa1n06x4               g037(.a(new_n128), .b(new_n97), .out0(new_n133));
  norp02aa1n02x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  norp02aa1n02x5               g039(.a(new_n134), .b(new_n97), .o1(new_n135));
  aob012aa1n02x5               g040(.a(new_n135), .b(new_n127), .c(new_n133), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n132), .b(new_n136), .c(new_n131), .out0(\s[11] ));
  orn002aa1n02x5               g042(.a(\a[11] ), .b(\b[10] ), .o(new_n138));
  oai022aa1n02x5               g043(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n139));
  and002aa1n02x5               g044(.a(new_n132), .b(new_n131), .o(new_n140));
  aoai13aa1n02x5               g045(.a(new_n140), .b(new_n139), .c(new_n127), .d(new_n133), .o1(new_n141));
  xnrc02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .out0(new_n142));
  xobna2aa1n03x5               g047(.a(new_n142), .b(new_n141), .c(new_n138), .out0(\s[12] ));
  aoi012aa1n02x5               g048(.a(new_n98), .b(new_n100), .c(new_n101), .o1(new_n144));
  nona23aa1n02x4               g049(.a(new_n107), .b(new_n104), .c(new_n103), .d(new_n106), .out0(new_n145));
  tech160nm_fioai012aa1n03p5x5 g050(.a(new_n110), .b(new_n145), .c(new_n144), .o1(new_n146));
  nanb02aa1n06x5               g051(.a(new_n121), .b(new_n146), .out0(new_n147));
  nanb02aa1n02x5               g052(.a(new_n134), .b(new_n131), .out0(new_n148));
  nona23aa1n03x5               g053(.a(new_n132), .b(new_n133), .c(new_n142), .d(new_n148), .out0(new_n149));
  aoi022aa1n02x5               g054(.a(\b[9] ), .b(\a[10] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n150));
  oaoi03aa1n02x5               g055(.a(\a[12] ), .b(\b[11] ), .c(new_n138), .o1(new_n151));
  aoi013aa1n02x4               g056(.a(new_n151), .b(new_n132), .c(new_n139), .d(new_n150), .o1(new_n152));
  aoai13aa1n03x5               g057(.a(new_n152), .b(new_n149), .c(new_n147), .d(new_n126), .o1(new_n153));
  norp02aa1n03x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand42aa1n03x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  nano23aa1n03x5               g061(.a(new_n148), .b(new_n142), .c(new_n132), .d(new_n133), .out0(new_n157));
  nanp03aa1n02x5               g062(.a(new_n132), .b(new_n139), .c(new_n150), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n151), .b(new_n158), .out0(new_n159));
  aoi112aa1n02x5               g064(.a(new_n156), .b(new_n159), .c(new_n127), .d(new_n157), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n160), .b(new_n153), .c(new_n156), .o1(\s[13] ));
  inv000aa1d42x5               g066(.a(\a[13] ), .o1(new_n162));
  inv000aa1d42x5               g067(.a(\b[12] ), .o1(new_n163));
  oaoi03aa1n03x5               g068(.a(new_n162), .b(new_n163), .c(new_n153), .o1(new_n164));
  xnrb03aa1n03x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n12x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nand42aa1n10x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nona23aa1d18x5               g072(.a(new_n167), .b(new_n155), .c(new_n154), .d(new_n166), .out0(new_n168));
  inv000aa1n02x5               g073(.a(new_n168), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n159), .c(new_n127), .d(new_n157), .o1(new_n170));
  aoai13aa1n12x5               g075(.a(new_n167), .b(new_n166), .c(new_n162), .d(new_n163), .o1(new_n171));
  norp02aa1n03x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n04x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n171), .out0(\s[15] ));
  inv000aa1n02x5               g080(.a(new_n172), .o1(new_n176));
  inv000aa1n02x5               g081(.a(new_n173), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n176), .b(new_n177), .c(new_n170), .d(new_n171), .o1(new_n178));
  nor022aa1n08x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand42aa1n03x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n178), .b(new_n181), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n171), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n174), .b(new_n183), .c(new_n153), .d(new_n169), .o1(new_n184));
  nona22aa1n02x4               g089(.a(new_n184), .b(new_n181), .c(new_n172), .out0(new_n185));
  nanp02aa1n02x5               g090(.a(new_n182), .b(new_n185), .o1(\s[16] ));
  nona23aa1n03x5               g091(.a(new_n180), .b(new_n173), .c(new_n172), .d(new_n179), .out0(new_n187));
  norp02aa1n06x5               g092(.a(new_n187), .b(new_n168), .o1(new_n188));
  norb02aa1n06x5               g093(.a(new_n188), .b(new_n149), .out0(new_n189));
  nand22aa1n03x5               g094(.a(new_n127), .b(new_n189), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n179), .o1(new_n191));
  aoai13aa1n09x5               g096(.a(new_n191), .b(new_n177), .c(new_n171), .d(new_n176), .o1(new_n192));
  aoi022aa1n06x5               g097(.a(new_n159), .b(new_n188), .c(new_n192), .d(new_n180), .o1(new_n193));
  xorc02aa1n02x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n190), .c(new_n193), .out0(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  nand02aa1n02x5               g101(.a(new_n157), .b(new_n188), .o1(new_n197));
  aoai13aa1n06x5               g102(.a(new_n193), .b(new_n197), .c(new_n147), .d(new_n126), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  tech160nm_fiaoi012aa1n05x5   g104(.a(new_n199), .b(new_n198), .c(new_n194), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n196), .out0(\s[18] ));
  nona32aa1n02x4               g106(.a(new_n169), .b(new_n181), .c(new_n177), .d(new_n172), .out0(new_n202));
  nand42aa1n02x5               g107(.a(new_n192), .b(new_n180), .o1(new_n203));
  oai012aa1n06x5               g108(.a(new_n203), .b(new_n202), .c(new_n152), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\a[17] ), .o1(new_n205));
  xroi22aa1d06x4               g110(.a(new_n205), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n204), .c(new_n127), .d(new_n189), .o1(new_n207));
  nand42aa1n03x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  oai022aa1d24x5               g113(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n209));
  nanp02aa1n02x5               g114(.a(new_n209), .b(new_n208), .o1(new_n210));
  nor042aa1n02x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanp02aa1n04x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n09x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n207), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g120(.a(new_n207), .b(new_n210), .o1(new_n216));
  xnrc02aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .out0(new_n217));
  aoai13aa1n02x5               g122(.a(new_n217), .b(new_n211), .c(new_n216), .d(new_n212), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n210), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n213), .b(new_n219), .c(new_n198), .d(new_n206), .o1(new_n220));
  nona22aa1n02x4               g125(.a(new_n220), .b(new_n217), .c(new_n211), .out0(new_n221));
  nanp02aa1n02x5               g126(.a(new_n218), .b(new_n221), .o1(\s[20] ));
  nanb03aa1d18x5               g127(.a(new_n217), .b(new_n206), .c(new_n213), .out0(new_n223));
  aoi013aa1n06x4               g128(.a(new_n211), .b(new_n209), .c(new_n208), .d(new_n212), .o1(new_n224));
  oaoi03aa1n12x5               g129(.a(\a[20] ), .b(\b[19] ), .c(new_n224), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n223), .c(new_n190), .d(new_n193), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  nanp02aa1n02x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  norp02aa1n02x5               g136(.a(\b[21] ), .b(\a[22] ), .o1(new_n232));
  nanp02aa1n04x5               g137(.a(\b[21] ), .b(\a[22] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n02x7               g140(.a(new_n235), .b(new_n229), .c(new_n227), .d(new_n231), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n223), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n231), .b(new_n225), .c(new_n198), .d(new_n237), .o1(new_n238));
  nona22aa1n02x4               g143(.a(new_n238), .b(new_n235), .c(new_n229), .out0(new_n239));
  nanp02aa1n02x5               g144(.a(new_n236), .b(new_n239), .o1(\s[22] ));
  nano23aa1n06x5               g145(.a(new_n229), .b(new_n232), .c(new_n233), .d(new_n230), .out0(new_n241));
  nano32aa1n02x4               g146(.a(new_n217), .b(new_n206), .c(new_n241), .d(new_n213), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n204), .c(new_n127), .d(new_n189), .o1(new_n243));
  oaih22aa1n06x5               g148(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n244));
  aoi022aa1n06x5               g149(.a(new_n225), .b(new_n241), .c(new_n233), .d(new_n244), .o1(new_n245));
  nor042aa1n02x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  nanp02aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  xnbna2aa1n03x5               g153(.a(new_n248), .b(new_n243), .c(new_n245), .out0(\s[23] ));
  nand22aa1n03x5               g154(.a(new_n243), .b(new_n245), .o1(new_n250));
  norp02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  nanb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(new_n253));
  aoai13aa1n02x5               g158(.a(new_n253), .b(new_n246), .c(new_n250), .d(new_n247), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n245), .o1(new_n255));
  aoai13aa1n02x5               g160(.a(new_n248), .b(new_n255), .c(new_n198), .d(new_n242), .o1(new_n256));
  nona22aa1n02x4               g161(.a(new_n256), .b(new_n253), .c(new_n246), .out0(new_n257));
  nanp02aa1n02x5               g162(.a(new_n254), .b(new_n257), .o1(\s[24] ));
  nano23aa1n06x5               g163(.a(new_n246), .b(new_n251), .c(new_n252), .d(new_n247), .out0(new_n259));
  nano22aa1n03x7               g164(.a(new_n223), .b(new_n241), .c(new_n259), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n204), .c(new_n127), .d(new_n189), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(new_n259), .b(new_n241), .o1(new_n262));
  inv040aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n02x5               g168(.a(new_n247), .b(new_n246), .c(new_n244), .d(new_n233), .o1(new_n264));
  oaoi03aa1n06x5               g169(.a(\a[24] ), .b(\b[23] ), .c(new_n264), .o1(new_n265));
  aoi012aa1n12x5               g170(.a(new_n265), .b(new_n225), .c(new_n263), .o1(new_n266));
  xorc02aa1n12x5               g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  xnbna2aa1n03x5               g172(.a(new_n267), .b(new_n261), .c(new_n266), .out0(\s[25] ));
  nand02aa1n03x5               g173(.a(new_n261), .b(new_n266), .o1(new_n269));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[25] ), .b(\a[26] ), .out0(new_n271));
  aoai13aa1n02x5               g176(.a(new_n271), .b(new_n270), .c(new_n269), .d(new_n267), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n266), .o1(new_n273));
  aoai13aa1n03x5               g178(.a(new_n267), .b(new_n273), .c(new_n198), .d(new_n260), .o1(new_n274));
  nona22aa1n02x4               g179(.a(new_n274), .b(new_n271), .c(new_n270), .out0(new_n275));
  nanp02aa1n02x5               g180(.a(new_n272), .b(new_n275), .o1(\s[26] ));
  norb02aa1n02x5               g181(.a(new_n267), .b(new_n271), .out0(new_n277));
  nano32aa1d12x5               g182(.a(new_n223), .b(new_n277), .c(new_n241), .d(new_n259), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n204), .c(new_n127), .d(new_n189), .o1(new_n279));
  orn002aa1n02x5               g184(.a(\a[20] ), .b(\b[19] ), .o(new_n280));
  and002aa1n02x5               g185(.a(\b[19] ), .b(\a[20] ), .o(new_n281));
  oaoi13aa1n06x5               g186(.a(new_n262), .b(new_n280), .c(new_n224), .d(new_n281), .o1(new_n282));
  inv000aa1d42x5               g187(.a(\a[26] ), .o1(new_n283));
  inv000aa1d42x5               g188(.a(\b[25] ), .o1(new_n284));
  oaoi03aa1n02x5               g189(.a(new_n283), .b(new_n284), .c(new_n270), .o1(new_n285));
  inv000aa1n02x5               g190(.a(new_n285), .o1(new_n286));
  oaoi13aa1n04x5               g191(.a(new_n286), .b(new_n277), .c(new_n282), .d(new_n265), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[27] ), .b(\b[26] ), .out0(new_n288));
  xnbna2aa1n03x5               g193(.a(new_n288), .b(new_n287), .c(new_n279), .out0(\s[27] ));
  nanp02aa1n06x5               g194(.a(new_n287), .b(new_n279), .o1(new_n290));
  norp02aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o1(new_n291));
  norp02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .o1(new_n292));
  nanp02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .o1(new_n293));
  nanb02aa1n02x5               g198(.a(new_n292), .b(new_n293), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n291), .c(new_n290), .d(new_n288), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n277), .b(new_n265), .c(new_n225), .d(new_n263), .o1(new_n296));
  nanp02aa1n03x5               g201(.a(new_n296), .b(new_n285), .o1(new_n297));
  aoai13aa1n02x5               g202(.a(new_n288), .b(new_n297), .c(new_n198), .d(new_n278), .o1(new_n298));
  nona22aa1n02x4               g203(.a(new_n298), .b(new_n294), .c(new_n291), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n295), .b(new_n299), .o1(\s[28] ));
  norb02aa1n03x5               g205(.a(new_n288), .b(new_n294), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n297), .c(new_n198), .d(new_n278), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n301), .o1(new_n303));
  oai012aa1n02x5               g208(.a(new_n293), .b(new_n292), .c(new_n291), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n303), .c(new_n287), .d(new_n279), .o1(new_n305));
  norp02aa1n02x5               g210(.a(\b[28] ), .b(\a[29] ), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(\b[28] ), .b(\a[29] ), .o1(new_n307));
  norb02aa1n02x5               g212(.a(new_n307), .b(new_n306), .out0(new_n308));
  oai022aa1n02x5               g213(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n309));
  aboi22aa1n03x5               g214(.a(new_n306), .b(new_n307), .c(new_n309), .d(new_n293), .out0(new_n310));
  aoi022aa1n03x5               g215(.a(new_n305), .b(new_n308), .c(new_n302), .d(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g216(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g217(.a(new_n294), .b(new_n288), .c(new_n308), .out0(new_n313));
  nanb02aa1n03x5               g218(.a(new_n313), .b(new_n290), .out0(new_n314));
  aoi013aa1n02x4               g219(.a(new_n306), .b(new_n309), .c(new_n293), .d(new_n307), .o1(new_n315));
  aoai13aa1n02x7               g220(.a(new_n315), .b(new_n313), .c(new_n287), .d(new_n279), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .out0(new_n317));
  aoi113aa1n02x5               g222(.a(new_n317), .b(new_n306), .c(new_n309), .d(new_n307), .e(new_n293), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n316), .d(new_n317), .o1(\s[30] ));
  nanp03aa1n02x5               g224(.a(new_n301), .b(new_n308), .c(new_n317), .o1(new_n320));
  nanb02aa1n03x5               g225(.a(new_n320), .b(new_n290), .out0(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  aoai13aa1n02x7               g229(.a(new_n323), .b(new_n320), .c(new_n287), .d(new_n279), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n321), .b(new_n324), .c(new_n325), .d(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g231(.a(new_n144), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi112aa1n02x5               g232(.a(new_n106), .b(new_n105), .c(new_n102), .d(new_n108), .o1(new_n328));
  aoib12aa1n02x5               g233(.a(new_n328), .b(new_n146), .c(new_n103), .out0(\s[4] ));
  norb02aa1n02x5               g234(.a(new_n119), .b(new_n118), .out0(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n330), .b(new_n109), .c(new_n110), .out0(\s[5] ));
  aoi012aa1n02x5               g236(.a(new_n118), .b(new_n146), .c(new_n119), .o1(new_n332));
  xnrb03aa1n02x5               g237(.a(new_n332), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g238(.a(new_n117), .b(new_n123), .c(new_n146), .d(new_n330), .o1(new_n334));
  xnrc02aa1n02x5               g239(.a(new_n334), .b(new_n122), .out0(\s[7] ));
  oaoi03aa1n02x5               g240(.a(\a[7] ), .b(\b[6] ), .c(new_n334), .o1(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g242(.a(new_n133), .b(new_n147), .c(new_n126), .out0(\s[9] ));
endmodule


