// Benchmark "adder" written by ABC on Thu Jul 18 01:06:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n337, new_n339,
    new_n341, new_n342, new_n343, new_n344, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor042aa1n06x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n06x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand42aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  tech160nm_fiaoi012aa1n04x5   g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  inv000aa1d42x5               g008(.a(\b[3] ), .o1(new_n104));
  nanb02aa1n02x5               g009(.a(\a[4] ), .b(new_n104), .out0(new_n105));
  nand02aa1n08x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(new_n105), .b(new_n106), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[3] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[2] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(new_n109), .b(new_n108), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(new_n110), .b(new_n111), .o1(new_n112));
  nor043aa1n02x5               g017(.a(new_n103), .b(new_n107), .c(new_n112), .o1(new_n113));
  nor042aa1n03x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nor042aa1n04x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  aoi012aa1n12x5               g020(.a(new_n114), .b(new_n115), .c(new_n106), .o1(new_n116));
  inv000aa1n02x5               g021(.a(new_n116), .o1(new_n117));
  nor002aa1d32x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nand22aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor002aa1d32x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nand22aa1n03x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nona23aa1n09x5               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  nor042aa1n06x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  nanp02aa1n24x5               g028(.a(\b[7] ), .b(\a[8] ), .o1(new_n124));
  nor042aa1n12x5               g029(.a(\b[6] ), .b(\a[7] ), .o1(new_n125));
  nanp02aa1n12x5               g030(.a(\b[6] ), .b(\a[7] ), .o1(new_n126));
  nona23aa1n02x4               g031(.a(new_n126), .b(new_n124), .c(new_n123), .d(new_n125), .out0(new_n127));
  nor002aa1n02x5               g032(.a(new_n127), .b(new_n122), .o1(new_n128));
  oai012aa1n06x5               g033(.a(new_n128), .b(new_n113), .c(new_n117), .o1(new_n129));
  nano23aa1d15x5               g034(.a(new_n123), .b(new_n125), .c(new_n126), .d(new_n124), .out0(new_n130));
  and002aa1n12x5               g035(.a(\b[5] ), .b(\a[6] ), .o(new_n131));
  oab012aa1d24x5               g036(.a(new_n131), .b(new_n118), .c(new_n120), .out0(new_n132));
  ao0012aa1n03x5               g037(.a(new_n123), .b(new_n125), .c(new_n124), .o(new_n133));
  aoi012aa1d18x5               g038(.a(new_n133), .b(new_n130), .c(new_n132), .o1(new_n134));
  xorc02aa1n12x5               g039(.a(\a[9] ), .b(\b[8] ), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  aoai13aa1n02x5               g041(.a(new_n99), .b(new_n136), .c(new_n129), .d(new_n134), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  inv000aa1n02x5               g043(.a(new_n100), .o1(new_n139));
  aob012aa1n03x5               g044(.a(new_n139), .b(new_n101), .c(new_n102), .out0(new_n140));
  norb02aa1n03x5               g045(.a(new_n106), .b(new_n114), .out0(new_n141));
  norb02aa1n06x5               g046(.a(new_n111), .b(new_n115), .out0(new_n142));
  nand23aa1n04x5               g047(.a(new_n140), .b(new_n141), .c(new_n142), .o1(new_n143));
  nano23aa1n06x5               g048(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n144));
  nand22aa1n03x5               g049(.a(new_n130), .b(new_n144), .o1(new_n145));
  aoai13aa1n12x5               g050(.a(new_n134), .b(new_n145), .c(new_n143), .d(new_n116), .o1(new_n146));
  tech160nm_fioaoi03aa1n03p5x5 g051(.a(new_n97), .b(new_n98), .c(new_n146), .o1(new_n147));
  oaoi03aa1n03x5               g052(.a(\a[10] ), .b(\b[9] ), .c(new_n147), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g054(.a(\b[10] ), .b(\a[11] ), .o1(new_n150));
  nand02aa1d04x5               g055(.a(\b[10] ), .b(\a[11] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  nor042aa1n04x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  nand02aa1d04x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(new_n155));
  aoai13aa1n02x5               g060(.a(new_n155), .b(new_n150), .c(new_n148), .d(new_n152), .o1(new_n156));
  nor042aa1n06x5               g061(.a(\b[9] ), .b(\a[10] ), .o1(new_n157));
  nand02aa1n04x5               g062(.a(\b[9] ), .b(\a[10] ), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n152), .b(new_n157), .c(new_n137), .d(new_n158), .o1(new_n159));
  nona22aa1n02x4               g064(.a(new_n159), .b(new_n155), .c(new_n150), .out0(new_n160));
  nanp02aa1n02x5               g065(.a(new_n156), .b(new_n160), .o1(\s[12] ));
  norb02aa1n06x4               g066(.a(new_n158), .b(new_n157), .out0(new_n162));
  nano23aa1n06x5               g067(.a(new_n150), .b(new_n153), .c(new_n154), .d(new_n151), .out0(new_n163));
  nand23aa1n02x5               g068(.a(new_n163), .b(new_n135), .c(new_n162), .o1(new_n164));
  aoai13aa1n12x5               g069(.a(new_n158), .b(new_n157), .c(new_n97), .d(new_n98), .o1(new_n165));
  inv000aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  tech160nm_fiaoi012aa1n02p5x5 g071(.a(new_n153), .b(new_n150), .c(new_n154), .o1(new_n167));
  aobi12aa1n03x5               g072(.a(new_n167), .b(new_n163), .c(new_n166), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n164), .c(new_n129), .d(new_n134), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nand02aa1n06x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  xnrb03aa1n03x5               g078(.a(new_n173), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nona23aa1n03x5               g079(.a(new_n154), .b(new_n151), .c(new_n150), .d(new_n153), .out0(new_n175));
  nano22aa1n02x5               g080(.a(new_n175), .b(new_n135), .c(new_n162), .out0(new_n176));
  oai012aa1n06x5               g081(.a(new_n167), .b(new_n175), .c(new_n165), .o1(new_n177));
  nor002aa1d32x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nand02aa1n06x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nona23aa1d18x5               g084(.a(new_n179), .b(new_n172), .c(new_n171), .d(new_n178), .out0(new_n180));
  inv000aa1n02x5               g085(.a(new_n180), .o1(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n177), .c(new_n146), .d(new_n176), .o1(new_n182));
  tech160nm_fioai012aa1n03p5x5 g087(.a(new_n179), .b(new_n178), .c(new_n171), .o1(new_n183));
  nor002aa1n06x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  nand42aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nanb02aa1n02x5               g090(.a(new_n184), .b(new_n185), .out0(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n182), .c(new_n183), .out0(\s[15] ));
  nand22aa1n03x5               g093(.a(new_n182), .b(new_n183), .o1(new_n189));
  nor002aa1n06x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nand02aa1n03x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nanb02aa1n02x5               g096(.a(new_n190), .b(new_n191), .out0(new_n192));
  aoai13aa1n02x5               g097(.a(new_n192), .b(new_n184), .c(new_n189), .d(new_n187), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(new_n189), .b(new_n187), .o1(new_n194));
  nona22aa1n02x4               g099(.a(new_n194), .b(new_n192), .c(new_n184), .out0(new_n195));
  nanp02aa1n02x5               g100(.a(new_n195), .b(new_n193), .o1(\s[16] ));
  nona23aa1n03x5               g101(.a(new_n191), .b(new_n185), .c(new_n184), .d(new_n190), .out0(new_n197));
  nor022aa1n04x5               g102(.a(new_n197), .b(new_n180), .o1(new_n198));
  nand02aa1n02x5               g103(.a(new_n176), .b(new_n198), .o1(new_n199));
  aoi012aa1n02x5               g104(.a(new_n190), .b(new_n184), .c(new_n191), .o1(new_n200));
  tech160nm_fioai012aa1n04x5   g105(.a(new_n200), .b(new_n197), .c(new_n183), .o1(new_n201));
  aoi012aa1n06x5               g106(.a(new_n201), .b(new_n177), .c(new_n198), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n129), .d(new_n134), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g109(.a(\a[17] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(\b[16] ), .b(new_n205), .out0(new_n206));
  nano23aa1n06x5               g111(.a(new_n184), .b(new_n190), .c(new_n191), .d(new_n185), .out0(new_n207));
  nano22aa1n12x5               g112(.a(new_n164), .b(new_n181), .c(new_n207), .out0(new_n208));
  nanb02aa1n12x5               g113(.a(new_n180), .b(new_n207), .out0(new_n209));
  oabi12aa1n09x5               g114(.a(new_n201), .b(new_n168), .c(new_n209), .out0(new_n210));
  xorc02aa1n02x5               g115(.a(\a[17] ), .b(\b[16] ), .out0(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n210), .c(new_n146), .d(new_n208), .o1(new_n212));
  xnrc02aa1n02x5               g117(.a(\b[17] ), .b(\a[18] ), .out0(new_n213));
  xobna2aa1n03x5               g118(.a(new_n213), .b(new_n212), .c(new_n206), .out0(\s[18] ));
  inv000aa1d42x5               g119(.a(\a[18] ), .o1(new_n215));
  xroi22aa1d04x5               g120(.a(new_n205), .b(\b[16] ), .c(new_n215), .d(\b[17] ), .out0(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n210), .c(new_n146), .d(new_n208), .o1(new_n217));
  oai022aa1n02x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  oaib12aa1n02x5               g123(.a(new_n218), .b(new_n215), .c(\b[17] ), .out0(new_n219));
  nor002aa1n06x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nand42aa1n02x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  nanb02aa1n02x5               g126(.a(new_n220), .b(new_n221), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n217), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand22aa1n02x5               g130(.a(new_n217), .b(new_n219), .o1(new_n226));
  nor002aa1n03x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nand02aa1n03x5               g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  nanb02aa1n02x5               g133(.a(new_n227), .b(new_n228), .out0(new_n229));
  aoai13aa1n02x5               g134(.a(new_n229), .b(new_n220), .c(new_n226), .d(new_n223), .o1(new_n230));
  oaoi03aa1n02x5               g135(.a(\a[18] ), .b(\b[17] ), .c(new_n206), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n223), .b(new_n231), .c(new_n203), .d(new_n216), .o1(new_n232));
  nona22aa1n02x4               g137(.a(new_n232), .b(new_n229), .c(new_n220), .out0(new_n233));
  nanp02aa1n02x5               g138(.a(new_n230), .b(new_n233), .o1(\s[20] ));
  nanp02aa1n06x5               g139(.a(new_n146), .b(new_n208), .o1(new_n235));
  nano23aa1n06x5               g140(.a(new_n220), .b(new_n227), .c(new_n228), .d(new_n221), .out0(new_n236));
  nanb03aa1n02x5               g141(.a(new_n213), .b(new_n236), .c(new_n211), .out0(new_n237));
  tech160nm_fiao0012aa1n02p5x5 g142(.a(new_n227), .b(new_n220), .c(new_n228), .o(new_n238));
  tech160nm_fiaoi012aa1n05x5   g143(.a(new_n238), .b(new_n236), .c(new_n231), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n237), .c(new_n235), .d(new_n202), .o1(new_n240));
  xorb03aa1n03x5               g145(.a(new_n240), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[20] ), .b(\a[21] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  tech160nm_fixnrc02aa1n04x5   g149(.a(\b[21] ), .b(\a[22] ), .out0(new_n245));
  aoai13aa1n02x7               g150(.a(new_n245), .b(new_n242), .c(new_n240), .d(new_n244), .o1(new_n246));
  nanp02aa1n04x5               g151(.a(new_n240), .b(new_n244), .o1(new_n247));
  nona22aa1n03x5               g152(.a(new_n247), .b(new_n245), .c(new_n242), .out0(new_n248));
  nanp02aa1n03x5               g153(.a(new_n248), .b(new_n246), .o1(\s[22] ));
  nor042aa1n03x5               g154(.a(new_n245), .b(new_n243), .o1(new_n250));
  nand23aa1n03x5               g155(.a(new_n216), .b(new_n250), .c(new_n236), .o1(new_n251));
  nona23aa1n09x5               g156(.a(new_n228), .b(new_n221), .c(new_n220), .d(new_n227), .out0(new_n252));
  oabi12aa1n06x5               g157(.a(new_n238), .b(new_n252), .c(new_n219), .out0(new_n253));
  inv000aa1d42x5               g158(.a(\a[22] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\b[21] ), .o1(new_n255));
  oao003aa1n03x5               g160(.a(new_n254), .b(new_n255), .c(new_n242), .carry(new_n256));
  aoi012aa1n02x5               g161(.a(new_n256), .b(new_n253), .c(new_n250), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n251), .c(new_n235), .d(new_n202), .o1(new_n258));
  xorb03aa1n02x5               g163(.a(new_n258), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(\b[22] ), .b(\a[23] ), .o1(new_n261));
  nanb02aa1n02x5               g166(.a(new_n260), .b(new_n261), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  nor042aa1n06x5               g168(.a(\b[23] ), .b(\a[24] ), .o1(new_n264));
  nand42aa1n03x5               g169(.a(\b[23] ), .b(\a[24] ), .o1(new_n265));
  nanb02aa1n02x5               g170(.a(new_n264), .b(new_n265), .out0(new_n266));
  aoai13aa1n02x7               g171(.a(new_n266), .b(new_n260), .c(new_n258), .d(new_n263), .o1(new_n267));
  nanp02aa1n04x5               g172(.a(new_n258), .b(new_n263), .o1(new_n268));
  nona22aa1n03x5               g173(.a(new_n268), .b(new_n266), .c(new_n260), .out0(new_n269));
  nanp02aa1n03x5               g174(.a(new_n269), .b(new_n267), .o1(\s[24] ));
  nona23aa1n09x5               g175(.a(new_n265), .b(new_n261), .c(new_n260), .d(new_n264), .out0(new_n271));
  inv020aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  nano22aa1n03x7               g177(.a(new_n237), .b(new_n250), .c(new_n272), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n210), .c(new_n146), .d(new_n208), .o1(new_n274));
  oai012aa1n02x5               g179(.a(new_n265), .b(new_n264), .c(new_n260), .o1(new_n275));
  oaib12aa1n02x5               g180(.a(new_n275), .b(new_n271), .c(new_n256), .out0(new_n276));
  nano22aa1n03x7               g181(.a(new_n239), .b(new_n250), .c(new_n272), .out0(new_n277));
  nona22aa1n03x5               g182(.a(new_n274), .b(new_n276), .c(new_n277), .out0(new_n278));
  xorb03aa1n02x5               g183(.a(new_n278), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n02x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[25] ), .b(\b[24] ), .out0(new_n281));
  tech160nm_fixnrc02aa1n05x5   g186(.a(\b[25] ), .b(\a[26] ), .out0(new_n282));
  aoai13aa1n02x5               g187(.a(new_n282), .b(new_n280), .c(new_n278), .d(new_n281), .o1(new_n283));
  aobi12aa1n03x7               g188(.a(new_n275), .b(new_n272), .c(new_n256), .out0(new_n284));
  nona32aa1n09x5               g189(.a(new_n253), .b(new_n271), .c(new_n245), .d(new_n243), .out0(new_n285));
  nanp02aa1n02x5               g190(.a(new_n285), .b(new_n284), .o1(new_n286));
  aoai13aa1n02x5               g191(.a(new_n281), .b(new_n286), .c(new_n203), .d(new_n273), .o1(new_n287));
  nona22aa1n02x4               g192(.a(new_n287), .b(new_n282), .c(new_n280), .out0(new_n288));
  nanp02aa1n02x5               g193(.a(new_n283), .b(new_n288), .o1(\s[26] ));
  norb02aa1n09x5               g194(.a(new_n281), .b(new_n282), .out0(new_n290));
  nano22aa1n03x7               g195(.a(new_n251), .b(new_n272), .c(new_n290), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n210), .c(new_n146), .d(new_n208), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\a[26] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[25] ), .o1(new_n294));
  tech160nm_fioaoi03aa1n02p5x5 g199(.a(new_n293), .b(new_n294), .c(new_n280), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  oaoi13aa1n12x5               g201(.a(new_n296), .b(new_n290), .c(new_n277), .d(new_n276), .o1(new_n297));
  xorc02aa1n02x5               g202(.a(\a[27] ), .b(\b[26] ), .out0(new_n298));
  xnbna2aa1n03x5               g203(.a(new_n298), .b(new_n297), .c(new_n292), .out0(\s[27] ));
  nanp02aa1n03x5               g204(.a(new_n297), .b(new_n292), .o1(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  tech160nm_fixorc02aa1n03p5x5 g206(.a(\a[28] ), .b(\b[27] ), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n301), .c(new_n300), .d(new_n298), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n290), .o1(new_n305));
  aoai13aa1n06x5               g210(.a(new_n295), .b(new_n305), .c(new_n285), .d(new_n284), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n298), .b(new_n306), .c(new_n203), .d(new_n291), .o1(new_n307));
  nona22aa1n02x4               g212(.a(new_n307), .b(new_n303), .c(new_n301), .out0(new_n308));
  nanp02aa1n03x5               g213(.a(new_n304), .b(new_n308), .o1(\s[28] ));
  and002aa1n02x5               g214(.a(new_n302), .b(new_n298), .o(new_n310));
  aoai13aa1n02x5               g215(.a(new_n310), .b(new_n306), .c(new_n203), .d(new_n291), .o1(new_n311));
  oai022aa1n02x5               g216(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n312));
  aob012aa1n02x5               g217(.a(new_n312), .b(\b[27] ), .c(\a[28] ), .out0(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .out0(new_n314));
  aoi012aa1n02x7               g219(.a(new_n314), .b(new_n311), .c(new_n313), .o1(new_n315));
  aobi12aa1n03x5               g220(.a(new_n310), .b(new_n297), .c(new_n292), .out0(new_n316));
  nano22aa1n03x7               g221(.a(new_n316), .b(new_n313), .c(new_n314), .out0(new_n317));
  nor002aa1n02x5               g222(.a(new_n315), .b(new_n317), .o1(\s[29] ));
  xorb03aa1n02x5               g223(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g224(.a(new_n314), .b(new_n298), .c(new_n302), .out0(new_n320));
  aoai13aa1n02x5               g225(.a(new_n320), .b(new_n306), .c(new_n203), .d(new_n291), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .carry(new_n322));
  xnrc02aa1n02x5               g227(.a(\b[29] ), .b(\a[30] ), .out0(new_n323));
  aoi012aa1n03x5               g228(.a(new_n323), .b(new_n321), .c(new_n322), .o1(new_n324));
  aobi12aa1n03x5               g229(.a(new_n320), .b(new_n297), .c(new_n292), .out0(new_n325));
  nano22aa1n03x7               g230(.a(new_n325), .b(new_n322), .c(new_n323), .out0(new_n326));
  nor002aa1n02x5               g231(.a(new_n324), .b(new_n326), .o1(\s[30] ));
  nano23aa1n02x4               g232(.a(new_n323), .b(new_n314), .c(new_n302), .d(new_n298), .out0(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n306), .c(new_n203), .d(new_n291), .o1(new_n329));
  oao003aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .c(new_n322), .carry(new_n330));
  xnrc02aa1n02x5               g235(.a(\b[30] ), .b(\a[31] ), .out0(new_n331));
  aoi012aa1n03x5               g236(.a(new_n331), .b(new_n329), .c(new_n330), .o1(new_n332));
  aobi12aa1n03x5               g237(.a(new_n328), .b(new_n297), .c(new_n292), .out0(new_n333));
  nano22aa1n03x7               g238(.a(new_n333), .b(new_n330), .c(new_n331), .out0(new_n334));
  nor002aa1n02x5               g239(.a(new_n332), .b(new_n334), .o1(\s[31] ));
  xnbna2aa1n03x5               g240(.a(new_n103), .b(new_n111), .c(new_n110), .out0(\s[3] ));
  aoi112aa1n02x5               g241(.a(new_n115), .b(new_n141), .c(new_n140), .d(new_n142), .o1(new_n337));
  oaoi13aa1n02x5               g242(.a(new_n337), .b(new_n105), .c(new_n113), .d(new_n117), .o1(\s[4] ));
  nanb02aa1n02x5               g243(.a(new_n120), .b(new_n121), .out0(new_n339));
  xobna2aa1n03x5               g244(.a(new_n339), .b(new_n143), .c(new_n116), .out0(\s[5] ));
  oabi12aa1n02x5               g245(.a(new_n339), .b(new_n113), .c(new_n117), .out0(new_n341));
  aoib12aa1n02x5               g246(.a(new_n120), .b(new_n119), .c(new_n118), .out0(new_n342));
  inv000aa1d42x5               g247(.a(new_n132), .o1(new_n343));
  aoai13aa1n02x5               g248(.a(new_n343), .b(new_n122), .c(new_n143), .d(new_n116), .o1(new_n344));
  aboi22aa1n03x5               g249(.a(new_n118), .b(new_n344), .c(new_n341), .d(new_n342), .out0(\s[6] ));
  xorb03aa1n02x5               g250(.a(new_n344), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g251(.a(new_n125), .b(new_n344), .c(new_n126), .o1(new_n347));
  xnrb03aa1n02x5               g252(.a(new_n347), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g253(.a(new_n146), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


