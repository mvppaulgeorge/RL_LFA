// Benchmark "adder" written by ABC on Thu Jul 18 04:41:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n348, new_n349, new_n351, new_n352, new_n354,
    new_n355, new_n357, new_n358, new_n359, new_n360, new_n362, new_n363,
    new_n365;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n12x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  orn002aa1n24x5               g002(.a(\a[2] ), .b(\b[1] ), .o(new_n98));
  nanp02aa1n06x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  aob012aa1n12x5               g004(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(new_n100));
  inv040aa1d32x5               g005(.a(\a[3] ), .o1(new_n101));
  inv030aa1d28x5               g006(.a(\b[2] ), .o1(new_n102));
  nand02aa1d06x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand02aa1d04x5               g009(.a(new_n103), .b(new_n104), .o1(new_n105));
  aoi012aa1n03x5               g010(.a(new_n105), .b(new_n100), .c(new_n98), .o1(new_n106));
  oai022aa1n02x5               g011(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n107));
  norp02aa1n03x5               g012(.a(new_n106), .b(new_n107), .o1(new_n108));
  nand02aa1d28x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand42aa1n16x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  oai112aa1n06x5               g015(.a(new_n109), .b(new_n110), .c(\b[5] ), .d(\a[6] ), .o1(new_n111));
  aoi022aa1d24x5               g016(.a(\b[5] ), .b(\a[6] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n112));
  oai022aa1n03x5               g017(.a(\a[5] ), .b(\b[4] ), .c(\b[6] ), .d(\a[7] ), .o1(new_n113));
  nor042aa1d18x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  aoi012aa1n12x5               g019(.a(new_n114), .b(\a[7] ), .c(\b[6] ), .o1(new_n115));
  nona23aa1n03x5               g020(.a(new_n115), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n116));
  nand42aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1n06x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  inv030aa1n02x5               g023(.a(new_n118), .o1(new_n119));
  nand02aa1n03x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nanb03aa1n03x5               g025(.a(new_n114), .b(new_n109), .c(new_n120), .out0(new_n121));
  oaih22aa1d12x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  nano32aa1n03x7               g027(.a(new_n121), .b(new_n122), .c(new_n119), .d(new_n117), .out0(new_n123));
  tech160nm_fiaoi012aa1n02p5x5 g028(.a(new_n114), .b(new_n118), .c(new_n109), .o1(new_n124));
  norb02aa1n09x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  tech160nm_fioai012aa1n05x5   g030(.a(new_n125), .b(new_n108), .c(new_n116), .o1(new_n126));
  nanp02aa1n06x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  aoi012aa1n02x5               g032(.a(new_n97), .b(new_n126), .c(new_n127), .o1(new_n128));
  nor022aa1n12x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1d12x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  norb02aa1n02x5               g036(.a(new_n127), .b(new_n97), .out0(new_n132));
  oai022aa1d24x5               g037(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  aoi122aa1n02x5               g038(.a(new_n133), .b(\b[9] ), .c(\a[10] ), .d(new_n126), .e(new_n132), .o1(new_n134));
  oabi12aa1n02x5               g039(.a(new_n134), .b(new_n128), .c(new_n131), .out0(\s[10] ));
  oai012aa1n02x5               g040(.a(new_n130), .b(new_n129), .c(new_n97), .o1(new_n136));
  nano23aa1n02x4               g041(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n127), .out0(new_n137));
  nanp02aa1n03x5               g042(.a(new_n126), .b(new_n137), .o1(new_n138));
  xnrc02aa1n12x5               g043(.a(\b[10] ), .b(\a[11] ), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n138), .c(new_n136), .out0(\s[11] ));
  nor042aa1d18x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand22aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  inv000aa1d42x5               g049(.a(\a[11] ), .o1(new_n145));
  aob012aa1n03x5               g050(.a(new_n140), .b(new_n138), .c(new_n136), .out0(new_n146));
  oaib12aa1n06x5               g051(.a(new_n146), .b(\b[10] ), .c(new_n145), .out0(new_n147));
  norp02aa1n04x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nona23aa1n02x4               g053(.a(new_n146), .b(new_n143), .c(new_n142), .d(new_n148), .out0(new_n149));
  aob012aa1n03x5               g054(.a(new_n149), .b(new_n147), .c(new_n144), .out0(\s[12] ));
  nona22aa1n02x4               g055(.a(new_n137), .b(new_n139), .c(new_n144), .out0(new_n151));
  inv000aa1n02x5               g056(.a(new_n151), .o1(new_n152));
  nand22aa1n03x5               g057(.a(new_n126), .b(new_n152), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(\b[10] ), .b(\a[11] ), .o1(new_n154));
  nanb03aa1n06x5               g059(.a(new_n142), .b(new_n143), .c(new_n154), .out0(new_n155));
  oai112aa1n06x5               g060(.a(new_n133), .b(new_n130), .c(\b[10] ), .d(\a[11] ), .o1(new_n156));
  tech160nm_fiaoi012aa1n03p5x5 g061(.a(new_n142), .b(new_n148), .c(new_n143), .o1(new_n157));
  tech160nm_fioai012aa1n05x5   g062(.a(new_n157), .b(new_n156), .c(new_n155), .o1(new_n158));
  nanb02aa1n06x5               g063(.a(new_n158), .b(new_n153), .out0(new_n159));
  nor002aa1d32x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand22aa1n09x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nanb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  oai112aa1n02x5               g068(.a(new_n157), .b(new_n162), .c(new_n156), .d(new_n155), .o1(new_n164));
  aboi22aa1n03x5               g069(.a(new_n164), .b(new_n153), .c(new_n159), .d(new_n163), .out0(\s[13] ));
  inv000aa1d42x5               g070(.a(new_n160), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n163), .b(new_n158), .c(new_n126), .d(new_n152), .o1(new_n167));
  nor002aa1n12x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand22aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  oai022aa1d24x5               g075(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n171));
  nanb03aa1n02x5               g076(.a(new_n171), .b(new_n167), .c(new_n169), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n170), .c(new_n166), .d(new_n167), .o1(\s[14] ));
  nano23aa1n06x5               g078(.a(new_n160), .b(new_n168), .c(new_n169), .d(new_n161), .out0(new_n174));
  oaoi03aa1n02x5               g079(.a(\a[14] ), .b(\b[13] ), .c(new_n166), .o1(new_n175));
  nor002aa1d32x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nand22aa1n04x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanb02aa1n06x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  inv040aa1d30x5               g083(.a(new_n178), .o1(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n175), .c(new_n159), .d(new_n174), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n175), .c(new_n159), .d(new_n174), .o1(new_n181));
  norb02aa1n03x4               g086(.a(new_n180), .b(new_n181), .out0(\s[15] ));
  inv000aa1d42x5               g087(.a(new_n176), .o1(new_n183));
  nor002aa1d32x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand02aa1n06x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  norb03aa1n02x5               g091(.a(new_n185), .b(new_n176), .c(new_n184), .out0(new_n187));
  nanp02aa1n03x5               g092(.a(new_n180), .b(new_n187), .o1(new_n188));
  aoai13aa1n03x5               g093(.a(new_n188), .b(new_n186), .c(new_n183), .d(new_n180), .o1(\s[16] ));
  nano32aa1n03x7               g094(.a(new_n151), .b(new_n186), .c(new_n174), .d(new_n179), .out0(new_n190));
  nanp02aa1n04x5               g095(.a(new_n126), .b(new_n190), .o1(new_n191));
  oa0022aa1n09x5               g096(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n105), .c(new_n100), .d(new_n98), .o1(new_n193));
  nano23aa1n02x5               g098(.a(new_n111), .b(new_n113), .c(new_n115), .d(new_n112), .out0(new_n194));
  nanp02aa1n06x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  nona23aa1n02x4               g100(.a(new_n130), .b(new_n127), .c(new_n97), .d(new_n129), .out0(new_n196));
  nona23aa1n09x5               g101(.a(new_n169), .b(new_n161), .c(new_n160), .d(new_n168), .out0(new_n197));
  nona23aa1n12x5               g102(.a(new_n185), .b(new_n177), .c(new_n176), .d(new_n184), .out0(new_n198));
  nor042aa1n06x5               g103(.a(new_n198), .b(new_n197), .o1(new_n199));
  nona32aa1n09x5               g104(.a(new_n199), .b(new_n196), .c(new_n144), .d(new_n139), .out0(new_n200));
  aoi022aa1d24x5               g105(.a(\b[14] ), .b(\a[15] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n201));
  tech160nm_fiaoi012aa1n03p5x5 g106(.a(new_n176), .b(new_n171), .c(new_n201), .o1(new_n202));
  oaoi03aa1n03x5               g107(.a(\a[16] ), .b(\b[15] ), .c(new_n202), .o1(new_n203));
  aoi012aa1n09x5               g108(.a(new_n203), .b(new_n158), .c(new_n199), .o1(new_n204));
  aoai13aa1n12x5               g109(.a(new_n204), .b(new_n200), .c(new_n195), .d(new_n125), .o1(new_n205));
  tech160nm_fixorc02aa1n02p5x5 g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  norb02aa1n02x5               g111(.a(new_n185), .b(new_n202), .out0(new_n207));
  oabi12aa1n02x5               g112(.a(new_n206), .b(\a[16] ), .c(\b[15] ), .out0(new_n208));
  aoi112aa1n02x5               g113(.a(new_n208), .b(new_n207), .c(new_n158), .d(new_n199), .o1(new_n209));
  aoi022aa1n02x5               g114(.a(new_n205), .b(new_n206), .c(new_n191), .d(new_n209), .o1(\s[17] ));
  nor042aa1n03x5               g115(.a(\b[16] ), .b(\a[17] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  inv000aa1d42x5               g117(.a(\a[17] ), .o1(new_n213));
  oaib12aa1n06x5               g118(.a(new_n205), .b(new_n213), .c(\b[16] ), .out0(new_n214));
  tech160nm_fixorc02aa1n02p5x5 g119(.a(\a[18] ), .b(\b[17] ), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n214), .c(new_n212), .out0(\s[18] ));
  inv000aa1d42x5               g121(.a(\a[18] ), .o1(new_n217));
  xroi22aa1d04x5               g122(.a(new_n213), .b(\b[16] ), .c(new_n217), .d(\b[17] ), .out0(new_n218));
  nand02aa1d06x5               g123(.a(new_n205), .b(new_n218), .o1(new_n219));
  oao003aa1n03x5               g124(.a(\a[18] ), .b(\b[17] ), .c(new_n212), .carry(new_n220));
  xorc02aa1n12x5               g125(.a(\a[19] ), .b(\b[18] ), .out0(new_n221));
  xnbna2aa1n03x5               g126(.a(new_n221), .b(new_n219), .c(new_n220), .out0(\s[19] ));
  xnrc02aa1n02x5               g127(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  xnrc02aa1n02x5               g128(.a(\b[19] ), .b(\a[20] ), .out0(new_n224));
  nor042aa1n09x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  inv030aa1n02x5               g130(.a(new_n225), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n221), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n226), .b(new_n227), .c(new_n219), .d(new_n220), .o1(new_n228));
  norp02aa1n04x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  and002aa1n03x5               g134(.a(\b[19] ), .b(\a[20] ), .o(new_n230));
  norp03aa1n02x5               g135(.a(new_n230), .b(new_n229), .c(new_n225), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n231), .b(new_n227), .c(new_n219), .d(new_n220), .o1(new_n232));
  aob012aa1n03x5               g137(.a(new_n232), .b(new_n228), .c(new_n224), .out0(\s[20] ));
  nano32aa1n03x7               g138(.a(new_n224), .b(new_n221), .c(new_n215), .d(new_n206), .out0(new_n234));
  oaih22aa1n04x5               g139(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n235));
  aoi112aa1n03x5               g140(.a(new_n230), .b(new_n229), .c(\a[19] ), .d(\b[18] ), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n225), .b(\a[18] ), .c(\b[17] ), .o1(new_n237));
  nand23aa1n03x5               g142(.a(new_n236), .b(new_n235), .c(new_n237), .o1(new_n238));
  oab012aa1n04x5               g143(.a(new_n229), .b(new_n226), .c(new_n230), .out0(new_n239));
  nanp02aa1n02x5               g144(.a(new_n238), .b(new_n239), .o1(new_n240));
  xorc02aa1n12x5               g145(.a(\a[21] ), .b(\b[20] ), .out0(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n240), .c(new_n205), .d(new_n234), .o1(new_n242));
  nano22aa1n02x4               g147(.a(new_n241), .b(new_n238), .c(new_n239), .out0(new_n243));
  aobi12aa1n02x5               g148(.a(new_n243), .b(new_n205), .c(new_n234), .out0(new_n244));
  norb02aa1n03x4               g149(.a(new_n242), .b(new_n244), .out0(\s[21] ));
  nor042aa1n04x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[22] ), .b(\b[21] ), .out0(new_n248));
  inv000aa1d42x5               g153(.a(\a[22] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\b[21] ), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n246), .b(new_n249), .c(new_n250), .o1(new_n251));
  oai112aa1n03x5               g156(.a(new_n242), .b(new_n251), .c(new_n250), .d(new_n249), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n248), .c(new_n242), .d(new_n247), .o1(\s[22] ));
  nand02aa1d06x5               g158(.a(new_n248), .b(new_n241), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  nano32aa1n02x4               g160(.a(new_n224), .b(new_n255), .c(new_n218), .d(new_n221), .out0(new_n256));
  tech160nm_fioaoi03aa1n03p5x5 g161(.a(new_n249), .b(new_n250), .c(new_n246), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n254), .c(new_n238), .d(new_n239), .o1(new_n258));
  tech160nm_fixorc02aa1n04x5   g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n258), .c(new_n205), .d(new_n256), .o1(new_n260));
  nanb02aa1n02x5               g165(.a(new_n259), .b(new_n257), .out0(new_n261));
  aoi122aa1n02x7               g166(.a(new_n261), .b(new_n240), .c(new_n255), .d(new_n205), .e(new_n256), .o1(new_n262));
  norb02aa1n03x4               g167(.a(new_n260), .b(new_n262), .out0(\s[23] ));
  nor042aa1n06x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  nor002aa1n02x5               g170(.a(\b[23] ), .b(\a[24] ), .o1(new_n266));
  nand42aa1n10x5               g171(.a(\b[23] ), .b(\a[24] ), .o1(new_n267));
  norb02aa1n02x5               g172(.a(new_n267), .b(new_n266), .out0(new_n268));
  nona23aa1n03x5               g173(.a(new_n260), .b(new_n267), .c(new_n266), .d(new_n264), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n268), .c(new_n265), .d(new_n260), .o1(\s[24] ));
  inv000aa1n02x5               g175(.a(new_n234), .o1(new_n271));
  nano22aa1n03x7               g176(.a(new_n254), .b(new_n259), .c(new_n268), .out0(new_n272));
  norb02aa1n02x5               g177(.a(new_n272), .b(new_n271), .out0(new_n273));
  and002aa1n02x5               g178(.a(new_n259), .b(new_n268), .o(new_n274));
  nanp02aa1n02x5               g179(.a(new_n258), .b(new_n274), .o1(new_n275));
  aoi012aa1n02x5               g180(.a(new_n266), .b(new_n264), .c(new_n267), .o1(new_n276));
  nand02aa1n02x5               g181(.a(new_n275), .b(new_n276), .o1(new_n277));
  tech160nm_fixorc02aa1n03p5x5 g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n205), .d(new_n273), .o1(new_n279));
  inv000aa1n02x5               g184(.a(new_n276), .o1(new_n280));
  nona22aa1n02x4               g185(.a(new_n275), .b(new_n280), .c(new_n278), .out0(new_n281));
  aoi012aa1n02x5               g186(.a(new_n281), .b(new_n205), .c(new_n273), .o1(new_n282));
  norb02aa1n03x4               g187(.a(new_n279), .b(new_n282), .out0(\s[25] ));
  norp02aa1n02x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .out0(new_n286));
  and002aa1n02x5               g191(.a(\b[25] ), .b(\a[26] ), .o(new_n287));
  oai022aa1n02x5               g192(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n288));
  nona22aa1n03x5               g193(.a(new_n279), .b(new_n287), .c(new_n288), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n286), .c(new_n285), .d(new_n279), .o1(\s[26] ));
  and002aa1n02x5               g195(.a(new_n286), .b(new_n278), .o(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n280), .c(new_n258), .d(new_n274), .o1(new_n292));
  inv040aa1n03x5               g197(.a(new_n292), .o1(new_n293));
  nand03aa1n02x5               g198(.a(new_n234), .b(new_n272), .c(new_n291), .o1(new_n294));
  aob012aa1n02x5               g199(.a(new_n288), .b(\b[25] ), .c(\a[26] ), .out0(new_n295));
  aoai13aa1n04x5               g200(.a(new_n295), .b(new_n294), .c(new_n191), .d(new_n204), .o1(new_n296));
  norp02aa1n02x5               g201(.a(\b[26] ), .b(\a[27] ), .o1(new_n297));
  and002aa1n24x5               g202(.a(\b[26] ), .b(\a[27] ), .o(new_n298));
  norp02aa1n02x5               g203(.a(new_n298), .b(new_n297), .o1(new_n299));
  nano22aa1n03x7               g204(.a(new_n271), .b(new_n272), .c(new_n291), .out0(new_n300));
  inv000aa1n06x5               g205(.a(new_n297), .o1(new_n301));
  oaib12aa1n02x5               g206(.a(new_n295), .b(new_n298), .c(new_n301), .out0(new_n302));
  aoi112aa1n02x7               g207(.a(new_n293), .b(new_n302), .c(new_n205), .d(new_n300), .o1(new_n303));
  oaoi13aa1n02x7               g208(.a(new_n303), .b(new_n299), .c(new_n293), .d(new_n296), .o1(\s[27] ));
  inv000aa1d42x5               g209(.a(new_n298), .o1(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(new_n296), .c(new_n293), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n287), .o1(new_n307));
  aoi022aa1n09x5               g212(.a(new_n205), .b(new_n300), .c(new_n307), .d(new_n288), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n301), .b(new_n298), .c(new_n308), .d(new_n292), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[28] ), .b(\b[27] ), .out0(new_n310));
  norp02aa1n02x5               g215(.a(new_n310), .b(new_n297), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n306), .d(new_n311), .o1(\s[28] ));
  inv000aa1d42x5               g217(.a(\a[27] ), .o1(new_n313));
  inv000aa1d42x5               g218(.a(\a[28] ), .o1(new_n314));
  xroi22aa1d06x4               g219(.a(new_n313), .b(\b[26] ), .c(new_n314), .d(\b[27] ), .out0(new_n315));
  oai012aa1n02x5               g220(.a(new_n315), .b(new_n296), .c(new_n293), .o1(new_n316));
  inv000aa1n06x5               g221(.a(new_n315), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[28] ), .b(\b[27] ), .c(new_n301), .carry(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n308), .d(new_n292), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .out0(new_n320));
  norb02aa1n02x5               g225(.a(new_n318), .b(new_n320), .out0(new_n321));
  aoi022aa1n03x5               g226(.a(new_n319), .b(new_n320), .c(new_n316), .d(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g228(.a(new_n310), .b(new_n320), .c(new_n299), .o(new_n324));
  oai012aa1n02x5               g229(.a(new_n324), .b(new_n296), .c(new_n293), .o1(new_n325));
  inv000aa1n02x5               g230(.a(new_n324), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\b[28] ), .o1(new_n327));
  inv000aa1d42x5               g232(.a(\a[29] ), .o1(new_n328));
  oaib12aa1n02x5               g233(.a(new_n318), .b(\b[28] ), .c(new_n328), .out0(new_n329));
  oaib12aa1n02x5               g234(.a(new_n329), .b(new_n327), .c(\a[29] ), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n326), .c(new_n308), .d(new_n292), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .out0(new_n332));
  oaoi13aa1n02x5               g237(.a(new_n332), .b(new_n329), .c(new_n328), .d(new_n327), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n331), .b(new_n332), .c(new_n325), .d(new_n333), .o1(\s[30] ));
  nano22aa1n02x4               g239(.a(new_n317), .b(new_n320), .c(new_n332), .out0(new_n335));
  oai012aa1n02x5               g240(.a(new_n335), .b(new_n296), .c(new_n293), .o1(new_n336));
  aoi022aa1n02x5               g241(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n337));
  norb02aa1n02x5               g242(.a(\b[30] ), .b(\a[31] ), .out0(new_n338));
  obai22aa1n02x7               g243(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n339));
  aoi112aa1n02x5               g244(.a(new_n339), .b(new_n338), .c(new_n329), .d(new_n337), .o1(new_n340));
  xorc02aa1n02x5               g245(.a(\a[31] ), .b(\b[30] ), .out0(new_n341));
  inv000aa1n02x5               g246(.a(new_n335), .o1(new_n342));
  norp02aa1n02x5               g247(.a(\b[29] ), .b(\a[30] ), .o1(new_n343));
  aoi012aa1n02x5               g248(.a(new_n343), .b(new_n329), .c(new_n337), .o1(new_n344));
  aoai13aa1n03x5               g249(.a(new_n344), .b(new_n342), .c(new_n308), .d(new_n292), .o1(new_n345));
  aoi022aa1n03x5               g250(.a(new_n345), .b(new_n341), .c(new_n336), .d(new_n340), .o1(\s[31] ));
  xobna2aa1n03x5               g251(.a(new_n105), .b(new_n100), .c(new_n98), .out0(\s[3] ));
  xorc02aa1n02x5               g252(.a(\a[4] ), .b(\b[3] ), .out0(new_n348));
  norb02aa1n02x5               g253(.a(new_n103), .b(new_n348), .out0(new_n349));
  aboi22aa1n03x5               g254(.a(new_n106), .b(new_n349), .c(new_n193), .d(new_n348), .out0(\s[4] ));
  nanp02aa1n02x5               g255(.a(\b[3] ), .b(\a[4] ), .o1(new_n351));
  xorc02aa1n02x5               g256(.a(\a[5] ), .b(\b[4] ), .out0(new_n352));
  xobna2aa1n03x5               g257(.a(new_n352), .b(new_n193), .c(new_n351), .out0(\s[5] ));
  aob012aa1n03x5               g258(.a(new_n352), .b(new_n193), .c(new_n351), .out0(new_n354));
  xorc02aa1n02x5               g259(.a(\a[6] ), .b(\b[5] ), .out0(new_n355));
  xobna2aa1n03x5               g260(.a(new_n355), .b(new_n354), .c(new_n110), .out0(\s[6] ));
  aobi12aa1n02x5               g261(.a(new_n355), .b(new_n354), .c(new_n110), .out0(new_n357));
  aboi22aa1n03x5               g262(.a(new_n357), .b(new_n117), .c(new_n119), .d(new_n120), .out0(new_n358));
  nano22aa1n02x4               g263(.a(new_n118), .b(new_n117), .c(new_n120), .out0(new_n359));
  nanb02aa1n06x5               g264(.a(new_n357), .b(new_n359), .out0(new_n360));
  norb02aa1n02x5               g265(.a(new_n360), .b(new_n358), .out0(\s[7] ));
  norb02aa1n02x5               g266(.a(new_n109), .b(new_n114), .out0(new_n362));
  nona23aa1n02x4               g267(.a(new_n360), .b(new_n109), .c(new_n118), .d(new_n114), .out0(new_n363));
  aoai13aa1n02x5               g268(.a(new_n363), .b(new_n362), .c(new_n119), .d(new_n360), .o1(\s[8] ));
  norb03aa1n02x5               g269(.a(new_n124), .b(new_n123), .c(new_n132), .out0(new_n365));
  aoi022aa1n02x5               g270(.a(new_n126), .b(new_n132), .c(new_n195), .d(new_n365), .o1(\s[9] ));
endmodule


