// Benchmark "adder" written by ABC on Wed Jul 17 21:02:57 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n323, new_n324, new_n325,
    new_n327, new_n328, new_n330, new_n331, new_n332, new_n333, new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  tech160nm_fixnrc02aa1n04x5   g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norp02aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai012aa1n04x7               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  tech160nm_fixnrc02aa1n05x5   g009(.a(\b[3] ), .b(\a[4] ), .out0(new_n105));
  nor042aa1n02x5               g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n103), .c(new_n99), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nor042aa1n06x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand42aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  norb02aa1n03x5               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  aoi022aa1d24x5               g016(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n112));
  norp02aa1n12x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  aoi012aa1n02x7               g018(.a(new_n113), .b(\a[4] ), .c(\b[3] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  norp02aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nona22aa1n02x4               g021(.a(new_n114), .b(new_n115), .c(new_n116), .out0(new_n117));
  nano32aa1n03x7               g022(.a(new_n117), .b(new_n111), .c(new_n112), .d(new_n108), .out0(new_n118));
  oai012aa1n02x7               g023(.a(new_n110), .b(new_n115), .c(new_n109), .o1(new_n119));
  nona23aa1n06x5               g024(.a(new_n112), .b(new_n110), .c(new_n115), .d(new_n109), .out0(new_n120));
  and002aa1n12x5               g025(.a(\b[5] ), .b(\a[6] ), .o(new_n121));
  nor043aa1n06x5               g026(.a(new_n121), .b(new_n113), .c(new_n116), .o1(new_n122));
  oai012aa1n12x5               g027(.a(new_n119), .b(new_n120), .c(new_n122), .o1(new_n123));
  nand42aa1n16x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n97), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n123), .c(new_n107), .d(new_n118), .o1(new_n126));
  nor042aa1n04x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n20x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  oai022aa1d18x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  nanb03aa1n02x5               g035(.a(new_n130), .b(new_n126), .c(new_n128), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n129), .c(new_n98), .d(new_n126), .o1(\s[10] ));
  nano23aa1d18x5               g037(.a(new_n97), .b(new_n127), .c(new_n128), .d(new_n124), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n123), .c(new_n107), .d(new_n118), .o1(new_n134));
  oai012aa1n02x5               g039(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n135));
  nor002aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand02aa1n06x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n134), .c(new_n135), .out0(\s[11] ));
  aobi12aa1n02x5               g044(.a(new_n138), .b(new_n134), .c(new_n135), .out0(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  nor042aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n143), .b(new_n141), .out0(new_n144));
  oai012aa1n02x5               g049(.a(new_n144), .b(new_n140), .c(new_n136), .o1(new_n145));
  oai022aa1d18x5               g050(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n146));
  oai013aa1n02x4               g051(.a(new_n145), .b(new_n142), .c(new_n140), .d(new_n146), .o1(\s[12] ));
  nano23aa1n09x5               g052(.a(new_n136), .b(new_n143), .c(new_n141), .d(new_n137), .out0(new_n148));
  nand22aa1n12x5               g053(.a(new_n148), .b(new_n133), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n123), .c(new_n107), .d(new_n118), .o1(new_n151));
  aoi022aa1d24x5               g056(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n152));
  aoai13aa1n12x5               g057(.a(new_n141), .b(new_n146), .c(new_n130), .d(new_n152), .o1(new_n153));
  nor002aa1d32x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nanp02aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n151), .c(new_n153), .out0(\s[13] ));
  inv000aa1d42x5               g062(.a(new_n154), .o1(new_n158));
  aob012aa1n02x5               g063(.a(new_n156), .b(new_n151), .c(new_n153), .out0(new_n159));
  nor002aa1n20x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n04x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  nona23aa1n02x4               g067(.a(new_n159), .b(new_n161), .c(new_n160), .d(new_n154), .out0(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n162), .c(new_n158), .d(new_n159), .o1(\s[14] ));
  nona23aa1n12x5               g069(.a(new_n161), .b(new_n155), .c(new_n154), .d(new_n160), .out0(new_n165));
  oai012aa1n12x5               g070(.a(new_n161), .b(new_n160), .c(new_n154), .o1(new_n166));
  oai012aa1d24x5               g071(.a(new_n166), .b(new_n153), .c(new_n165), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  tech160nm_fioai012aa1n05x5   g073(.a(new_n168), .b(new_n151), .c(new_n165), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand02aa1n06x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  nor042aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n12x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  norb02aa1n02x5               g081(.a(new_n172), .b(new_n171), .out0(new_n177));
  oai022aa1n02x5               g082(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n178));
  aoi122aa1n02x5               g083(.a(new_n178), .b(\b[15] ), .c(\a[16] ), .d(new_n169), .e(new_n177), .o1(new_n179));
  oabi12aa1n02x7               g084(.a(new_n179), .b(new_n173), .c(new_n176), .out0(\s[16] ));
  nano23aa1n03x7               g085(.a(new_n154), .b(new_n160), .c(new_n161), .d(new_n155), .out0(new_n181));
  nano23aa1d15x5               g086(.a(new_n171), .b(new_n174), .c(new_n175), .d(new_n172), .out0(new_n182));
  nano22aa1n12x5               g087(.a(new_n149), .b(new_n181), .c(new_n182), .out0(new_n183));
  aoai13aa1n12x5               g088(.a(new_n183), .b(new_n123), .c(new_n107), .d(new_n118), .o1(new_n184));
  aoi022aa1d18x5               g089(.a(new_n167), .b(new_n182), .c(new_n175), .d(new_n178), .o1(new_n185));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n184), .out0(\s[17] ));
  nor042aa1n06x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  nand42aa1n10x5               g094(.a(new_n185), .b(new_n184), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n190), .b(new_n186), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[18] ), .b(\b[17] ), .out0(new_n192));
  nanp02aa1n04x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  oai022aa1d18x5               g098(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n194));
  nanb03aa1n03x5               g099(.a(new_n194), .b(new_n191), .c(new_n193), .out0(new_n195));
  aoai13aa1n02x5               g100(.a(new_n195), .b(new_n192), .c(new_n189), .d(new_n191), .o1(\s[18] ));
  nanp02aa1n02x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  norp02aa1n02x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nano23aa1n06x5               g103(.a(new_n188), .b(new_n198), .c(new_n193), .d(new_n197), .out0(new_n199));
  oaoi03aa1n02x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n200));
  tech160nm_fixorc02aa1n03p5x5 g105(.a(\a[19] ), .b(\b[18] ), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n202));
  aoi112aa1n02x5               g107(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n203));
  norb02aa1n03x4               g108(.a(new_n202), .b(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[18] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  xorc02aa1n02x5               g113(.a(\a[20] ), .b(\b[19] ), .out0(new_n209));
  nanp02aa1n02x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  oai022aa1n02x5               g115(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n211));
  norb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  tech160nm_finand02aa1n05x5   g117(.a(new_n202), .b(new_n212), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n208), .d(new_n202), .o1(\s[20] ));
  and003aa1n06x5               g119(.a(new_n199), .b(new_n209), .c(new_n201), .o(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  oai112aa1n02x5               g121(.a(new_n194), .b(new_n193), .c(new_n207), .d(new_n206), .o1(new_n217));
  aboi22aa1n03x5               g122(.a(new_n211), .b(new_n217), .c(\a[20] ), .d(\b[19] ), .out0(new_n218));
  inv000aa1n02x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n04x5               g124(.a(new_n219), .b(new_n216), .c(new_n185), .d(new_n184), .o1(new_n220));
  nor042aa1n03x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  nanp02aa1n04x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1n06x4               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  aoi112aa1n02x5               g128(.a(new_n223), .b(new_n218), .c(new_n190), .d(new_n215), .o1(new_n224));
  aoi012aa1n02x5               g129(.a(new_n224), .b(new_n220), .c(new_n223), .o1(\s[21] ));
  xnrc02aa1n02x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n221), .c(new_n220), .d(new_n222), .o1(new_n227));
  nand22aa1n03x5               g132(.a(new_n220), .b(new_n223), .o1(new_n228));
  nand42aa1n02x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\a[22] ), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\b[21] ), .o1(new_n231));
  aoi012aa1n06x5               g136(.a(new_n221), .b(new_n230), .c(new_n231), .o1(new_n232));
  nanp03aa1n02x5               g137(.a(new_n228), .b(new_n229), .c(new_n232), .o1(new_n233));
  nanp02aa1n02x5               g138(.a(new_n233), .b(new_n227), .o1(\s[22] ));
  nanb02aa1n06x5               g139(.a(new_n226), .b(new_n223), .out0(new_n235));
  nano32aa1n03x7               g140(.a(new_n235), .b(new_n199), .c(new_n201), .d(new_n209), .out0(new_n236));
  nanb02aa1n02x5               g141(.a(new_n211), .b(new_n217), .out0(new_n237));
  oai012aa1n02x5               g142(.a(new_n222), .b(\b[21] ), .c(\a[22] ), .o1(new_n238));
  nano23aa1n03x7               g143(.a(new_n238), .b(new_n221), .c(new_n210), .d(new_n229), .out0(new_n239));
  nanp02aa1n02x5               g144(.a(new_n237), .b(new_n239), .o1(new_n240));
  oaib12aa1n02x5               g145(.a(new_n240), .b(new_n232), .c(new_n229), .out0(new_n241));
  tech160nm_fixorc02aa1n03p5x5 g146(.a(\a[23] ), .b(\b[22] ), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n241), .c(new_n190), .d(new_n236), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n229), .b(new_n232), .out0(new_n244));
  nona22aa1n02x4               g149(.a(new_n240), .b(new_n244), .c(new_n242), .out0(new_n245));
  aoi012aa1n02x5               g150(.a(new_n245), .b(new_n190), .c(new_n236), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n243), .b(new_n246), .out0(\s[23] ));
  nor042aa1n03x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  inv000aa1n03x5               g153(.a(new_n248), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[24] ), .b(\b[23] ), .out0(new_n250));
  oai022aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n251));
  aoi012aa1n02x5               g156(.a(new_n251), .b(\a[24] ), .c(\b[23] ), .o1(new_n252));
  tech160nm_finand02aa1n03p5x5 g157(.a(new_n243), .b(new_n252), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n250), .c(new_n249), .d(new_n243), .o1(\s[24] ));
  norb02aa1n02x5               g159(.a(new_n223), .b(new_n226), .out0(new_n255));
  and002aa1n02x5               g160(.a(new_n250), .b(new_n242), .o(new_n256));
  nano22aa1n03x7               g161(.a(new_n216), .b(new_n256), .c(new_n255), .out0(new_n257));
  aoai13aa1n09x5               g162(.a(new_n256), .b(new_n244), .c(new_n237), .d(new_n239), .o1(new_n258));
  oaoi03aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(new_n258), .b(new_n260), .o1(new_n261));
  xnrc02aa1n12x5               g166(.a(\b[24] ), .b(\a[25] ), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n261), .c(new_n190), .d(new_n257), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n261), .c(new_n190), .d(new_n257), .o1(new_n265));
  norb02aa1n03x4               g170(.a(new_n264), .b(new_n265), .out0(\s[25] ));
  nor042aa1n03x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  inv000aa1n03x5               g172(.a(new_n267), .o1(new_n268));
  xorc02aa1n02x5               g173(.a(\a[26] ), .b(\b[25] ), .out0(new_n269));
  oai022aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n270));
  aoi012aa1n02x5               g175(.a(new_n270), .b(\a[26] ), .c(\b[25] ), .o1(new_n271));
  tech160nm_finand02aa1n05x5   g176(.a(new_n264), .b(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n269), .c(new_n268), .d(new_n264), .o1(\s[26] ));
  norb02aa1n09x5               g178(.a(new_n269), .b(new_n262), .out0(new_n274));
  nand03aa1n02x5               g179(.a(new_n236), .b(new_n256), .c(new_n274), .o1(new_n275));
  tech160nm_fiaoi012aa1n05x5   g180(.a(new_n275), .b(new_n185), .c(new_n184), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n275), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n274), .o1(new_n278));
  oaoi03aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .c(new_n268), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoai13aa1n12x5               g185(.a(new_n280), .b(new_n278), .c(new_n258), .d(new_n260), .o1(new_n281));
  xorc02aa1n02x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n281), .c(new_n190), .d(new_n277), .o1(new_n283));
  norp02aa1n02x5               g188(.a(new_n279), .b(new_n282), .o1(new_n284));
  aoai13aa1n02x5               g189(.a(new_n284), .b(new_n278), .c(new_n258), .d(new_n260), .o1(new_n285));
  oa0012aa1n03x5               g190(.a(new_n283), .b(new_n285), .c(new_n276), .o(\s[27] ));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  xorc02aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .out0(new_n289));
  oai022aa1d24x5               g194(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(\a[28] ), .c(\b[27] ), .o1(new_n291));
  tech160nm_finand02aa1n03p5x5 g196(.a(new_n283), .b(new_n291), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n289), .c(new_n288), .d(new_n283), .o1(\s[28] ));
  xorc02aa1n02x5               g198(.a(\a[29] ), .b(\b[28] ), .out0(new_n294));
  and002aa1n02x5               g199(.a(new_n289), .b(new_n282), .o(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n281), .c(new_n190), .d(new_n277), .o1(new_n296));
  inv000aa1d42x5               g201(.a(\b[27] ), .o1(new_n297));
  oaib12aa1n09x5               g202(.a(new_n290), .b(new_n297), .c(\a[28] ), .out0(new_n298));
  nanp03aa1n03x5               g203(.a(new_n296), .b(new_n298), .c(new_n294), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n298), .o1(new_n300));
  oaoi13aa1n02x5               g205(.a(new_n300), .b(new_n295), .c(new_n276), .d(new_n281), .o1(new_n301));
  oai012aa1n03x5               g206(.a(new_n299), .b(new_n301), .c(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g208(.a(new_n282), .b(new_n294), .c(new_n289), .o(new_n304));
  tech160nm_fioaoi03aa1n03p5x5 g209(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .o1(new_n305));
  oaoi13aa1n02x5               g210(.a(new_n305), .b(new_n304), .c(new_n276), .d(new_n281), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  aoai13aa1n02x5               g212(.a(new_n304), .b(new_n281), .c(new_n190), .d(new_n277), .o1(new_n308));
  norb02aa1n03x5               g213(.a(new_n307), .b(new_n305), .out0(new_n309));
  nand42aa1n02x5               g214(.a(new_n308), .b(new_n309), .o1(new_n310));
  oaih12aa1n02x5               g215(.a(new_n310), .b(new_n306), .c(new_n307), .o1(\s[30] ));
  and003aa1n02x5               g216(.a(new_n295), .b(new_n307), .c(new_n294), .o(new_n312));
  aoi012aa1n02x7               g217(.a(new_n309), .b(\a[30] ), .c(\b[29] ), .o1(new_n313));
  oaoi13aa1n02x5               g218(.a(new_n313), .b(new_n312), .c(new_n276), .d(new_n281), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[31] ), .b(\b[30] ), .out0(new_n315));
  aoai13aa1n02x5               g220(.a(new_n312), .b(new_n281), .c(new_n190), .d(new_n277), .o1(new_n316));
  norb02aa1n02x5               g221(.a(new_n315), .b(new_n313), .out0(new_n317));
  nand42aa1n02x5               g222(.a(new_n316), .b(new_n317), .o1(new_n318));
  oai012aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n321));
  aob012aa1n02x5               g226(.a(new_n107), .b(new_n321), .c(new_n105), .out0(\s[4] ));
  aob012aa1n02x5               g227(.a(new_n107), .b(\b[3] ), .c(\a[4] ), .out0(new_n323));
  nanb02aa1n02x5               g228(.a(new_n113), .b(new_n108), .out0(new_n324));
  nanp03aa1n02x5               g229(.a(new_n107), .b(new_n108), .c(new_n114), .o1(new_n325));
  aobi12aa1n02x5               g230(.a(new_n325), .b(new_n324), .c(new_n323), .out0(\s[5] ));
  obai22aa1n02x7               g231(.a(new_n325), .b(new_n113), .c(new_n121), .d(new_n116), .out0(new_n327));
  nanp02aa1n02x5               g232(.a(new_n325), .b(new_n122), .o1(new_n328));
  nanp02aa1n02x5               g233(.a(new_n327), .b(new_n328), .o1(\s[6] ));
  inv000aa1d42x5               g234(.a(new_n115), .o1(new_n330));
  nanp03aa1n03x5               g235(.a(new_n328), .b(new_n112), .c(new_n330), .o1(new_n331));
  xnrc02aa1n02x5               g236(.a(\b[6] ), .b(\a[7] ), .out0(new_n332));
  aoai13aa1n02x5               g237(.a(new_n332), .b(new_n121), .c(new_n325), .d(new_n122), .o1(new_n333));
  and002aa1n02x5               g238(.a(new_n331), .b(new_n333), .o(\s[7] ));
  xnbna2aa1n03x5               g239(.a(new_n111), .b(new_n331), .c(new_n330), .out0(\s[8] ));
  aoi112aa1n02x5               g240(.a(new_n125), .b(new_n123), .c(new_n107), .d(new_n118), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n126), .b(new_n336), .out0(\s[9] ));
endmodule


