// Benchmark "adder" written by ABC on Wed Jul 17 19:02:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n329, new_n330, new_n332, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  oai022aa1d24x5               g002(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n98));
  xorc02aa1n12x5               g003(.a(\a[7] ), .b(\b[6] ), .out0(new_n99));
  aoi022aa1n06x5               g004(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n100));
  orn002aa1n12x5               g005(.a(\a[7] ), .b(\b[6] ), .o(new_n101));
  oaoi03aa1n09x5               g006(.a(\a[8] ), .b(\b[7] ), .c(new_n101), .o1(new_n102));
  aoi013aa1n09x5               g007(.a(new_n102), .b(new_n99), .c(new_n100), .d(new_n98), .o1(new_n103));
  nor002aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  inv000aa1n02x5               g009(.a(new_n104), .o1(new_n105));
  nanp02aa1n04x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  aob012aa1n02x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .out0(new_n108));
  nor042aa1n03x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  nand02aa1n03x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  norb02aa1n03x5               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  nor042aa1n02x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nand42aa1n02x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  norb02aa1n03x5               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  nand03aa1n04x5               g019(.a(new_n108), .b(new_n111), .c(new_n114), .o1(new_n115));
  tech160nm_fiaoi012aa1n04x5   g020(.a(new_n109), .b(new_n112), .c(new_n110), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nanp03aa1n02x5               g022(.a(new_n99), .b(new_n100), .c(new_n117), .o1(new_n118));
  aoai13aa1n12x5               g023(.a(new_n103), .b(new_n118), .c(new_n115), .d(new_n116), .o1(new_n119));
  xorc02aa1n02x5               g024(.a(\a[9] ), .b(\b[8] ), .out0(new_n120));
  nanp02aa1n02x5               g025(.a(new_n119), .b(new_n120), .o1(new_n121));
  oaib12aa1n02x5               g026(.a(new_n121), .b(\b[8] ), .c(new_n97), .out0(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1n10x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  nor042aa1n06x5               g029(.a(\b[10] ), .b(\a[11] ), .o1(new_n125));
  norb02aa1n06x5               g030(.a(new_n124), .b(new_n125), .out0(new_n126));
  oai022aa1d24x5               g031(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  aoi022aa1n02x5               g033(.a(new_n121), .b(new_n128), .c(\b[9] ), .d(\a[10] ), .o1(new_n129));
  nand42aa1n03x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nano22aa1n02x4               g035(.a(new_n125), .b(new_n130), .c(new_n124), .out0(new_n131));
  aoai13aa1n06x5               g036(.a(new_n131), .b(new_n127), .c(new_n119), .d(new_n120), .o1(new_n132));
  oa0012aa1n02x5               g037(.a(new_n132), .b(new_n129), .c(new_n126), .o(\s[11] ));
  oai012aa1n02x5               g038(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  aoi012aa1n02x5               g040(.a(new_n104), .b(new_n106), .c(new_n107), .o1(new_n136));
  nona23aa1n09x5               g041(.a(new_n113), .b(new_n110), .c(new_n109), .d(new_n112), .out0(new_n137));
  oai012aa1n03x5               g042(.a(new_n116), .b(new_n137), .c(new_n136), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n98), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(\b[6] ), .b(\a[7] ), .o1(new_n140));
  nanp03aa1n02x5               g045(.a(new_n100), .b(new_n101), .c(new_n140), .o1(new_n141));
  nano23aa1n02x4               g046(.a(new_n102), .b(new_n141), .c(new_n139), .d(new_n117), .out0(new_n142));
  nand42aa1n02x5               g047(.a(new_n142), .b(new_n138), .o1(new_n143));
  aoi022aa1d24x5               g048(.a(\b[9] ), .b(\a[10] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n144));
  inv000aa1d42x5               g049(.a(\a[12] ), .o1(new_n145));
  inv000aa1d42x5               g050(.a(\b[11] ), .o1(new_n146));
  oao003aa1n03x5               g051(.a(new_n145), .b(new_n146), .c(new_n125), .carry(new_n147));
  aoi013aa1n09x5               g052(.a(new_n147), .b(new_n126), .c(new_n127), .d(new_n144), .o1(new_n148));
  and002aa1n02x5               g053(.a(\b[8] ), .b(\a[9] ), .o(new_n149));
  nand42aa1n03x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nano32aa1n03x7               g055(.a(new_n125), .b(new_n150), .c(new_n130), .d(new_n124), .out0(new_n151));
  oaoi03aa1n09x5               g056(.a(new_n145), .b(new_n146), .c(new_n125), .o1(new_n152));
  nona23aa1d18x5               g057(.a(new_n151), .b(new_n152), .c(new_n127), .d(new_n149), .out0(new_n153));
  aoai13aa1n02x5               g058(.a(new_n148), .b(new_n153), .c(new_n143), .d(new_n103), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g060(.a(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(\b[12] ), .o1(new_n157));
  oaoi03aa1n02x5               g062(.a(new_n156), .b(new_n157), .c(new_n154), .o1(new_n158));
  xnrb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g064(.a(new_n148), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n153), .o1(new_n161));
  nor002aa1n02x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nor022aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nano23aa1n03x7               g070(.a(new_n162), .b(new_n164), .c(new_n165), .d(new_n163), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n160), .c(new_n119), .d(new_n161), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n165), .b(new_n164), .c(new_n156), .d(new_n157), .o1(new_n168));
  nor002aa1n16x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand42aa1n10x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nanb02aa1d24x5               g075(.a(new_n169), .b(new_n170), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n167), .c(new_n168), .out0(\s[15] ));
  nanp02aa1n02x5               g078(.a(new_n167), .b(new_n168), .o1(new_n174));
  orn002aa1n02x5               g079(.a(\a[16] ), .b(\b[15] ), .o(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(new_n175), .b(new_n176), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n169), .c(new_n174), .d(new_n170), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(new_n174), .b(new_n172), .o1(new_n179));
  nona22aa1n02x4               g084(.a(new_n179), .b(new_n177), .c(new_n169), .out0(new_n180));
  nanp02aa1n02x5               g085(.a(new_n180), .b(new_n178), .o1(\s[16] ));
  nona23aa1n02x4               g086(.a(new_n165), .b(new_n163), .c(new_n162), .d(new_n164), .out0(new_n182));
  norp03aa1n02x5               g087(.a(new_n182), .b(new_n171), .c(new_n177), .o1(new_n183));
  nanb02aa1n03x5               g088(.a(new_n153), .b(new_n183), .out0(new_n184));
  inv000aa1d42x5               g089(.a(new_n169), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n170), .o1(new_n186));
  aoai13aa1n02x5               g091(.a(new_n175), .b(new_n186), .c(new_n168), .d(new_n185), .o1(new_n187));
  aboi22aa1n03x5               g092(.a(new_n148), .b(new_n183), .c(new_n187), .d(new_n176), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n184), .c(new_n143), .d(new_n103), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g095(.a(\a[18] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[16] ), .o1(new_n193));
  oaoi03aa1n03x5               g098(.a(new_n192), .b(new_n193), .c(new_n189), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[17] ), .c(new_n191), .out0(\s[18] ));
  nona22aa1n03x5               g100(.a(new_n166), .b(new_n177), .c(new_n171), .out0(new_n196));
  nor042aa1n04x5               g101(.a(new_n153), .b(new_n196), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n187), .b(new_n176), .o1(new_n198));
  oai012aa1n12x5               g103(.a(new_n198), .b(new_n148), .c(new_n196), .o1(new_n199));
  xroi22aa1d06x4               g104(.a(new_n192), .b(\b[16] ), .c(new_n191), .d(\b[17] ), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n199), .c(new_n119), .d(new_n197), .o1(new_n201));
  nand02aa1d04x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  oai022aa1d18x5               g107(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n203), .b(new_n202), .o1(new_n204));
  nor002aa1n10x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand22aa1n06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  norb02aa1n09x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n201), .c(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n03p5x5 g114(.a(new_n201), .b(new_n204), .o1(new_n210));
  xnrc02aa1n02x5               g115(.a(\b[19] ), .b(\a[20] ), .out0(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n205), .c(new_n210), .d(new_n206), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n204), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n207), .b(new_n213), .c(new_n189), .d(new_n200), .o1(new_n214));
  nona22aa1n03x5               g119(.a(new_n214), .b(new_n211), .c(new_n205), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n212), .b(new_n215), .o1(\s[20] ));
  nanb03aa1d18x5               g121(.a(new_n211), .b(new_n200), .c(new_n207), .out0(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n199), .c(new_n119), .d(new_n197), .o1(new_n219));
  inv000aa1d48x5               g124(.a(new_n205), .o1(new_n220));
  orn002aa1n24x5               g125(.a(\a[20] ), .b(\b[19] ), .o(new_n221));
  and002aa1n12x5               g126(.a(\b[19] ), .b(\a[20] ), .o(new_n222));
  nanp03aa1d12x5               g127(.a(new_n203), .b(new_n202), .c(new_n206), .o1(new_n223));
  aoai13aa1n12x5               g128(.a(new_n221), .b(new_n222), .c(new_n223), .d(new_n220), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  norp02aa1n04x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  nand42aa1n03x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  norb02aa1n06x4               g132(.a(new_n227), .b(new_n226), .out0(new_n228));
  xnbna2aa1n03x5               g133(.a(new_n228), .b(new_n219), .c(new_n225), .out0(\s[21] ));
  nand42aa1n03x5               g134(.a(new_n219), .b(new_n225), .o1(new_n230));
  nor042aa1n04x5               g135(.a(\b[21] ), .b(\a[22] ), .o1(new_n231));
  nand42aa1n06x5               g136(.a(\b[21] ), .b(\a[22] ), .o1(new_n232));
  norb02aa1n15x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n226), .c(new_n230), .d(new_n228), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n228), .b(new_n224), .c(new_n189), .d(new_n218), .o1(new_n236));
  nona22aa1n03x5               g141(.a(new_n236), .b(new_n234), .c(new_n226), .out0(new_n237));
  nanp02aa1n02x5               g142(.a(new_n235), .b(new_n237), .o1(\s[22] ));
  nano23aa1n09x5               g143(.a(new_n226), .b(new_n231), .c(new_n232), .d(new_n227), .out0(new_n239));
  nano32aa1n02x4               g144(.a(new_n211), .b(new_n200), .c(new_n239), .d(new_n207), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n199), .c(new_n119), .d(new_n197), .o1(new_n241));
  oai022aa1n06x5               g146(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n242));
  aoi022aa1n02x5               g147(.a(new_n224), .b(new_n239), .c(new_n232), .d(new_n242), .o1(new_n243));
  norp02aa1n04x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  nand02aa1n03x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  norb02aa1n06x4               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  xnbna2aa1n03x5               g151(.a(new_n246), .b(new_n241), .c(new_n243), .out0(\s[23] ));
  nand22aa1n03x5               g152(.a(new_n241), .b(new_n243), .o1(new_n248));
  nor002aa1n02x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  nanb02aa1n02x5               g155(.a(new_n249), .b(new_n250), .out0(new_n251));
  aoai13aa1n02x5               g156(.a(new_n251), .b(new_n244), .c(new_n248), .d(new_n245), .o1(new_n252));
  inv000aa1n02x5               g157(.a(new_n243), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n246), .b(new_n253), .c(new_n189), .d(new_n240), .o1(new_n254));
  nona22aa1n03x5               g159(.a(new_n254), .b(new_n251), .c(new_n244), .out0(new_n255));
  nanp02aa1n02x5               g160(.a(new_n252), .b(new_n255), .o1(\s[24] ));
  nano23aa1n06x5               g161(.a(new_n244), .b(new_n249), .c(new_n250), .d(new_n245), .out0(new_n257));
  nano22aa1n03x7               g162(.a(new_n217), .b(new_n239), .c(new_n257), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n199), .c(new_n119), .d(new_n197), .o1(new_n259));
  nano32aa1n09x5               g164(.a(new_n251), .b(new_n246), .c(new_n233), .d(new_n228), .out0(new_n260));
  aoai13aa1n02x5               g165(.a(new_n245), .b(new_n244), .c(new_n242), .d(new_n232), .o1(new_n261));
  oaoi03aa1n09x5               g166(.a(\a[24] ), .b(\b[23] ), .c(new_n261), .o1(new_n262));
  aoi012aa1d24x5               g167(.a(new_n262), .b(new_n224), .c(new_n260), .o1(new_n263));
  tech160nm_fixorc02aa1n04x5   g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n259), .c(new_n263), .out0(\s[25] ));
  nand22aa1n02x5               g170(.a(new_n259), .b(new_n263), .o1(new_n266));
  norp02aa1n02x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n266), .d(new_n264), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n263), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n264), .b(new_n270), .c(new_n189), .d(new_n258), .o1(new_n271));
  nona22aa1n02x5               g176(.a(new_n271), .b(new_n268), .c(new_n267), .out0(new_n272));
  nanp02aa1n02x5               g177(.a(new_n269), .b(new_n272), .o1(\s[26] ));
  norb02aa1n03x5               g178(.a(new_n264), .b(new_n268), .out0(new_n274));
  nano32aa1d12x5               g179(.a(new_n217), .b(new_n274), .c(new_n239), .d(new_n257), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n199), .c(new_n119), .d(new_n197), .o1(new_n276));
  aoi013aa1n02x4               g181(.a(new_n205), .b(new_n203), .c(new_n202), .d(new_n206), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(new_n257), .b(new_n239), .o1(new_n278));
  oaoi13aa1n02x5               g183(.a(new_n278), .b(new_n221), .c(new_n277), .d(new_n222), .o1(new_n279));
  inv000aa1d42x5               g184(.a(\a[26] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(\b[25] ), .o1(new_n281));
  tech160nm_fioaoi03aa1n03p5x5 g186(.a(new_n280), .b(new_n281), .c(new_n267), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  oaoi13aa1n04x5               g188(.a(new_n283), .b(new_n274), .c(new_n279), .d(new_n262), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n284), .c(new_n276), .out0(\s[27] ));
  tech160nm_finand02aa1n03p5x5 g191(.a(new_n284), .b(new_n276), .o1(new_n287));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  norp02aa1n02x5               g193(.a(\b[27] ), .b(\a[28] ), .o1(new_n289));
  nand42aa1n03x5               g194(.a(\b[27] ), .b(\a[28] ), .o1(new_n290));
  nanb02aa1n09x5               g195(.a(new_n289), .b(new_n290), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n288), .c(new_n287), .d(new_n285), .o1(new_n292));
  oaib12aa1n06x5               g197(.a(new_n282), .b(new_n263), .c(new_n274), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n285), .b(new_n293), .c(new_n189), .d(new_n275), .o1(new_n294));
  nona22aa1n03x5               g199(.a(new_n294), .b(new_n291), .c(new_n288), .out0(new_n295));
  nanp02aa1n03x5               g200(.a(new_n292), .b(new_n295), .o1(\s[28] ));
  norb02aa1n03x5               g201(.a(new_n285), .b(new_n291), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n293), .c(new_n189), .d(new_n275), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n297), .o1(new_n299));
  oai012aa1n02x5               g204(.a(new_n290), .b(new_n289), .c(new_n288), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n299), .c(new_n284), .d(new_n276), .o1(new_n301));
  norp02aa1n02x5               g206(.a(\b[28] ), .b(\a[29] ), .o1(new_n302));
  nanp02aa1n02x5               g207(.a(\b[28] ), .b(\a[29] ), .o1(new_n303));
  norb02aa1n02x5               g208(.a(new_n303), .b(new_n302), .out0(new_n304));
  oai022aa1n02x5               g209(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n305));
  aboi22aa1n03x5               g210(.a(new_n302), .b(new_n303), .c(new_n305), .d(new_n290), .out0(new_n306));
  aoi022aa1n03x5               g211(.a(new_n301), .b(new_n304), .c(new_n298), .d(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g213(.a(new_n291), .b(new_n285), .c(new_n304), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n293), .c(new_n189), .d(new_n275), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n309), .o1(new_n311));
  aoi013aa1n02x4               g216(.a(new_n302), .b(new_n305), .c(new_n290), .d(new_n303), .o1(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n311), .c(new_n284), .d(new_n276), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  aoi113aa1n02x5               g219(.a(new_n314), .b(new_n302), .c(new_n305), .d(new_n303), .e(new_n290), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n310), .d(new_n315), .o1(\s[30] ));
  nanp03aa1n02x5               g221(.a(new_n297), .b(new_n304), .c(new_n314), .o1(new_n317));
  nanb02aa1n03x5               g222(.a(new_n317), .b(new_n287), .out0(new_n318));
  xorc02aa1n02x5               g223(.a(\a[31] ), .b(\b[30] ), .out0(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n320), .b(new_n317), .c(new_n284), .d(new_n276), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n318), .b(new_n321), .c(new_n322), .d(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n136), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi112aa1n02x5               g229(.a(new_n112), .b(new_n111), .c(new_n108), .d(new_n114), .o1(new_n325));
  aoib12aa1n02x5               g230(.a(new_n325), .b(new_n138), .c(new_n109), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n138), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  xorc02aa1n02x5               g232(.a(\a[5] ), .b(\b[4] ), .out0(new_n328));
  nanp02aa1n02x5               g233(.a(new_n138), .b(new_n328), .o1(new_n329));
  oa0012aa1n02x5               g234(.a(new_n329), .b(\b[4] ), .c(\a[5] ), .o(new_n330));
  xnrb03aa1n02x5               g235(.a(new_n330), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi022aa1n02x5               g236(.a(new_n329), .b(new_n139), .c(\a[6] ), .d(\b[5] ), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aobi12aa1n02x5               g238(.a(new_n101), .b(new_n332), .c(new_n140), .out0(new_n334));
  xnrb03aa1n02x5               g239(.a(new_n334), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g240(.a(new_n119), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


