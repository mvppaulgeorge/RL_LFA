// Benchmark "adder" written by ABC on Thu Jul 18 09:32:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n318, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n342, new_n343, new_n344,
    new_n346, new_n348, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n357, new_n358, new_n360, new_n361;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand03aa1n03x5               g003(.a(new_n98), .b(\a[1] ), .c(\b[0] ), .o1(new_n99));
  nor042aa1n04x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nand02aa1n08x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norb02aa1n12x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  nor042aa1d18x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1d28x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano22aa1n03x7               g009(.a(new_n103), .b(new_n98), .c(new_n104), .out0(new_n105));
  oai112aa1n06x5               g010(.a(new_n105), .b(new_n102), .c(new_n99), .d(new_n97), .o1(new_n106));
  tech160nm_fioai012aa1n04x5   g011(.a(new_n101), .b(new_n103), .c(new_n100), .o1(new_n107));
  nand02aa1d10x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nor002aa1n03x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nand02aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nano23aa1n06x5               g016(.a(new_n110), .b(new_n109), .c(new_n111), .d(new_n108), .out0(new_n112));
  norp02aa1n24x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1d28x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanb02aa1n03x5               g019(.a(new_n113), .b(new_n114), .out0(new_n115));
  nor002aa1d32x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand22aa1n12x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nanb02aa1n12x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  nona22aa1n09x5               g023(.a(new_n112), .b(new_n115), .c(new_n118), .out0(new_n119));
  norb02aa1n06x4               g024(.a(new_n114), .b(new_n113), .out0(new_n120));
  nano22aa1n03x7               g025(.a(new_n116), .b(new_n108), .c(new_n117), .out0(new_n121));
  oaih22aa1n04x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  nor042aa1n02x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  oa0012aa1n03x5               g028(.a(new_n114), .b(new_n116), .c(new_n113), .o(new_n124));
  aoi113aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(new_n121), .d(new_n122), .e(new_n120), .o1(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n119), .c(new_n106), .d(new_n107), .o1(new_n126));
  nor022aa1n04x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n16x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n09x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  nand42aa1n03x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n130), .b(new_n126), .c(new_n131), .out0(\s[10] ));
  nand42aa1n16x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nano22aa1n02x4               g039(.a(new_n134), .b(new_n128), .c(new_n133), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n130), .c(new_n126), .d(new_n131), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n134), .b(new_n133), .out0(new_n137));
  aoai13aa1n02x5               g042(.a(new_n128), .b(new_n130), .c(new_n126), .d(new_n131), .o1(new_n138));
  aobi12aa1n02x5               g043(.a(new_n136), .b(new_n138), .c(new_n137), .out0(\s[11] ));
  inv000aa1d42x5               g044(.a(new_n134), .o1(new_n140));
  norp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1n10x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  nona23aa1n02x4               g048(.a(new_n136), .b(new_n142), .c(new_n141), .d(new_n134), .out0(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n143), .c(new_n140), .d(new_n136), .o1(\s[12] ));
  aoi013aa1n06x4               g050(.a(new_n124), .b(new_n121), .c(new_n122), .d(new_n120), .o1(new_n146));
  aoai13aa1n12x5               g051(.a(new_n146), .b(new_n119), .c(new_n106), .d(new_n107), .o1(new_n147));
  nano23aa1n03x7               g052(.a(new_n141), .b(new_n134), .c(new_n142), .d(new_n133), .out0(new_n148));
  norb02aa1n03x5               g053(.a(new_n131), .b(new_n123), .out0(new_n149));
  and003aa1n02x5               g054(.a(new_n148), .b(new_n129), .c(new_n149), .o(new_n150));
  nanp02aa1n03x5               g055(.a(new_n147), .b(new_n150), .o1(new_n151));
  aoi012aa1n02x5               g056(.a(new_n134), .b(\a[10] ), .c(\b[9] ), .o1(new_n152));
  nano22aa1n03x5               g057(.a(new_n141), .b(new_n133), .c(new_n142), .out0(new_n153));
  oai112aa1n03x5               g058(.a(new_n153), .b(new_n152), .c(new_n127), .d(new_n123), .o1(new_n154));
  oai012aa1n02x5               g059(.a(new_n142), .b(new_n141), .c(new_n134), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n154), .b(new_n155), .o1(new_n156));
  nanb02aa1n03x5               g061(.a(new_n156), .b(new_n151), .out0(new_n157));
  nor042aa1n09x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nanp02aa1n02x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(new_n160));
  and003aa1n02x5               g065(.a(new_n154), .b(new_n160), .c(new_n155), .o(new_n161));
  aboi22aa1n03x5               g066(.a(new_n160), .b(new_n157), .c(new_n161), .d(new_n151), .out0(\s[13] ));
  inv000aa1d42x5               g067(.a(new_n158), .o1(new_n163));
  nanb02aa1n03x5               g068(.a(new_n160), .b(new_n157), .out0(new_n164));
  nor002aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nanp02aa1n04x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  oaih22aa1d12x5               g072(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n168));
  nanb03aa1n02x5               g073(.a(new_n168), .b(new_n164), .c(new_n166), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n167), .c(new_n163), .d(new_n164), .o1(\s[14] ));
  nano23aa1n06x5               g075(.a(new_n158), .b(new_n165), .c(new_n166), .d(new_n159), .out0(new_n171));
  aoai13aa1n02x5               g076(.a(new_n171), .b(new_n156), .c(new_n147), .d(new_n150), .o1(new_n172));
  oaoi03aa1n02x5               g077(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  xorc02aa1n12x5               g079(.a(\a[15] ), .b(\b[14] ), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n172), .c(new_n174), .out0(\s[15] ));
  orn002aa1n02x5               g081(.a(\a[15] ), .b(\b[14] ), .o(new_n177));
  aob012aa1n03x5               g082(.a(new_n175), .b(new_n172), .c(new_n174), .out0(new_n178));
  xorc02aa1n02x5               g083(.a(\a[16] ), .b(\b[15] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n175), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\a[16] ), .o1(new_n181));
  nanb02aa1n12x5               g086(.a(\b[15] ), .b(new_n181), .out0(new_n182));
  nanp02aa1n02x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  and003aa1n02x5               g088(.a(new_n177), .b(new_n182), .c(new_n183), .o(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n180), .c(new_n172), .d(new_n174), .o1(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n179), .c(new_n178), .d(new_n177), .o1(\s[16] ));
  nand23aa1n06x5               g091(.a(new_n171), .b(new_n175), .c(new_n179), .o1(new_n187));
  nano32aa1n06x5               g092(.a(new_n187), .b(new_n149), .c(new_n148), .d(new_n129), .out0(new_n188));
  nand02aa1n03x5               g093(.a(new_n147), .b(new_n188), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(\b[14] ), .b(\a[15] ), .o1(new_n190));
  nanp03aa1n02x5               g095(.a(new_n182), .b(new_n190), .c(new_n183), .o1(new_n191));
  oai112aa1n02x5               g096(.a(new_n168), .b(new_n166), .c(\b[14] ), .d(\a[15] ), .o1(new_n192));
  oaoi03aa1n02x5               g097(.a(\a[16] ), .b(\b[15] ), .c(new_n177), .o1(new_n193));
  oab012aa1n02x4               g098(.a(new_n193), .b(new_n192), .c(new_n191), .out0(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n187), .c(new_n154), .d(new_n155), .o1(new_n195));
  inv000aa1n06x5               g100(.a(new_n195), .o1(new_n196));
  nand22aa1n09x5               g101(.a(new_n189), .b(new_n196), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  norp02aa1n02x5               g103(.a(new_n193), .b(new_n198), .o1(new_n199));
  oai012aa1n02x5               g104(.a(new_n199), .b(new_n192), .c(new_n191), .o1(new_n200));
  aoib12aa1n02x5               g105(.a(new_n200), .b(new_n156), .c(new_n187), .out0(new_n201));
  aoi022aa1n02x5               g106(.a(new_n197), .b(new_n198), .c(new_n189), .d(new_n201), .o1(\s[17] ));
  nor002aa1d32x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n02x5               g109(.a(new_n198), .b(new_n195), .c(new_n147), .d(new_n188), .o1(new_n205));
  xorc02aa1n12x5               g110(.a(\a[18] ), .b(\b[17] ), .out0(new_n206));
  nand42aa1n02x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nor002aa1n02x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  norp02aa1n03x5               g113(.a(new_n208), .b(new_n203), .o1(new_n209));
  nanp03aa1n02x5               g114(.a(new_n205), .b(new_n207), .c(new_n209), .o1(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n206), .c(new_n204), .d(new_n205), .o1(\s[18] ));
  and002aa1n02x5               g116(.a(new_n206), .b(new_n198), .o(new_n212));
  oaoi03aa1n02x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n213));
  xorc02aa1n02x5               g118(.a(\a[19] ), .b(\b[18] ), .out0(new_n214));
  aoai13aa1n06x5               g119(.a(new_n214), .b(new_n213), .c(new_n197), .d(new_n212), .o1(new_n215));
  aoi112aa1n02x5               g120(.a(new_n214), .b(new_n213), .c(new_n197), .d(new_n212), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n215), .b(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g123(.a(\a[19] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(\b[18] ), .o1(new_n220));
  nand02aa1d12x5               g125(.a(new_n220), .b(new_n219), .o1(new_n221));
  nor042aa1n03x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand42aa1n06x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  nano22aa1n02x4               g129(.a(new_n222), .b(new_n221), .c(new_n223), .out0(new_n225));
  nanp02aa1n03x5               g130(.a(new_n215), .b(new_n225), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n224), .c(new_n221), .d(new_n215), .o1(\s[20] ));
  nand42aa1n03x5               g132(.a(\b[18] ), .b(\a[19] ), .o1(new_n228));
  nano32aa1n03x7               g133(.a(new_n222), .b(new_n221), .c(new_n223), .d(new_n228), .out0(new_n229));
  nand23aa1n06x5               g134(.a(new_n229), .b(new_n198), .c(new_n206), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  nano22aa1n03x7               g136(.a(new_n222), .b(new_n228), .c(new_n223), .out0(new_n232));
  oai012aa1n03x5               g137(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .o1(new_n233));
  nona22aa1n09x5               g138(.a(new_n232), .b(new_n209), .c(new_n233), .out0(new_n234));
  oaoi03aa1n09x5               g139(.a(\a[20] ), .b(\b[19] ), .c(new_n221), .o1(new_n235));
  inv000aa1n02x5               g140(.a(new_n235), .o1(new_n236));
  nanp02aa1n02x5               g141(.a(new_n234), .b(new_n236), .o1(new_n237));
  tech160nm_fixorc02aa1n02p5x5 g142(.a(\a[21] ), .b(\b[20] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n237), .c(new_n197), .d(new_n231), .o1(new_n239));
  nona22aa1n02x4               g144(.a(new_n234), .b(new_n235), .c(new_n238), .out0(new_n240));
  aoi012aa1n02x5               g145(.a(new_n240), .b(new_n197), .c(new_n231), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n239), .b(new_n241), .out0(\s[21] ));
  norp02aa1n02x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  xorc02aa1n02x5               g149(.a(\a[22] ), .b(\b[21] ), .out0(new_n245));
  oai022aa1n02x5               g150(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(\a[22] ), .c(\b[21] ), .o1(new_n247));
  nanp02aa1n03x5               g152(.a(new_n239), .b(new_n247), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n248), .b(new_n245), .c(new_n244), .d(new_n239), .o1(\s[22] ));
  nand02aa1n02x5               g154(.a(new_n245), .b(new_n238), .o1(new_n250));
  nano32aa1n02x4               g155(.a(new_n250), .b(new_n229), .c(new_n206), .d(new_n198), .out0(new_n251));
  inv000aa1d42x5               g156(.a(\b[21] ), .o1(new_n252));
  oaib12aa1n02x5               g157(.a(new_n246), .b(new_n252), .c(\a[22] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n250), .c(new_n234), .d(new_n236), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n197), .d(new_n251), .o1(new_n256));
  aoai13aa1n02x5               g161(.a(new_n251), .b(new_n195), .c(new_n147), .d(new_n188), .o1(new_n257));
  oab012aa1n02x4               g162(.a(new_n233), .b(new_n203), .c(new_n208), .out0(new_n258));
  inv000aa1d42x5               g163(.a(\b[20] ), .o1(new_n259));
  xroi22aa1d04x5               g164(.a(new_n252), .b(\a[22] ), .c(new_n259), .d(\a[21] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n235), .c(new_n258), .d(new_n232), .o1(new_n261));
  nano32aa1n02x4               g166(.a(new_n255), .b(new_n257), .c(new_n261), .d(new_n253), .out0(new_n262));
  norb02aa1n02x5               g167(.a(new_n256), .b(new_n262), .out0(\s[23] ));
  nor042aa1n03x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  inv020aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .out0(new_n266));
  oai022aa1n02x5               g171(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n267));
  aoi012aa1n02x5               g172(.a(new_n267), .b(\a[24] ), .c(\b[23] ), .o1(new_n268));
  nanp02aa1n03x5               g173(.a(new_n256), .b(new_n268), .o1(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n266), .c(new_n265), .d(new_n256), .o1(\s[24] ));
  tech160nm_fixnrc02aa1n04x5   g175(.a(\b[23] ), .b(\a[24] ), .out0(new_n271));
  norb02aa1n12x5               g176(.a(new_n255), .b(new_n271), .out0(new_n272));
  nano22aa1n02x4               g177(.a(new_n230), .b(new_n272), .c(new_n260), .out0(new_n273));
  inv000aa1d42x5               g178(.a(new_n272), .o1(new_n274));
  tech160nm_fioaoi03aa1n02p5x5 g179(.a(\a[24] ), .b(\b[23] ), .c(new_n265), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n274), .c(new_n261), .d(new_n253), .o1(new_n277));
  tech160nm_fixorc02aa1n03p5x5 g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n197), .d(new_n273), .o1(new_n279));
  aoi112aa1n02x5               g184(.a(new_n278), .b(new_n275), .c(new_n254), .d(new_n272), .o1(new_n280));
  aobi12aa1n02x5               g185(.a(new_n280), .b(new_n273), .c(new_n197), .out0(new_n281));
  norb02aa1n03x4               g186(.a(new_n279), .b(new_n281), .out0(\s[25] ));
  norp02aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[26] ), .b(\b[25] ), .out0(new_n285));
  oai022aa1n02x5               g190(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n286));
  aoi012aa1n02x5               g191(.a(new_n286), .b(\a[26] ), .c(\b[25] ), .o1(new_n287));
  nanp02aa1n03x5               g192(.a(new_n279), .b(new_n287), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n285), .c(new_n284), .d(new_n279), .o1(\s[26] ));
  and002aa1n02x5               g194(.a(new_n285), .b(new_n278), .o(new_n290));
  nano32aa1n03x7               g195(.a(new_n230), .b(new_n290), .c(new_n260), .d(new_n272), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n195), .c(new_n147), .d(new_n188), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n290), .b(new_n275), .c(new_n254), .d(new_n272), .o1(new_n293));
  aob012aa1n02x5               g198(.a(new_n286), .b(\b[25] ), .c(\a[26] ), .out0(new_n294));
  nand23aa1n06x5               g199(.a(new_n292), .b(new_n293), .c(new_n294), .o1(new_n295));
  xorc02aa1n12x5               g200(.a(\a[27] ), .b(\b[26] ), .out0(new_n296));
  inv000aa1d42x5               g201(.a(new_n296), .o1(new_n297));
  and003aa1n02x5               g202(.a(new_n293), .b(new_n297), .c(new_n294), .o(new_n298));
  aoi022aa1n02x5               g203(.a(new_n298), .b(new_n292), .c(new_n295), .d(new_n296), .o1(\s[27] ));
  norp02aa1n02x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n295), .b(new_n296), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .out0(new_n303));
  aobi12aa1n02x7               g208(.a(new_n294), .b(new_n277), .c(new_n290), .out0(new_n304));
  oai022aa1n02x5               g209(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n305));
  aoi012aa1n02x5               g210(.a(new_n305), .b(\a[28] ), .c(\b[27] ), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n306), .b(new_n297), .c(new_n304), .d(new_n292), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n302), .d(new_n301), .o1(\s[28] ));
  and002aa1n02x5               g213(.a(new_n303), .b(new_n296), .o(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  aob012aa1n09x5               g215(.a(new_n305), .b(\b[27] ), .c(\a[28] ), .out0(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[28] ), .b(\a[29] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n311), .b(new_n312), .out0(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n310), .c(new_n304), .d(new_n292), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n311), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n312), .b(new_n315), .c(new_n295), .d(new_n309), .o1(new_n316));
  nanp02aa1n03x5               g221(.a(new_n316), .b(new_n314), .o1(\s[29] ));
  nanp02aa1n02x5               g222(.a(\b[0] ), .b(\a[1] ), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g224(.a(new_n312), .b(new_n296), .c(new_n303), .out0(new_n320));
  oaoi03aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .o1(new_n321));
  norp02aa1n02x5               g226(.a(\b[29] ), .b(\a[30] ), .o1(new_n322));
  nanp02aa1n02x5               g227(.a(\b[29] ), .b(\a[30] ), .o1(new_n323));
  nanb02aa1n02x5               g228(.a(new_n322), .b(new_n323), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n321), .c(new_n295), .d(new_n320), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n320), .o1(new_n326));
  nanp02aa1n02x5               g231(.a(\b[28] ), .b(\a[29] ), .o1(new_n327));
  oai012aa1n02x5               g232(.a(new_n311), .b(\b[28] ), .c(\a[29] ), .o1(new_n328));
  aoi012aa1n02x5               g233(.a(new_n324), .b(new_n328), .c(new_n327), .o1(new_n329));
  aoai13aa1n02x5               g234(.a(new_n329), .b(new_n326), .c(new_n304), .d(new_n292), .o1(new_n330));
  nanp02aa1n03x5               g235(.a(new_n325), .b(new_n330), .o1(\s[30] ));
  nano23aa1n02x5               g236(.a(new_n324), .b(new_n312), .c(new_n303), .d(new_n296), .out0(new_n332));
  nanp02aa1n03x5               g237(.a(new_n295), .b(new_n332), .o1(new_n333));
  inv000aa1n02x5               g238(.a(new_n332), .o1(new_n334));
  nano22aa1n02x4               g239(.a(new_n322), .b(new_n327), .c(new_n323), .out0(new_n335));
  oai022aa1n02x5               g240(.a(\a[30] ), .b(\b[29] ), .c(\b[30] ), .d(\a[31] ), .o1(new_n336));
  aoi122aa1n03x5               g241(.a(new_n336), .b(\b[30] ), .c(\a[31] ), .d(new_n328), .e(new_n335), .o1(new_n337));
  aoai13aa1n02x5               g242(.a(new_n337), .b(new_n334), .c(new_n304), .d(new_n292), .o1(new_n338));
  aoi012aa1n02x5               g243(.a(new_n322), .b(new_n328), .c(new_n335), .o1(new_n339));
  xorc02aa1n02x5               g244(.a(\a[31] ), .b(\b[30] ), .out0(new_n340));
  aoai13aa1n03x5               g245(.a(new_n338), .b(new_n340), .c(new_n333), .d(new_n339), .o1(\s[31] ));
  oai012aa1n02x5               g246(.a(new_n105), .b(new_n99), .c(new_n97), .o1(new_n342));
  oai012aa1n02x5               g247(.a(new_n98), .b(new_n97), .c(new_n318), .o1(new_n343));
  oaib12aa1n02x5               g248(.a(new_n343), .b(new_n103), .c(new_n104), .out0(new_n344));
  and002aa1n02x5               g249(.a(new_n342), .b(new_n344), .o(\s[3] ));
  inv000aa1d42x5               g250(.a(new_n103), .o1(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n102), .b(new_n342), .c(new_n346), .out0(\s[4] ));
  norb02aa1n02x5               g252(.a(new_n111), .b(new_n110), .out0(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n348), .b(new_n106), .c(new_n107), .out0(\s[5] ));
  norb02aa1n02x5               g254(.a(new_n108), .b(new_n109), .out0(new_n350));
  nanp02aa1n02x5               g255(.a(new_n106), .b(new_n107), .o1(new_n351));
  aoi012aa1n02x5               g256(.a(new_n110), .b(new_n351), .c(new_n111), .o1(new_n352));
  norb03aa1n02x5               g257(.a(new_n108), .b(new_n110), .c(new_n109), .out0(new_n353));
  aob012aa1n02x5               g258(.a(new_n353), .b(new_n351), .c(new_n348), .out0(new_n354));
  oai012aa1n02x5               g259(.a(new_n354), .b(new_n352), .c(new_n350), .o1(\s[6] ));
  xnbna2aa1n03x5               g260(.a(new_n118), .b(new_n354), .c(new_n108), .out0(\s[7] ));
  aoai13aa1n02x5               g261(.a(new_n115), .b(new_n116), .c(new_n354), .d(new_n121), .o1(new_n357));
  nona22aa1n02x4               g262(.a(new_n114), .b(new_n116), .c(new_n113), .out0(new_n358));
  aoai13aa1n02x5               g263(.a(new_n357), .b(new_n358), .c(new_n354), .d(new_n121), .o1(\s[8] ));
  nanb02aa1n02x5               g264(.a(new_n119), .b(new_n351), .out0(new_n360));
  aoi113aa1n02x5               g265(.a(new_n149), .b(new_n124), .c(new_n121), .d(new_n122), .e(new_n120), .o1(new_n361));
  aoi022aa1n02x5               g266(.a(new_n361), .b(new_n360), .c(new_n147), .d(new_n149), .o1(\s[9] ));
endmodule


