// Benchmark "adder" written by ABC on Wed Jul 17 20:40:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n355, new_n357, new_n360, new_n361,
    new_n363, new_n364, new_n366, new_n368, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n08x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand42aa1n06x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  norb03aa1n09x5               g004(.a(new_n98), .b(new_n97), .c(new_n99), .out0(new_n100));
  inv030aa1n04x5               g005(.a(new_n100), .o1(new_n101));
  tech160nm_fixnrc02aa1n04x5   g006(.a(\b[3] ), .b(\a[4] ), .out0(new_n102));
  nor042aa1n09x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb03aa1n12x5               g009(.a(new_n103), .b(new_n104), .c(new_n98), .out0(new_n105));
  nona22aa1n09x5               g010(.a(new_n101), .b(new_n105), .c(new_n102), .out0(new_n106));
  inv000aa1d42x5               g011(.a(new_n103), .o1(new_n107));
  oao003aa1n02x5               g012(.a(\a[4] ), .b(\b[3] ), .c(new_n107), .carry(new_n108));
  xnrc02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .out0(new_n109));
  tech160nm_fixorc02aa1n03p5x5 g014(.a(\a[5] ), .b(\b[4] ), .out0(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .out0(new_n111));
  nor042aa1n06x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand42aa1n06x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  norb02aa1n02x7               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  nona23aa1n06x5               g019(.a(new_n114), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n115));
  xorc02aa1n12x5               g020(.a(\a[8] ), .b(\b[7] ), .out0(new_n116));
  nand42aa1n03x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nano22aa1n02x4               g022(.a(new_n112), .b(new_n117), .c(new_n113), .out0(new_n118));
  norp02aa1n04x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  oab012aa1n04x5               g024(.a(new_n119), .b(\a[6] ), .c(\b[5] ), .out0(new_n120));
  inv000aa1n02x5               g025(.a(new_n120), .o1(new_n121));
  inv040aa1n06x5               g026(.a(new_n112), .o1(new_n122));
  oaoi03aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  aoi013aa1n06x4               g028(.a(new_n123), .b(new_n118), .c(new_n116), .d(new_n121), .o1(new_n124));
  aoai13aa1n12x5               g029(.a(new_n124), .b(new_n115), .c(new_n106), .d(new_n108), .o1(new_n125));
  xnrc02aa1n12x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  inv000aa1d42x5               g031(.a(new_n126), .o1(new_n127));
  nor002aa1n02x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nor002aa1n12x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1n06x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n128), .c(new_n125), .d(new_n127), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n129), .o1(new_n133));
  oai112aa1n02x5               g038(.a(new_n133), .b(new_n130), .c(\b[8] ), .d(\a[9] ), .o1(new_n134));
  aoai13aa1n02x5               g039(.a(new_n132), .b(new_n134), .c(new_n127), .d(new_n125), .o1(\s[10] ));
  oai013aa1n09x5               g040(.a(new_n108), .b(new_n100), .c(new_n105), .d(new_n102), .o1(new_n136));
  xorc02aa1n02x5               g041(.a(\a[6] ), .b(\b[5] ), .out0(new_n137));
  nano32aa1n03x7               g042(.a(new_n111), .b(new_n110), .c(new_n137), .d(new_n114), .out0(new_n138));
  nanp03aa1n02x5               g043(.a(new_n118), .b(new_n116), .c(new_n121), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n123), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(new_n139), .b(new_n140), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n126), .b(new_n131), .o1(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n141), .c(new_n138), .d(new_n136), .o1(new_n143));
  oai012aa1n02x5               g048(.a(new_n130), .b(new_n129), .c(new_n128), .o1(new_n144));
  tech160nm_fixorc02aa1n03p5x5 g049(.a(\a[11] ), .b(\b[10] ), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n143), .c(new_n144), .out0(\s[11] ));
  inv040aa1d32x5               g051(.a(\a[11] ), .o1(new_n147));
  inv000aa1d42x5               g052(.a(\b[10] ), .o1(new_n148));
  nanp02aa1n04x5               g053(.a(new_n148), .b(new_n147), .o1(new_n149));
  aob012aa1n02x5               g054(.a(new_n145), .b(new_n143), .c(new_n144), .out0(new_n150));
  norp02aa1n02x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nand42aa1n03x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  norb02aa1n03x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  nano22aa1n02x4               g058(.a(new_n151), .b(new_n149), .c(new_n152), .out0(new_n154));
  nanp02aa1n02x5               g059(.a(new_n150), .b(new_n154), .o1(new_n155));
  aoai13aa1n02x5               g060(.a(new_n155), .b(new_n153), .c(new_n149), .d(new_n150), .o1(\s[12] ));
  nona23aa1d18x5               g061(.a(new_n153), .b(new_n145), .c(new_n126), .d(new_n131), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nand42aa1n02x5               g063(.a(\b[10] ), .b(\a[11] ), .o1(new_n159));
  nano22aa1n02x4               g064(.a(new_n151), .b(new_n159), .c(new_n152), .out0(new_n160));
  oai012aa1n02x5               g065(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .o1(new_n161));
  oab012aa1n04x5               g066(.a(new_n161), .b(new_n128), .c(new_n129), .out0(new_n162));
  oaoi03aa1n12x5               g067(.a(\a[12] ), .b(\b[11] ), .c(new_n149), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  aob012aa1n02x5               g069(.a(new_n164), .b(new_n162), .c(new_n160), .out0(new_n165));
  nor002aa1n10x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n165), .c(new_n125), .d(new_n158), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n163), .b(new_n168), .c(new_n162), .d(new_n160), .o1(new_n170));
  aobi12aa1n02x5               g075(.a(new_n170), .b(new_n125), .c(new_n158), .out0(new_n171));
  norb02aa1n02x5               g076(.a(new_n169), .b(new_n171), .out0(\s[13] ));
  inv000aa1d42x5               g077(.a(new_n166), .o1(new_n173));
  nor042aa1n02x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nand42aa1n02x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  oai022aa1n02x5               g081(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n177));
  nanb03aa1n02x5               g082(.a(new_n177), .b(new_n169), .c(new_n175), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n176), .c(new_n173), .d(new_n169), .o1(\s[14] ));
  nano23aa1n06x5               g084(.a(new_n166), .b(new_n174), .c(new_n175), .d(new_n167), .out0(new_n180));
  nanp03aa1n02x5               g085(.a(new_n125), .b(new_n158), .c(new_n180), .o1(new_n181));
  aoi022aa1n02x5               g086(.a(new_n165), .b(new_n180), .c(new_n175), .d(new_n177), .o1(new_n182));
  nor002aa1n03x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  nanp02aa1n02x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norb02aa1n02x5               g089(.a(new_n184), .b(new_n183), .out0(new_n185));
  aob012aa1n03x5               g090(.a(new_n185), .b(new_n181), .c(new_n182), .out0(new_n186));
  oai012aa1n06x5               g091(.a(new_n175), .b(new_n174), .c(new_n166), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(new_n185), .b(new_n188), .c(new_n165), .d(new_n180), .o1(new_n189));
  aobi12aa1n02x5               g094(.a(new_n186), .b(new_n189), .c(new_n181), .out0(\s[15] ));
  inv000aa1n02x5               g095(.a(new_n183), .o1(new_n191));
  xnrc02aa1n12x5               g096(.a(\b[15] ), .b(\a[16] ), .out0(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\a[16] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[15] ), .o1(new_n195));
  aoi012aa1n02x5               g100(.a(new_n183), .b(new_n194), .c(new_n195), .o1(new_n196));
  oai112aa1n02x5               g101(.a(new_n186), .b(new_n196), .c(new_n195), .d(new_n194), .o1(new_n197));
  aoai13aa1n02x5               g102(.a(new_n197), .b(new_n193), .c(new_n191), .d(new_n186), .o1(\s[16] ));
  nano22aa1n12x5               g103(.a(new_n192), .b(new_n191), .c(new_n184), .out0(new_n199));
  nano22aa1d15x5               g104(.a(new_n157), .b(new_n180), .c(new_n199), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n141), .c(new_n136), .d(new_n138), .o1(new_n201));
  oaoi03aa1n02x5               g106(.a(new_n194), .b(new_n195), .c(new_n183), .o1(new_n202));
  aoai13aa1n04x5               g107(.a(new_n180), .b(new_n163), .c(new_n162), .d(new_n160), .o1(new_n203));
  aob012aa1n06x5               g108(.a(new_n199), .b(new_n203), .c(new_n187), .out0(new_n204));
  nand23aa1n06x5               g109(.a(new_n201), .b(new_n202), .c(new_n204), .o1(new_n205));
  tech160nm_fixorc02aa1n03p5x5 g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  nano22aa1n02x4               g111(.a(new_n206), .b(new_n204), .c(new_n202), .out0(new_n207));
  aoi022aa1n02x5               g112(.a(new_n207), .b(new_n201), .c(new_n205), .d(new_n206), .o1(\s[17] ));
  nor002aa1d32x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n199), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n202), .b(new_n211), .c(new_n203), .d(new_n187), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n206), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n213));
  nor042aa1n04x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  nand42aa1n06x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  norb02aa1n02x7               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  nona23aa1n02x4               g121(.a(new_n213), .b(new_n215), .c(new_n214), .d(new_n209), .out0(new_n217));
  aoai13aa1n02x5               g122(.a(new_n217), .b(new_n216), .c(new_n210), .d(new_n213), .o1(\s[18] ));
  and002aa1n02x5               g123(.a(new_n206), .b(new_n216), .o(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n220));
  oaoi03aa1n02x5               g125(.a(\a[18] ), .b(\b[17] ), .c(new_n210), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[19] ), .b(\b[18] ), .out0(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n220), .c(new_n222), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g130(.a(\a[19] ), .o1(new_n226));
  inv040aa1d28x5               g131(.a(\b[18] ), .o1(new_n227));
  nand02aa1d24x5               g132(.a(new_n227), .b(new_n226), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n223), .b(new_n221), .c(new_n205), .d(new_n219), .o1(new_n229));
  nor042aa1n02x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nanp02aa1n04x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n223), .o1(new_n233));
  nano22aa1n02x4               g138(.a(new_n230), .b(new_n228), .c(new_n231), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n233), .c(new_n220), .d(new_n222), .o1(new_n235));
  aoai13aa1n02x5               g140(.a(new_n235), .b(new_n232), .c(new_n229), .d(new_n228), .o1(\s[20] ));
  nand42aa1n02x5               g141(.a(\b[18] ), .b(\a[19] ), .o1(new_n237));
  nano32aa1n02x4               g142(.a(new_n230), .b(new_n228), .c(new_n231), .d(new_n237), .out0(new_n238));
  nand23aa1n06x5               g143(.a(new_n238), .b(new_n206), .c(new_n216), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n241));
  nano22aa1n03x7               g146(.a(new_n230), .b(new_n237), .c(new_n231), .out0(new_n242));
  oai012aa1n02x7               g147(.a(new_n215), .b(\b[18] ), .c(\a[19] ), .o1(new_n243));
  oab012aa1n04x5               g148(.a(new_n243), .b(new_n209), .c(new_n214), .out0(new_n244));
  nanp02aa1n02x5               g149(.a(new_n244), .b(new_n242), .o1(new_n245));
  oaoi03aa1n12x5               g150(.a(\a[20] ), .b(\b[19] ), .c(new_n228), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  nanp02aa1n02x5               g152(.a(new_n245), .b(new_n247), .o1(new_n248));
  nor022aa1n16x5               g153(.a(\b[20] ), .b(\a[21] ), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[20] ), .b(\a[21] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n250), .b(new_n249), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n248), .c(new_n205), .d(new_n240), .o1(new_n252));
  aoi112aa1n02x5               g157(.a(new_n246), .b(new_n251), .c(new_n244), .d(new_n242), .o1(new_n253));
  aobi12aa1n03x7               g158(.a(new_n252), .b(new_n253), .c(new_n241), .out0(\s[21] ));
  inv000aa1d42x5               g159(.a(new_n249), .o1(new_n255));
  nor042aa1n03x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  nanp02aa1n06x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n248), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n251), .o1(new_n260));
  norb03aa1n02x5               g165(.a(new_n257), .b(new_n249), .c(new_n256), .out0(new_n261));
  aoai13aa1n02x5               g166(.a(new_n261), .b(new_n260), .c(new_n241), .d(new_n259), .o1(new_n262));
  aoai13aa1n02x5               g167(.a(new_n262), .b(new_n258), .c(new_n252), .d(new_n255), .o1(\s[22] ));
  nano23aa1n06x5               g168(.a(new_n249), .b(new_n256), .c(new_n257), .d(new_n250), .out0(new_n264));
  norb02aa1n03x5               g169(.a(new_n264), .b(new_n239), .out0(new_n265));
  aoai13aa1n02x5               g170(.a(new_n265), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n266));
  aoai13aa1n12x5               g171(.a(new_n264), .b(new_n246), .c(new_n244), .d(new_n242), .o1(new_n267));
  oai012aa1n12x5               g172(.a(new_n257), .b(new_n256), .c(new_n249), .o1(new_n268));
  nand02aa1d06x5               g173(.a(new_n267), .b(new_n268), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[23] ), .b(\b[22] ), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n205), .d(new_n265), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n270), .o1(new_n272));
  and003aa1n02x5               g177(.a(new_n267), .b(new_n272), .c(new_n268), .o(new_n273));
  aobi12aa1n02x5               g178(.a(new_n271), .b(new_n273), .c(new_n266), .out0(\s[23] ));
  norp02aa1n02x5               g179(.a(\b[22] ), .b(\a[23] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[24] ), .b(\b[23] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n269), .o1(new_n278));
  oai022aa1n02x5               g183(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n279));
  aoi012aa1n02x5               g184(.a(new_n279), .b(\a[24] ), .c(\b[23] ), .o1(new_n280));
  aoai13aa1n02x7               g185(.a(new_n280), .b(new_n272), .c(new_n266), .d(new_n278), .o1(new_n281));
  aoai13aa1n02x5               g186(.a(new_n281), .b(new_n277), .c(new_n271), .d(new_n276), .o1(\s[24] ));
  nano32aa1n02x5               g187(.a(new_n239), .b(new_n277), .c(new_n264), .d(new_n270), .out0(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n284));
  and002aa1n02x7               g189(.a(new_n277), .b(new_n270), .o(new_n285));
  inv020aa1n02x5               g190(.a(new_n285), .o1(new_n286));
  aob012aa1n02x5               g191(.a(new_n279), .b(\b[23] ), .c(\a[24] ), .out0(new_n287));
  aoai13aa1n12x5               g192(.a(new_n287), .b(new_n286), .c(new_n267), .d(new_n268), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[25] ), .b(\b[24] ), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n288), .c(new_n205), .d(new_n283), .o1(new_n290));
  nand22aa1n03x5               g195(.a(new_n269), .b(new_n285), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n289), .o1(new_n292));
  and003aa1n02x5               g197(.a(new_n291), .b(new_n287), .c(new_n292), .o(new_n293));
  aobi12aa1n02x5               g198(.a(new_n290), .b(new_n293), .c(new_n284), .out0(\s[25] ));
  norp02aa1n02x5               g199(.a(\b[24] ), .b(\a[25] ), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[26] ), .b(\b[25] ), .out0(new_n297));
  inv000aa1d42x5               g202(.a(new_n288), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(\b[25] ), .b(\a[26] ), .o1(new_n299));
  oai022aa1n02x5               g204(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n300));
  norb02aa1n02x5               g205(.a(new_n299), .b(new_n300), .out0(new_n301));
  aoai13aa1n02x7               g206(.a(new_n301), .b(new_n292), .c(new_n284), .d(new_n298), .o1(new_n302));
  aoai13aa1n02x5               g207(.a(new_n302), .b(new_n297), .c(new_n290), .d(new_n296), .o1(\s[26] ));
  and002aa1n06x5               g208(.a(new_n297), .b(new_n289), .o(new_n304));
  inv000aa1n02x5               g209(.a(new_n304), .o1(new_n305));
  nano23aa1n06x5               g210(.a(new_n305), .b(new_n239), .c(new_n285), .d(new_n264), .out0(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n212), .c(new_n125), .d(new_n200), .o1(new_n307));
  nanp02aa1n02x5               g212(.a(new_n300), .b(new_n299), .o1(new_n308));
  aoai13aa1n04x5               g213(.a(new_n308), .b(new_n305), .c(new_n291), .d(new_n287), .o1(new_n309));
  tech160nm_fixorc02aa1n03p5x5 g214(.a(\a[27] ), .b(\b[26] ), .out0(new_n310));
  aoai13aa1n06x5               g215(.a(new_n310), .b(new_n309), .c(new_n205), .d(new_n306), .o1(new_n311));
  aoi122aa1n02x5               g216(.a(new_n310), .b(new_n299), .c(new_n300), .d(new_n288), .e(new_n304), .o1(new_n312));
  aobi12aa1n02x5               g217(.a(new_n311), .b(new_n312), .c(new_n307), .out0(\s[27] ));
  norp02aa1n02x5               g218(.a(\b[26] ), .b(\a[27] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .out0(new_n316));
  aoi022aa1d18x5               g221(.a(new_n288), .b(new_n304), .c(new_n299), .d(new_n300), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n310), .o1(new_n318));
  oai022aa1n02x5               g223(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n319), .b(\a[28] ), .c(\b[27] ), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n318), .c(new_n307), .d(new_n317), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n316), .c(new_n311), .d(new_n315), .o1(\s[28] ));
  and002aa1n02x5               g227(.a(new_n316), .b(new_n310), .o(new_n323));
  inv000aa1d42x5               g228(.a(new_n323), .o1(new_n324));
  aob012aa1n02x5               g229(.a(new_n319), .b(\b[27] ), .c(\a[28] ), .out0(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[28] ), .b(\a[29] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n325), .b(new_n326), .out0(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n324), .c(new_n307), .d(new_n317), .o1(new_n328));
  aoai13aa1n06x5               g233(.a(new_n325), .b(new_n324), .c(new_n307), .d(new_n317), .o1(new_n329));
  nanp02aa1n03x5               g234(.a(new_n329), .b(new_n326), .o1(new_n330));
  nanp02aa1n03x5               g235(.a(new_n330), .b(new_n328), .o1(\s[29] ));
  xorb03aa1n02x5               g236(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g237(.a(new_n326), .b(new_n310), .c(new_n316), .out0(new_n333));
  nanp02aa1n02x5               g238(.a(\b[28] ), .b(\a[29] ), .o1(new_n334));
  oai012aa1n02x5               g239(.a(new_n325), .b(\b[28] ), .c(\a[29] ), .o1(new_n335));
  nanp02aa1n02x5               g240(.a(new_n335), .b(new_n334), .o1(new_n336));
  aoai13aa1n06x5               g241(.a(new_n336), .b(new_n333), .c(new_n307), .d(new_n317), .o1(new_n337));
  norp02aa1n02x5               g242(.a(\b[29] ), .b(\a[30] ), .o1(new_n338));
  nanp02aa1n02x5               g243(.a(\b[29] ), .b(\a[30] ), .o1(new_n339));
  nanb02aa1n02x5               g244(.a(new_n338), .b(new_n339), .out0(new_n340));
  nanp02aa1n03x5               g245(.a(new_n337), .b(new_n340), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n340), .b(new_n335), .c(new_n334), .o1(new_n342));
  aoai13aa1n03x5               g247(.a(new_n342), .b(new_n333), .c(new_n307), .d(new_n317), .o1(new_n343));
  nanp02aa1n03x5               g248(.a(new_n341), .b(new_n343), .o1(\s[30] ));
  nano23aa1d12x5               g249(.a(new_n340), .b(new_n326), .c(new_n316), .d(new_n310), .out0(new_n345));
  aoai13aa1n02x5               g250(.a(new_n345), .b(new_n309), .c(new_n205), .d(new_n306), .o1(new_n346));
  inv000aa1d42x5               g251(.a(new_n345), .o1(new_n347));
  nano22aa1n02x4               g252(.a(new_n338), .b(new_n334), .c(new_n339), .out0(new_n348));
  oai022aa1n02x5               g253(.a(\a[30] ), .b(\b[29] ), .c(\b[30] ), .d(\a[31] ), .o1(new_n349));
  aoi122aa1n02x5               g254(.a(new_n349), .b(\b[30] ), .c(\a[31] ), .d(new_n335), .e(new_n348), .o1(new_n350));
  aoai13aa1n03x5               g255(.a(new_n350), .b(new_n347), .c(new_n307), .d(new_n317), .o1(new_n351));
  aoi012aa1n02x5               g256(.a(new_n338), .b(new_n335), .c(new_n348), .o1(new_n352));
  xorc02aa1n02x5               g257(.a(\a[31] ), .b(\b[30] ), .out0(new_n353));
  aoai13aa1n03x5               g258(.a(new_n351), .b(new_n353), .c(new_n346), .d(new_n352), .o1(\s[31] ));
  norb02aa1n02x5               g259(.a(new_n104), .b(new_n103), .out0(new_n355));
  xobna2aa1n03x5               g260(.a(new_n355), .b(new_n101), .c(new_n98), .out0(\s[3] ));
  oai112aa1n02x5               g261(.a(new_n355), .b(new_n98), .c(new_n99), .d(new_n97), .o1(new_n357));
  xobna2aa1n03x5               g262(.a(new_n102), .b(new_n357), .c(new_n107), .out0(\s[4] ));
  xnbna2aa1n03x5               g263(.a(new_n110), .b(new_n106), .c(new_n108), .out0(\s[5] ));
  aoai13aa1n02x5               g264(.a(new_n109), .b(new_n119), .c(new_n136), .d(new_n110), .o1(new_n360));
  oai012aa1n02x5               g265(.a(new_n137), .b(\b[4] ), .c(\a[5] ), .o1(new_n361));
  aoai13aa1n02x5               g266(.a(new_n360), .b(new_n361), .c(new_n110), .d(new_n136), .o1(\s[6] ));
  nanb02aa1n02x5               g267(.a(new_n120), .b(new_n117), .out0(new_n363));
  nanp03aa1n02x5               g268(.a(new_n136), .b(new_n137), .c(new_n110), .o1(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n114), .b(new_n364), .c(new_n363), .out0(\s[7] ));
  aob012aa1n02x5               g270(.a(new_n114), .b(new_n364), .c(new_n363), .out0(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n116), .b(new_n366), .c(new_n122), .out0(\s[8] ));
  nanp02aa1n02x5               g272(.a(new_n138), .b(new_n136), .o1(new_n368));
  aoi113aa1n02x5               g273(.a(new_n127), .b(new_n123), .c(new_n118), .d(new_n116), .e(new_n121), .o1(new_n369));
  aoi022aa1n02x5               g274(.a(new_n125), .b(new_n127), .c(new_n368), .d(new_n369), .o1(\s[9] ));
endmodule


