// Benchmark "adder" written by ABC on Wed Jul 17 17:24:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n325, new_n327,
    new_n328, new_n330;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n02x5               g001(.a(\b[3] ), .b(\a[4] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  nor002aa1n02x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  aoi012aa1n02x5               g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[1] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  oaoi03aa1n02x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n02x4               g010(.a(new_n105), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n106));
  tech160nm_fioai012aa1n04x5   g011(.a(new_n100), .b(new_n106), .c(new_n104), .o1(new_n107));
  oaih22aa1d12x5               g012(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(new_n108), .o1(new_n109));
  and002aa1n06x5               g014(.a(\b[6] ), .b(\a[7] ), .o(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand22aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor022aa1n06x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand22aa1n02x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  norp02aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nona23aa1n09x5               g020(.a(new_n114), .b(new_n112), .c(new_n115), .d(new_n113), .out0(new_n116));
  nano23aa1n06x5               g021(.a(new_n116), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n117));
  oai012aa1n02x5               g022(.a(new_n112), .b(new_n115), .c(new_n113), .o1(new_n118));
  oai013aa1n09x5               g023(.a(new_n118), .b(new_n116), .c(new_n109), .d(new_n110), .o1(new_n119));
  xorc02aa1n02x5               g024(.a(\a[9] ), .b(\b[8] ), .out0(new_n120));
  aoai13aa1n02x5               g025(.a(new_n120), .b(new_n119), .c(new_n117), .d(new_n107), .o1(new_n121));
  xorc02aa1n12x5               g026(.a(\a[10] ), .b(\b[9] ), .out0(new_n122));
  inv000aa1d42x5               g027(.a(new_n122), .o1(new_n123));
  oaoi13aa1n04x5               g028(.a(new_n123), .b(new_n121), .c(\a[9] ), .d(\b[8] ), .o1(new_n124));
  nor002aa1d24x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  oao003aa1n02x5               g030(.a(new_n101), .b(new_n102), .c(new_n103), .carry(new_n126));
  nano23aa1n02x4               g031(.a(new_n97), .b(new_n99), .c(new_n105), .d(new_n98), .out0(new_n127));
  aobi12aa1n02x5               g032(.a(new_n100), .b(new_n127), .c(new_n126), .out0(new_n128));
  nano23aa1n06x5               g033(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n129));
  nona23aa1n02x4               g034(.a(new_n129), .b(new_n111), .c(new_n108), .d(new_n110), .out0(new_n130));
  norb02aa1n02x5               g035(.a(new_n108), .b(new_n110), .out0(new_n131));
  aobi12aa1n02x5               g036(.a(new_n118), .b(new_n129), .c(new_n131), .out0(new_n132));
  oai012aa1n06x5               g037(.a(new_n132), .b(new_n128), .c(new_n130), .o1(new_n133));
  aoi112aa1n02x5               g038(.a(new_n122), .b(new_n125), .c(new_n133), .d(new_n120), .o1(new_n134));
  norp02aa1n02x5               g039(.a(new_n124), .b(new_n134), .o1(\s[10] ));
  inv000aa1d42x5               g040(.a(\a[10] ), .o1(new_n136));
  inv020aa1d32x5               g041(.a(\b[9] ), .o1(new_n137));
  oaoi03aa1n12x5               g042(.a(new_n136), .b(new_n137), .c(new_n125), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  nand42aa1n20x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  nor022aa1n06x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  oai022aa1n02x5               g047(.a(new_n124), .b(new_n139), .c(new_n142), .d(new_n141), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n140), .b(new_n142), .out0(new_n144));
  nano22aa1n02x4               g049(.a(new_n124), .b(new_n138), .c(new_n144), .out0(new_n145));
  nanb02aa1n02x5               g050(.a(new_n145), .b(new_n143), .out0(\s[11] ));
  norp02aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  tech160nm_finand02aa1n05x5   g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  tech160nm_fioai012aa1n02p5x5 g054(.a(new_n149), .b(new_n145), .c(new_n141), .o1(new_n150));
  nor043aa1n03x5               g055(.a(new_n145), .b(new_n149), .c(new_n141), .o1(new_n151));
  nanb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(\s[12] ));
  nano23aa1n02x4               g057(.a(new_n147), .b(new_n142), .c(new_n148), .d(new_n140), .out0(new_n153));
  nanp03aa1n03x5               g058(.a(new_n153), .b(new_n120), .c(new_n122), .o1(new_n154));
  nanb02aa1n06x5               g059(.a(new_n154), .b(new_n133), .out0(new_n155));
  nona23aa1n09x5               g060(.a(new_n140), .b(new_n148), .c(new_n147), .d(new_n142), .out0(new_n156));
  tech160nm_fioai012aa1n03p5x5 g061(.a(new_n148), .b(new_n147), .c(new_n142), .o1(new_n157));
  oai012aa1d24x5               g062(.a(new_n157), .b(new_n156), .c(new_n138), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  xorc02aa1n12x5               g064(.a(\a[13] ), .b(\b[12] ), .out0(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n155), .c(new_n159), .out0(\s[13] ));
  nor042aa1d18x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  inv020aa1n04x5               g067(.a(new_n162), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(new_n155), .b(new_n159), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(new_n164), .b(new_n160), .o1(new_n165));
  xorc02aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n165), .c(new_n163), .out0(\s[14] ));
  nanp02aa1n02x5               g072(.a(new_n166), .b(new_n160), .o1(new_n168));
  oaoi03aa1n12x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n04x5               g075(.a(new_n170), .b(new_n168), .c(new_n155), .d(new_n159), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor022aa1n08x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n10x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  nor002aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nand42aa1n06x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n173), .c(new_n171), .d(new_n175), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(new_n171), .b(new_n175), .o1(new_n180));
  nona22aa1n02x4               g085(.a(new_n180), .b(new_n178), .c(new_n173), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n181), .b(new_n179), .o1(\s[16] ));
  nano23aa1n03x5               g087(.a(new_n176), .b(new_n173), .c(new_n177), .d(new_n174), .out0(new_n183));
  nand23aa1n03x5               g088(.a(new_n183), .b(new_n160), .c(new_n166), .o1(new_n184));
  nor042aa1n03x5               g089(.a(new_n184), .b(new_n154), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n185), .b(new_n119), .c(new_n117), .d(new_n107), .o1(new_n186));
  norb02aa1n03x5               g091(.a(new_n183), .b(new_n168), .out0(new_n187));
  tech160nm_fiao0012aa1n02p5x5 g092(.a(new_n176), .b(new_n173), .c(new_n177), .o(new_n188));
  aoi012aa1n02x7               g093(.a(new_n188), .b(new_n183), .c(new_n169), .o1(new_n189));
  aobi12aa1n12x5               g094(.a(new_n189), .b(new_n187), .c(new_n158), .out0(new_n190));
  nand02aa1d08x5               g095(.a(new_n186), .b(new_n190), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[18] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  oaoi03aa1n02x5               g100(.a(new_n194), .b(new_n195), .c(new_n191), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  xroi22aa1d04x5               g102(.a(new_n194), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n198));
  norp02aa1n02x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  aoi013aa1n09x5               g105(.a(new_n199), .b(new_n200), .c(new_n194), .d(new_n195), .o1(new_n201));
  aob012aa1n03x5               g106(.a(new_n201), .b(new_n191), .c(new_n198), .out0(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanp02aa1n02x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  nor002aa1n03x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand22aa1n03x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n205), .c(new_n202), .d(new_n207), .o1(new_n211));
  nona22aa1n02x4               g116(.a(new_n200), .b(\b[16] ), .c(\a[17] ), .out0(new_n212));
  oaib12aa1n02x5               g117(.a(new_n212), .b(\b[17] ), .c(new_n193), .out0(new_n213));
  aoai13aa1n02x5               g118(.a(new_n207), .b(new_n213), .c(new_n191), .d(new_n198), .o1(new_n214));
  nona22aa1n02x4               g119(.a(new_n214), .b(new_n210), .c(new_n205), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n211), .b(new_n215), .o1(\s[20] ));
  nano23aa1n06x5               g121(.a(new_n208), .b(new_n205), .c(new_n209), .d(new_n206), .out0(new_n217));
  nanp02aa1n02x5               g122(.a(new_n198), .b(new_n217), .o1(new_n218));
  nona23aa1n09x5               g123(.a(new_n206), .b(new_n209), .c(new_n208), .d(new_n205), .out0(new_n219));
  oai012aa1n06x5               g124(.a(new_n209), .b(new_n208), .c(new_n205), .o1(new_n220));
  oai012aa1n18x5               g125(.a(new_n220), .b(new_n219), .c(new_n201), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n222), .b(new_n218), .c(new_n186), .d(new_n190), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xorc02aa1n02x5               g130(.a(\a[21] ), .b(\b[20] ), .out0(new_n226));
  xorc02aa1n02x5               g131(.a(\a[22] ), .b(\b[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n226), .o1(new_n229));
  aoi112aa1n02x5               g134(.a(new_n225), .b(new_n228), .c(new_n223), .d(new_n226), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(\s[22] ));
  inv000aa1d42x5               g136(.a(\a[21] ), .o1(new_n232));
  inv040aa1d32x5               g137(.a(\a[22] ), .o1(new_n233));
  xroi22aa1d06x4               g138(.a(new_n232), .b(\b[20] ), .c(new_n233), .d(\b[21] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(\b[21] ), .o1(new_n235));
  oao003aa1n02x5               g140(.a(new_n233), .b(new_n235), .c(new_n225), .carry(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n221), .c(new_n234), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n234), .o1(new_n238));
  nona22aa1n09x5               g143(.a(new_n191), .b(new_n218), .c(new_n238), .out0(new_n239));
  xnrc02aa1n02x5               g144(.a(\b[22] ), .b(\a[23] ), .out0(new_n240));
  xobna2aa1n03x5               g145(.a(new_n240), .b(new_n239), .c(new_n237), .out0(\s[23] ));
  and002aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o(new_n242));
  xorc02aa1n12x5               g147(.a(\a[24] ), .b(\b[23] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  inv000aa1n02x5               g149(.a(new_n220), .o1(new_n245));
  aoai13aa1n06x5               g150(.a(new_n234), .b(new_n245), .c(new_n217), .d(new_n213), .o1(new_n246));
  norp02aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  nona22aa1n02x4               g152(.a(new_n246), .b(new_n236), .c(new_n247), .out0(new_n248));
  inv040aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n244), .b(new_n242), .c(new_n239), .d(new_n249), .o1(new_n250));
  aoi112aa1n03x5               g155(.a(new_n244), .b(new_n242), .c(new_n239), .d(new_n249), .o1(new_n251));
  norb02aa1n03x4               g156(.a(new_n250), .b(new_n251), .out0(\s[24] ));
  oaib12aa1n03x5               g157(.a(new_n189), .b(new_n184), .c(new_n158), .out0(new_n253));
  norb02aa1n03x5               g158(.a(new_n243), .b(new_n240), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n218), .b(new_n254), .c(new_n234), .out0(new_n255));
  aoai13aa1n02x5               g160(.a(new_n255), .b(new_n253), .c(new_n133), .d(new_n185), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n254), .b(new_n236), .c(new_n221), .d(new_n234), .o1(new_n257));
  inv000aa1n03x5               g162(.a(new_n247), .o1(new_n258));
  oaoi03aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n258), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  nanp03aa1n03x5               g165(.a(new_n256), .b(new_n257), .c(new_n260), .o1(new_n261));
  xorb03aa1n02x5               g166(.a(new_n261), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  nor002aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .o1(new_n265));
  nand42aa1n03x5               g170(.a(\b[25] ), .b(\a[26] ), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n266), .b(new_n265), .out0(new_n267));
  inv040aa1n03x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n263), .c(new_n261), .d(new_n264), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n236), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n254), .o1(new_n271));
  aoai13aa1n04x5               g176(.a(new_n260), .b(new_n271), .c(new_n246), .d(new_n270), .o1(new_n272));
  aoai13aa1n02x5               g177(.a(new_n264), .b(new_n272), .c(new_n191), .d(new_n255), .o1(new_n273));
  nona22aa1n02x4               g178(.a(new_n273), .b(new_n268), .c(new_n263), .out0(new_n274));
  nanp02aa1n02x5               g179(.a(new_n269), .b(new_n274), .o1(\s[26] ));
  norb02aa1n03x5               g180(.a(new_n264), .b(new_n268), .out0(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  nano23aa1n06x5               g182(.a(new_n277), .b(new_n218), .c(new_n254), .d(new_n234), .out0(new_n278));
  aoai13aa1n04x5               g183(.a(new_n278), .b(new_n253), .c(new_n133), .d(new_n185), .o1(new_n279));
  oai012aa1n02x5               g184(.a(new_n266), .b(new_n265), .c(new_n263), .o1(new_n280));
  aobi12aa1n06x5               g185(.a(new_n280), .b(new_n272), .c(new_n276), .out0(new_n281));
  norp02aa1n02x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  norb02aa1n02x5               g188(.a(new_n283), .b(new_n282), .out0(new_n284));
  xnbna2aa1n03x5               g189(.a(new_n284), .b(new_n281), .c(new_n279), .out0(\s[27] ));
  norp02aa1n02x5               g190(.a(\b[27] ), .b(\a[28] ), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(\b[27] ), .b(\a[28] ), .o1(new_n287));
  norb02aa1n02x5               g192(.a(new_n287), .b(new_n286), .out0(new_n288));
  oai112aa1n03x5               g193(.a(new_n281), .b(new_n279), .c(\b[26] ), .d(\a[27] ), .o1(new_n289));
  aoi012aa1n03x5               g194(.a(new_n288), .b(new_n289), .c(new_n283), .o1(new_n290));
  aobi12aa1n06x5               g195(.a(new_n278), .b(new_n186), .c(new_n190), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n280), .b(new_n277), .c(new_n257), .d(new_n260), .o1(new_n292));
  nor043aa1n02x5               g197(.a(new_n292), .b(new_n291), .c(new_n282), .o1(new_n293));
  nano22aa1n03x7               g198(.a(new_n293), .b(new_n283), .c(new_n288), .out0(new_n294));
  nor002aa1n02x5               g199(.a(new_n290), .b(new_n294), .o1(\s[28] ));
  nano23aa1n02x4               g200(.a(new_n282), .b(new_n286), .c(new_n287), .d(new_n283), .out0(new_n296));
  oai012aa1n03x5               g201(.a(new_n296), .b(new_n292), .c(new_n291), .o1(new_n297));
  aoi012aa1n02x5               g202(.a(new_n286), .b(new_n282), .c(new_n287), .o1(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .out0(new_n299));
  tech160nm_fiaoi012aa1n05x5   g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n296), .b(new_n281), .c(new_n279), .out0(new_n301));
  nano22aa1n03x5               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g209(.a(new_n299), .b(new_n284), .c(new_n288), .out0(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(new_n292), .c(new_n291), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  aobi12aa1n02x7               g214(.a(new_n305), .b(new_n281), .c(new_n279), .out0(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n307), .c(new_n308), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[30] ));
  nano23aa1n02x4               g217(.a(new_n308), .b(new_n299), .c(new_n288), .d(new_n284), .out0(new_n313));
  oai012aa1n03x5               g218(.a(new_n313), .b(new_n292), .c(new_n291), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n314), .c(new_n315), .o1(new_n317));
  aobi12aa1n02x7               g222(.a(new_n313), .b(new_n281), .c(new_n279), .out0(new_n318));
  nano22aa1n03x5               g223(.a(new_n318), .b(new_n315), .c(new_n316), .out0(new_n319));
  norp02aa1n03x5               g224(.a(new_n317), .b(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g225(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g226(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g228(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g229(.a(\a[5] ), .b(\b[4] ), .c(new_n128), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norp02aa1n02x5               g231(.a(\b[5] ), .b(\a[6] ), .o1(new_n327));
  oai012aa1n02x5               g232(.a(new_n114), .b(new_n325), .c(new_n327), .o1(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g234(.a(\a[7] ), .b(\b[6] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g236(.a(new_n133), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


