// Benchmark "adder" written by ABC on Thu Jul 18 09:20:56 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n303, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n325, new_n326,
    new_n328, new_n329, new_n331, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n20x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor042aa1n04x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nand42aa1n03x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nor022aa1n16x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  tech160nm_fioai012aa1n03p5x5 g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  aoi022aa1d24x5               g010(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n106));
  nor042aa1n03x5               g011(.a(new_n106), .b(new_n105), .o1(new_n107));
  tech160nm_finand02aa1n03p5x5 g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nona23aa1n09x5               g013(.a(new_n101), .b(new_n108), .c(new_n103), .d(new_n102), .out0(new_n109));
  oaih12aa1n12x5               g014(.a(new_n104), .b(new_n109), .c(new_n107), .o1(new_n110));
  norp02aa1n12x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand22aa1n09x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1d18x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  xnrc02aa1n03x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nor043aa1n06x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[5] ), .o1(new_n119));
  oai022aa1n02x7               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  oaib12aa1n02x5               g025(.a(new_n120), .b(new_n119), .c(\a[6] ), .out0(new_n121));
  oai012aa1n02x5               g026(.a(new_n112), .b(new_n113), .c(new_n111), .o1(new_n122));
  oai012aa1n04x7               g027(.a(new_n122), .b(new_n115), .c(new_n121), .o1(new_n123));
  tech160nm_fiao0012aa1n02p5x5 g028(.a(new_n123), .b(new_n110), .c(new_n118), .o(new_n124));
  nand42aa1n06x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  aoai13aa1n02x5               g030(.a(new_n99), .b(new_n100), .c(new_n124), .d(new_n125), .o1(new_n126));
  inv000aa1n02x5               g031(.a(new_n98), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n125), .b(new_n100), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n123), .c(new_n110), .d(new_n118), .o1(new_n129));
  nona32aa1n02x4               g034(.a(new_n129), .b(new_n100), .c(new_n127), .d(new_n97), .out0(new_n130));
  nanp02aa1n02x5               g035(.a(new_n126), .b(new_n130), .o1(\s[10] ));
  nor042aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n06x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n06x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  inv000aa1d42x5               g039(.a(new_n134), .o1(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n130), .c(new_n98), .out0(\s[11] ));
  nor042aa1n02x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  tech160nm_finand02aa1n05x5   g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  aoi013aa1n02x4               g044(.a(new_n132), .b(new_n130), .c(new_n98), .d(new_n133), .o1(new_n140));
  xnrc02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(\s[12] ));
  nano32aa1n03x7               g046(.a(new_n99), .b(new_n139), .c(new_n128), .d(new_n134), .out0(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n123), .c(new_n110), .d(new_n118), .o1(new_n143));
  nano23aa1n03x7               g048(.a(new_n132), .b(new_n137), .c(new_n138), .d(new_n133), .out0(new_n144));
  oab012aa1n04x5               g049(.a(new_n127), .b(new_n97), .c(new_n100), .out0(new_n145));
  nanp02aa1n06x5               g050(.a(new_n144), .b(new_n145), .o1(new_n146));
  oai012aa1n02x7               g051(.a(new_n138), .b(new_n137), .c(new_n132), .o1(new_n147));
  nand02aa1d08x5               g052(.a(new_n146), .b(new_n147), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  norp02aa1n02x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nand42aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nanb02aa1n02x5               g056(.a(new_n150), .b(new_n151), .out0(new_n152));
  xobna2aa1n03x5               g057(.a(new_n152), .b(new_n143), .c(new_n149), .out0(\s[13] ));
  inv000aa1d42x5               g058(.a(\a[13] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(\b[12] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n143), .b(new_n149), .o1(new_n156));
  oaoi03aa1n03x5               g061(.a(new_n154), .b(new_n155), .c(new_n156), .o1(new_n157));
  xnrb03aa1n02x5               g062(.a(new_n157), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nanp02aa1n09x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(new_n161));
  nona22aa1n02x4               g066(.a(new_n156), .b(new_n152), .c(new_n161), .out0(new_n162));
  aoai13aa1n06x5               g067(.a(new_n160), .b(new_n159), .c(new_n154), .d(new_n155), .o1(new_n163));
  nor002aa1n16x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand02aa1n04x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n162), .c(new_n163), .out0(\s[15] ));
  inv000aa1d42x5               g072(.a(new_n164), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n161), .b(new_n152), .c(new_n143), .d(new_n149), .o1(new_n169));
  inv000aa1n02x5               g074(.a(new_n163), .o1(new_n170));
  oai012aa1n02x5               g075(.a(new_n166), .b(new_n169), .c(new_n170), .o1(new_n171));
  nor042aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand02aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  tech160nm_fiaoi012aa1n02p5x5 g079(.a(new_n174), .b(new_n171), .c(new_n168), .o1(new_n175));
  aobi12aa1n02x5               g080(.a(new_n166), .b(new_n162), .c(new_n163), .out0(new_n176));
  nano22aa1n02x4               g081(.a(new_n176), .b(new_n168), .c(new_n174), .out0(new_n177));
  norp02aa1n02x5               g082(.a(new_n175), .b(new_n177), .o1(\s[16] ));
  nano23aa1n02x5               g083(.a(new_n97), .b(new_n100), .c(new_n125), .d(new_n98), .out0(new_n179));
  nano23aa1n06x5               g084(.a(new_n164), .b(new_n172), .c(new_n173), .d(new_n165), .out0(new_n180));
  nano23aa1n03x5               g085(.a(new_n150), .b(new_n159), .c(new_n160), .d(new_n151), .out0(new_n181));
  nand02aa1n02x5               g086(.a(new_n181), .b(new_n180), .o1(new_n182));
  nano22aa1n03x7               g087(.a(new_n182), .b(new_n144), .c(new_n179), .out0(new_n183));
  aoai13aa1n12x5               g088(.a(new_n183), .b(new_n123), .c(new_n110), .d(new_n118), .o1(new_n184));
  inv030aa1n02x5               g089(.a(new_n182), .o1(new_n185));
  oai012aa1n02x5               g090(.a(new_n173), .b(new_n172), .c(new_n164), .o1(new_n186));
  aob012aa1n09x5               g091(.a(new_n186), .b(new_n180), .c(new_n170), .out0(new_n187));
  aoi012aa1d24x5               g092(.a(new_n187), .b(new_n148), .c(new_n185), .o1(new_n188));
  xorc02aa1n12x5               g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  xnbna2aa1n03x5               g094(.a(new_n189), .b(new_n184), .c(new_n188), .out0(\s[17] ));
  inv000aa1d42x5               g095(.a(\a[17] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[16] ), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(new_n192), .b(new_n191), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n189), .o1(new_n194));
  aoai13aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n184), .d(new_n188), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nand02aa1d10x5               g101(.a(new_n184), .b(new_n188), .o1(new_n197));
  nor022aa1n16x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nand02aa1n06x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  nona22aa1n03x5               g105(.a(new_n197), .b(new_n194), .c(new_n200), .out0(new_n201));
  aoai13aa1n12x5               g106(.a(new_n199), .b(new_n198), .c(new_n191), .d(new_n192), .o1(new_n202));
  nor022aa1n12x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand42aa1n08x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n201), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n03x5               g112(.a(new_n203), .o1(new_n208));
  aoi112aa1n03x5               g113(.a(new_n200), .b(new_n194), .c(new_n184), .d(new_n188), .o1(new_n209));
  inv000aa1n02x5               g114(.a(new_n202), .o1(new_n210));
  oai012aa1n03x5               g115(.a(new_n205), .b(new_n209), .c(new_n210), .o1(new_n211));
  nor022aa1n16x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand42aa1n06x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  tech160nm_fiaoi012aa1n05x5   g120(.a(new_n215), .b(new_n211), .c(new_n208), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n205), .o1(new_n217));
  tech160nm_fiaoi012aa1n05x5   g122(.a(new_n217), .b(new_n201), .c(new_n202), .o1(new_n218));
  nano22aa1n03x7               g123(.a(new_n218), .b(new_n208), .c(new_n215), .out0(new_n219));
  nor002aa1n02x5               g124(.a(new_n216), .b(new_n219), .o1(\s[20] ));
  nano23aa1n03x7               g125(.a(new_n203), .b(new_n212), .c(new_n213), .d(new_n204), .out0(new_n221));
  nanb03aa1n12x5               g126(.a(new_n200), .b(new_n221), .c(new_n189), .out0(new_n222));
  nona23aa1n09x5               g127(.a(new_n213), .b(new_n204), .c(new_n203), .d(new_n212), .out0(new_n223));
  oaoi03aa1n09x5               g128(.a(\a[20] ), .b(\b[19] ), .c(new_n208), .o1(new_n224));
  inv040aa1n02x5               g129(.a(new_n224), .o1(new_n225));
  oai012aa1n12x5               g130(.a(new_n225), .b(new_n223), .c(new_n202), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n222), .c(new_n184), .d(new_n188), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n233));
  aoi112aa1n02x7               g138(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n234));
  norb02aa1n03x4               g139(.a(new_n233), .b(new_n234), .out0(\s[22] ));
  inv030aa1d32x5               g140(.a(\a[21] ), .o1(new_n236));
  inv040aa1d32x5               g141(.a(\a[22] ), .o1(new_n237));
  xroi22aa1d06x4               g142(.a(new_n236), .b(\b[20] ), .c(new_n237), .d(\b[21] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n224), .c(new_n221), .d(new_n210), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\b[21] ), .o1(new_n240));
  oao003aa1n02x5               g145(.a(new_n237), .b(new_n240), .c(new_n230), .carry(new_n241));
  inv000aa1n02x5               g146(.a(new_n241), .o1(new_n242));
  nand22aa1n03x5               g147(.a(new_n239), .b(new_n242), .o1(new_n243));
  inv000aa1n02x5               g148(.a(new_n243), .o1(new_n244));
  inv000aa1n02x5               g149(.a(new_n238), .o1(new_n245));
  nona22aa1n06x5               g150(.a(new_n197), .b(new_n222), .c(new_n245), .out0(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[22] ), .b(\a[23] ), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  xnbna2aa1n03x5               g153(.a(new_n248), .b(new_n246), .c(new_n244), .out0(\s[23] ));
  orn002aa1n02x5               g154(.a(\a[23] ), .b(\b[22] ), .o(new_n250));
  tech160nm_fiaoi012aa1n05x5   g155(.a(new_n222), .b(new_n184), .c(new_n188), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n248), .b(new_n243), .c(new_n251), .d(new_n238), .o1(new_n252));
  tech160nm_fixnrc02aa1n04x5   g157(.a(\b[23] ), .b(\a[24] ), .out0(new_n253));
  tech160nm_fiaoi012aa1n02p5x5 g158(.a(new_n253), .b(new_n252), .c(new_n250), .o1(new_n254));
  tech160nm_fiaoi012aa1n02p5x5 g159(.a(new_n247), .b(new_n246), .c(new_n244), .o1(new_n255));
  nano22aa1n02x4               g160(.a(new_n255), .b(new_n250), .c(new_n253), .out0(new_n256));
  nor002aa1n02x5               g161(.a(new_n254), .b(new_n256), .o1(\s[24] ));
  nor042aa1n02x5               g162(.a(new_n253), .b(new_n247), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n258), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .c(new_n250), .carry(new_n260));
  aoai13aa1n04x5               g165(.a(new_n260), .b(new_n259), .c(new_n239), .d(new_n242), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  nona32aa1n06x5               g167(.a(new_n197), .b(new_n259), .c(new_n245), .d(new_n222), .out0(new_n263));
  xnrc02aa1n12x5               g168(.a(\b[24] ), .b(\a[25] ), .out0(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n263), .c(new_n262), .out0(\s[25] ));
  nor042aa1n03x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(new_n238), .b(new_n258), .o1(new_n269));
  aoi112aa1n02x5               g174(.a(new_n269), .b(new_n222), .c(new_n184), .d(new_n188), .o1(new_n270));
  oai012aa1n02x5               g175(.a(new_n265), .b(new_n270), .c(new_n261), .o1(new_n271));
  xnrc02aa1n02x5               g176(.a(\b[25] ), .b(\a[26] ), .out0(new_n272));
  aoi012aa1n02x7               g177(.a(new_n272), .b(new_n271), .c(new_n268), .o1(new_n273));
  aoi012aa1n06x5               g178(.a(new_n264), .b(new_n263), .c(new_n262), .o1(new_n274));
  nano22aa1n03x5               g179(.a(new_n274), .b(new_n268), .c(new_n272), .out0(new_n275));
  norp02aa1n03x5               g180(.a(new_n273), .b(new_n275), .o1(\s[26] ));
  xorc02aa1n12x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  nor002aa1n02x5               g182(.a(new_n272), .b(new_n264), .o1(new_n278));
  inv000aa1n02x5               g183(.a(new_n278), .o1(new_n279));
  nona32aa1d24x5               g184(.a(new_n197), .b(new_n279), .c(new_n269), .d(new_n222), .out0(new_n280));
  oao003aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .c(new_n268), .carry(new_n281));
  aobi12aa1n09x5               g186(.a(new_n281), .b(new_n261), .c(new_n278), .out0(new_n282));
  xnbna2aa1n06x5               g187(.a(new_n277), .b(new_n282), .c(new_n280), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  nano22aa1n06x5               g190(.a(new_n245), .b(new_n258), .c(new_n278), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n258), .b(new_n241), .c(new_n226), .d(new_n238), .o1(new_n287));
  aoai13aa1n04x5               g192(.a(new_n281), .b(new_n279), .c(new_n287), .d(new_n260), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n277), .b(new_n288), .c(new_n251), .d(new_n286), .o1(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[27] ), .b(\a[28] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n289), .c(new_n285), .o1(new_n291));
  aobi12aa1n06x5               g196(.a(new_n277), .b(new_n282), .c(new_n280), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n285), .c(new_n290), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[28] ));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  norb02aa1n02x5               g200(.a(new_n277), .b(new_n290), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n288), .c(new_n251), .d(new_n286), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n295), .b(new_n297), .c(new_n298), .o1(new_n299));
  aobi12aa1n06x5               g204(.a(new_n296), .b(new_n282), .c(new_n280), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n295), .c(new_n298), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[29] ));
  nanp02aa1n02x5               g207(.a(\b[0] ), .b(\a[1] ), .o1(new_n303));
  xorb03aa1n02x5               g208(.a(new_n303), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g209(.a(\b[29] ), .b(\a[30] ), .out0(new_n305));
  norb03aa1n02x5               g210(.a(new_n277), .b(new_n295), .c(new_n290), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n288), .c(new_n251), .d(new_n286), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n305), .b(new_n307), .c(new_n308), .o1(new_n309));
  aobi12aa1n06x5               g214(.a(new_n306), .b(new_n282), .c(new_n280), .out0(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n305), .c(new_n308), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[30] ));
  norb02aa1n02x5               g217(.a(new_n306), .b(new_n305), .out0(new_n313));
  aobi12aa1n06x5               g218(.a(new_n313), .b(new_n282), .c(new_n280), .out0(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  nano22aa1n03x5               g221(.a(new_n314), .b(new_n315), .c(new_n316), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n313), .b(new_n288), .c(new_n251), .d(new_n286), .o1(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n316), .b(new_n318), .c(new_n315), .o1(new_n319));
  norp02aa1n03x5               g224(.a(new_n319), .b(new_n317), .o1(\s[31] ));
  xnrb03aa1n02x5               g225(.a(new_n107), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi13aa1n02x5               g226(.a(new_n103), .b(new_n108), .c(new_n106), .d(new_n105), .o1(new_n322));
  xnrb03aa1n02x5               g227(.a(new_n322), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g228(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n06x5               g229(.a(new_n117), .b(new_n110), .out0(new_n325));
  tech160nm_fioai012aa1n03p5x5 g230(.a(new_n325), .b(\b[4] ), .c(\a[5] ), .o1(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n03x5               g232(.a(new_n116), .b(new_n326), .out0(new_n328));
  oaib12aa1n06x5               g233(.a(new_n328), .b(\a[6] ), .c(new_n119), .out0(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  orn002aa1n02x5               g235(.a(\a[8] ), .b(\b[7] ), .o(new_n331));
  tech160nm_fiaoi012aa1n05x5   g236(.a(new_n113), .b(new_n329), .c(new_n114), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n331), .c(new_n112), .out0(\s[8] ));
  xorb03aa1n02x5               g238(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


