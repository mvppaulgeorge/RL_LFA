// Benchmark "adder" written by ABC on Wed Jul 17 20:00:50 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n308, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n327, new_n329, new_n331, new_n332, new_n333,
    new_n335, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor002aa1n06x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai112aa1n06x5               g006(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n102));
  nand42aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  orn002aa1n06x5               g008(.a(\a[4] ), .b(\b[3] ), .o(new_n104));
  nand42aa1n02x5               g009(.a(new_n104), .b(new_n103), .o1(new_n105));
  aoi113aa1n03x7               g010(.a(new_n105), .b(new_n99), .c(new_n102), .d(new_n100), .e(new_n101), .o1(new_n106));
  nand42aa1n20x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand02aa1d08x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nano22aa1n06x5               g014(.a(new_n108), .b(new_n107), .c(new_n109), .out0(new_n110));
  xorc02aa1n02x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  nor002aa1d24x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nano23aa1n06x5               g019(.a(new_n113), .b(new_n112), .c(new_n114), .d(new_n103), .out0(new_n115));
  nand03aa1n02x5               g020(.a(new_n115), .b(new_n110), .c(new_n111), .o1(new_n116));
  inv000aa1d42x5               g021(.a(new_n112), .o1(new_n117));
  oai112aa1n02x5               g022(.a(new_n117), .b(new_n107), .c(\b[4] ), .d(\a[5] ), .o1(new_n118));
  inv040aa1d32x5               g023(.a(\a[8] ), .o1(new_n119));
  inv040aa1d28x5               g024(.a(\b[7] ), .o1(new_n120));
  oaoi03aa1n06x5               g025(.a(new_n119), .b(new_n120), .c(new_n108), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n121), .o1(new_n122));
  aoi013aa1n02x4               g027(.a(new_n122), .b(new_n110), .c(new_n118), .d(new_n111), .o1(new_n123));
  tech160nm_fioai012aa1n05x5   g028(.a(new_n123), .b(new_n116), .c(new_n106), .o1(new_n124));
  nand42aa1n16x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nanp03aa1n03x5               g030(.a(new_n124), .b(new_n98), .c(new_n125), .o1(new_n126));
  nor002aa1n16x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n20x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  norb03aa1d15x5               g035(.a(new_n128), .b(new_n97), .c(new_n127), .out0(new_n131));
  aoi022aa1n02x7               g036(.a(new_n126), .b(new_n131), .c(\b[9] ), .d(\a[10] ), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nand42aa1d28x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor002aa1d32x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1d16x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanb02aa1n12x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  aoai13aa1n03x5               g043(.a(new_n138), .b(new_n135), .c(new_n132), .d(new_n134), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n126), .b(new_n131), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n134), .b(new_n135), .out0(new_n141));
  nanp03aa1n02x5               g046(.a(new_n140), .b(new_n128), .c(new_n141), .o1(new_n142));
  nona22aa1n02x4               g047(.a(new_n142), .b(new_n138), .c(new_n135), .out0(new_n143));
  nanp02aa1n02x5               g048(.a(new_n139), .b(new_n143), .o1(\s[12] ));
  nanb02aa1n06x5               g049(.a(new_n99), .b(new_n100), .out0(new_n145));
  nanp02aa1n09x5               g050(.a(new_n102), .b(new_n101), .o1(new_n146));
  nano22aa1n03x7               g051(.a(new_n99), .b(new_n104), .c(new_n103), .out0(new_n147));
  oai012aa1n12x5               g052(.a(new_n147), .b(new_n146), .c(new_n145), .o1(new_n148));
  nanb03aa1d18x5               g053(.a(new_n108), .b(new_n109), .c(new_n107), .out0(new_n149));
  nanp02aa1n03x5               g054(.a(\b[7] ), .b(\a[8] ), .o1(new_n150));
  nand02aa1n03x5               g055(.a(new_n120), .b(new_n119), .o1(new_n151));
  nand02aa1n03x5               g056(.a(new_n151), .b(new_n150), .o1(new_n152));
  nona23aa1n09x5               g057(.a(new_n103), .b(new_n114), .c(new_n113), .d(new_n112), .out0(new_n153));
  nor043aa1n06x5               g058(.a(new_n153), .b(new_n152), .c(new_n149), .o1(new_n154));
  norb03aa1n03x5               g059(.a(new_n107), .b(new_n113), .c(new_n112), .out0(new_n155));
  oai013aa1n06x5               g060(.a(new_n121), .b(new_n155), .c(new_n149), .d(new_n152), .o1(new_n156));
  norb02aa1n15x5               g061(.a(new_n137), .b(new_n136), .out0(new_n157));
  nano22aa1d15x5               g062(.a(new_n135), .b(new_n128), .c(new_n134), .out0(new_n158));
  norb03aa1d15x5               g063(.a(new_n125), .b(new_n97), .c(new_n127), .out0(new_n159));
  nand23aa1d12x5               g064(.a(new_n158), .b(new_n159), .c(new_n157), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n06x5               g066(.a(new_n161), .b(new_n156), .c(new_n154), .d(new_n148), .o1(new_n162));
  nanb03aa1d24x5               g067(.a(new_n135), .b(new_n128), .c(new_n134), .out0(new_n163));
  aoi012aa1d24x5               g068(.a(new_n136), .b(new_n135), .c(new_n137), .o1(new_n164));
  oai013aa1d12x5               g069(.a(new_n164), .b(new_n131), .c(new_n163), .d(new_n138), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(new_n162), .b(new_n166), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d24x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nanp02aa1n04x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n169), .b(new_n167), .c(new_n170), .o1(new_n171));
  xnrb03aa1n02x5               g076(.a(new_n171), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nand22aa1n12x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nona23aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n169), .d(new_n173), .out0(new_n175));
  aoi012aa1d24x5               g080(.a(new_n173), .b(new_n169), .c(new_n174), .o1(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n175), .c(new_n162), .d(new_n166), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nanp02aa1n12x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  norb02aa1n12x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  nor042aa1n09x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand42aa1n06x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nanb02aa1n06x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n179), .c(new_n177), .d(new_n181), .o1(new_n185));
  aoi112aa1n02x5               g090(.a(new_n179), .b(new_n184), .c(new_n177), .d(new_n180), .o1(new_n186));
  nanb02aa1n02x5               g091(.a(new_n186), .b(new_n185), .out0(\s[16] ));
  nano23aa1n06x5               g092(.a(new_n169), .b(new_n173), .c(new_n174), .d(new_n170), .out0(new_n188));
  nano23aa1n06x5               g093(.a(new_n179), .b(new_n182), .c(new_n183), .d(new_n180), .out0(new_n189));
  nano22aa1d15x5               g094(.a(new_n160), .b(new_n188), .c(new_n189), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n156), .c(new_n154), .d(new_n148), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n181), .o1(new_n192));
  nor043aa1n06x5               g097(.a(new_n175), .b(new_n192), .c(new_n184), .o1(new_n193));
  tech160nm_fioai012aa1n04x5   g098(.a(new_n183), .b(new_n182), .c(new_n179), .o1(new_n194));
  oai013aa1n06x5               g099(.a(new_n194), .b(new_n192), .c(new_n176), .d(new_n184), .o1(new_n195));
  aoi012aa1d24x5               g100(.a(new_n195), .b(new_n165), .c(new_n193), .o1(new_n196));
  xnrc02aa1n12x5               g101(.a(\b[16] ), .b(\a[17] ), .out0(new_n197));
  xobna2aa1n03x5               g102(.a(new_n197), .b(new_n191), .c(new_n196), .out0(\s[17] ));
  orn002aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .o(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n197), .c(new_n191), .d(new_n196), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  tech160nm_fixnrc02aa1n02p5x5 g106(.a(\b[17] ), .b(\a[18] ), .out0(new_n202));
  nor042aa1n06x5               g107(.a(new_n202), .b(new_n197), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  nor042aa1n02x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  aoi112aa1n09x5               g110(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n206));
  norp02aa1n02x5               g111(.a(new_n206), .b(new_n205), .o1(new_n207));
  aoai13aa1n04x5               g112(.a(new_n207), .b(new_n204), .c(new_n191), .d(new_n196), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand02aa1n06x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nor042aa1d18x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d28x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1d27x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n211), .c(new_n208), .d(new_n212), .o1(new_n217));
  aoi112aa1n03x5               g122(.a(new_n211), .b(new_n216), .c(new_n208), .d(new_n212), .o1(new_n218));
  nanb02aa1n03x5               g123(.a(new_n218), .b(new_n217), .out0(\s[20] ));
  nano23aa1n02x5               g124(.a(new_n211), .b(new_n213), .c(new_n214), .d(new_n212), .out0(new_n220));
  nona22aa1n02x4               g125(.a(new_n220), .b(new_n202), .c(new_n197), .out0(new_n221));
  norb02aa1n03x5               g126(.a(new_n212), .b(new_n211), .out0(new_n222));
  oai112aa1n06x5               g127(.a(new_n222), .b(new_n215), .c(new_n206), .d(new_n205), .o1(new_n223));
  aoi012aa1n12x5               g128(.a(new_n213), .b(new_n211), .c(new_n214), .o1(new_n224));
  nand22aa1n12x5               g129(.a(new_n223), .b(new_n224), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n221), .c(new_n191), .d(new_n196), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n229), .c(new_n227), .d(new_n231), .o1(new_n233));
  aoi112aa1n03x4               g138(.a(new_n229), .b(new_n232), .c(new_n227), .d(new_n231), .o1(new_n234));
  nanb02aa1n03x5               g139(.a(new_n234), .b(new_n233), .out0(\s[22] ));
  nor042aa1n04x5               g140(.a(new_n232), .b(new_n230), .o1(new_n236));
  nand23aa1n03x5               g141(.a(new_n236), .b(new_n203), .c(new_n220), .o1(new_n237));
  norp02aa1n02x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nanp02aa1n02x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n238), .b(new_n229), .c(new_n239), .o1(new_n240));
  aobi12aa1n02x7               g145(.a(new_n240), .b(new_n225), .c(new_n236), .out0(new_n241));
  aoai13aa1n04x5               g146(.a(new_n241), .b(new_n237), .c(new_n191), .d(new_n196), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n04x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  nanp02aa1n04x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  nor042aa1d18x5               g150(.a(\b[23] ), .b(\a[24] ), .o1(new_n246));
  nanp02aa1n04x5               g151(.a(\b[23] ), .b(\a[24] ), .o1(new_n247));
  nanb02aa1n02x5               g152(.a(new_n246), .b(new_n247), .out0(new_n248));
  aoai13aa1n03x5               g153(.a(new_n248), .b(new_n244), .c(new_n242), .d(new_n245), .o1(new_n249));
  aoi112aa1n03x5               g154(.a(new_n244), .b(new_n248), .c(new_n242), .d(new_n245), .o1(new_n250));
  nanb02aa1n03x5               g155(.a(new_n250), .b(new_n249), .out0(\s[24] ));
  nona23aa1n09x5               g156(.a(new_n247), .b(new_n245), .c(new_n244), .d(new_n246), .out0(new_n252));
  inv030aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  nanb03aa1n02x5               g158(.a(new_n221), .b(new_n253), .c(new_n236), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n246), .o1(new_n255));
  nanp02aa1n02x5               g160(.a(new_n244), .b(new_n247), .o1(new_n256));
  oai112aa1n03x5               g161(.a(new_n256), .b(new_n255), .c(new_n252), .d(new_n240), .o1(new_n257));
  aoi013aa1n03x5               g162(.a(new_n257), .b(new_n225), .c(new_n236), .d(new_n253), .o1(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n254), .c(new_n191), .d(new_n196), .o1(new_n259));
  xorb03aa1n02x5               g164(.a(new_n259), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  xorc02aa1n12x5               g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[25] ), .b(\a[26] ), .out0(new_n263));
  aoai13aa1n03x5               g168(.a(new_n263), .b(new_n261), .c(new_n259), .d(new_n262), .o1(new_n264));
  aoi112aa1n03x5               g169(.a(new_n261), .b(new_n263), .c(new_n259), .d(new_n262), .o1(new_n265));
  nanb02aa1n03x5               g170(.a(new_n265), .b(new_n264), .out0(\s[26] ));
  nona22aa1n02x4               g171(.a(new_n128), .b(new_n127), .c(new_n97), .out0(new_n267));
  nanp03aa1n02x5               g172(.a(new_n267), .b(new_n158), .c(new_n157), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(new_n189), .b(new_n188), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n176), .o1(new_n270));
  aobi12aa1n02x7               g175(.a(new_n194), .b(new_n189), .c(new_n270), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n269), .c(new_n268), .d(new_n164), .o1(new_n272));
  norb02aa1n09x5               g177(.a(new_n262), .b(new_n263), .out0(new_n273));
  nano22aa1n03x7               g178(.a(new_n237), .b(new_n253), .c(new_n273), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n272), .c(new_n124), .d(new_n190), .o1(new_n275));
  inv040aa1n03x5               g180(.a(new_n236), .o1(new_n276));
  aoi112aa1n03x5               g181(.a(new_n276), .b(new_n252), .c(new_n223), .d(new_n224), .o1(new_n277));
  inv000aa1d42x5               g182(.a(\a[26] ), .o1(new_n278));
  inv000aa1d42x5               g183(.a(\b[25] ), .o1(new_n279));
  oao003aa1n02x5               g184(.a(new_n278), .b(new_n279), .c(new_n261), .carry(new_n280));
  oaoi13aa1n09x5               g185(.a(new_n280), .b(new_n273), .c(new_n277), .d(new_n257), .o1(new_n281));
  xorc02aa1n02x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n275), .out0(\s[27] ));
  nand42aa1n03x5               g188(.a(new_n281), .b(new_n275), .o1(new_n284));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  tech160nm_fixorc02aa1n03p5x5 g190(.a(\a[28] ), .b(\b[27] ), .out0(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n285), .c(new_n284), .d(new_n282), .o1(new_n288));
  nanp02aa1n06x5               g193(.a(new_n191), .b(new_n196), .o1(new_n289));
  nona32aa1n03x5               g194(.a(new_n225), .b(new_n252), .c(new_n232), .d(new_n230), .out0(new_n290));
  norp02aa1n02x5               g195(.a(new_n252), .b(new_n240), .o1(new_n291));
  nano22aa1n02x4               g196(.a(new_n291), .b(new_n255), .c(new_n256), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n273), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n280), .o1(new_n294));
  aoai13aa1n06x5               g199(.a(new_n294), .b(new_n293), .c(new_n290), .d(new_n292), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n282), .b(new_n295), .c(new_n289), .d(new_n274), .o1(new_n296));
  nona22aa1n02x5               g201(.a(new_n296), .b(new_n287), .c(new_n285), .out0(new_n297));
  nanp02aa1n03x5               g202(.a(new_n288), .b(new_n297), .o1(\s[28] ));
  and002aa1n02x5               g203(.a(new_n286), .b(new_n282), .o(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n295), .c(new_n289), .d(new_n274), .o1(new_n300));
  aoi112aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n301));
  oab012aa1n02x4               g206(.a(new_n301), .b(\a[28] ), .c(\b[27] ), .out0(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[28] ), .b(\a[29] ), .out0(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n300), .c(new_n302), .o1(new_n304));
  aobi12aa1n02x7               g209(.a(new_n299), .b(new_n281), .c(new_n275), .out0(new_n305));
  nano22aa1n03x5               g210(.a(new_n305), .b(new_n302), .c(new_n303), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n304), .b(new_n306), .o1(\s[29] ));
  nanp02aa1n02x5               g212(.a(\b[0] ), .b(\a[1] ), .o1(new_n308));
  xorb03aa1n02x5               g213(.a(new_n308), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g214(.a(new_n303), .b(new_n282), .c(new_n286), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n295), .c(new_n289), .d(new_n274), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n302), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[29] ), .b(\a[30] ), .out0(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n313), .b(new_n311), .c(new_n312), .o1(new_n314));
  aobi12aa1n02x7               g219(.a(new_n310), .b(new_n281), .c(new_n275), .out0(new_n315));
  nano22aa1n03x5               g220(.a(new_n315), .b(new_n312), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[30] ));
  nano23aa1n02x4               g222(.a(new_n313), .b(new_n303), .c(new_n286), .d(new_n282), .out0(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n295), .c(new_n289), .d(new_n274), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n320));
  xnrc02aa1n02x5               g225(.a(\b[30] ), .b(\a[31] ), .out0(new_n321));
  tech160nm_fiaoi012aa1n02p5x5 g226(.a(new_n321), .b(new_n319), .c(new_n320), .o1(new_n322));
  aobi12aa1n02x7               g227(.a(new_n318), .b(new_n281), .c(new_n275), .out0(new_n323));
  nano22aa1n03x5               g228(.a(new_n323), .b(new_n320), .c(new_n321), .out0(new_n324));
  norp02aa1n03x5               g229(.a(new_n322), .b(new_n324), .o1(\s[31] ));
  xnbna2aa1n03x5               g230(.a(new_n145), .b(new_n102), .c(new_n101), .out0(\s[3] ));
  aoi013aa1n02x4               g231(.a(new_n99), .b(new_n102), .c(new_n101), .d(new_n100), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n148), .b(new_n327), .c(new_n105), .out0(\s[4] ));
  nanb02aa1n02x5               g233(.a(new_n113), .b(new_n114), .out0(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n329), .b(new_n148), .c(new_n103), .out0(\s[5] ));
  aoi013aa1n02x4               g235(.a(new_n113), .b(new_n148), .c(new_n103), .d(new_n114), .o1(new_n331));
  nanb03aa1n02x5               g236(.a(new_n113), .b(new_n114), .c(new_n103), .out0(new_n332));
  oai012aa1n02x5               g237(.a(new_n155), .b(new_n106), .c(new_n332), .o1(new_n333));
  aoai13aa1n02x5               g238(.a(new_n333), .b(new_n331), .c(new_n107), .d(new_n117), .o1(\s[6] ));
  norb02aa1n02x5               g239(.a(new_n109), .b(new_n108), .out0(new_n335));
  xobna2aa1n03x5               g240(.a(new_n335), .b(new_n333), .c(new_n107), .out0(\s[7] ));
  aoi012aa1n02x5               g241(.a(new_n108), .b(new_n333), .c(new_n110), .o1(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n337), .b(new_n150), .c(new_n151), .out0(\s[8] ));
  xorb03aa1n02x5               g243(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


