// Benchmark "adder" written by ABC on Thu Jul 18 11:43:45 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n337,
    new_n338, new_n340, new_n343, new_n344, new_n346, new_n347, new_n349,
    new_n351;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1n08x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1n20x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nanb03aa1d18x5               g006(.a(new_n100), .b(new_n101), .c(new_n99), .out0(new_n102));
  nand02aa1d04x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  norp02aa1n04x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  norb03aa1n09x5               g009(.a(new_n101), .b(new_n104), .c(new_n103), .out0(new_n105));
  xnrc02aa1n12x5               g010(.a(\b[3] ), .b(\a[4] ), .out0(new_n106));
  inv030aa1n04x5               g011(.a(new_n100), .o1(new_n107));
  oao003aa1n12x5               g012(.a(\a[4] ), .b(\b[3] ), .c(new_n107), .carry(new_n108));
  oai013aa1d12x5               g013(.a(new_n108), .b(new_n105), .c(new_n102), .d(new_n106), .o1(new_n109));
  xorc02aa1n02x5               g014(.a(\a[6] ), .b(\b[5] ), .out0(new_n110));
  tech160nm_fixorc02aa1n05x5   g015(.a(\a[5] ), .b(\b[4] ), .out0(new_n111));
  xorc02aa1n12x5               g016(.a(\a[8] ), .b(\b[7] ), .out0(new_n112));
  nor042aa1n09x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  norb02aa1n09x5               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  nand42aa1n02x5               g020(.a(new_n112), .b(new_n115), .o1(new_n116));
  nano22aa1n03x7               g021(.a(new_n116), .b(new_n110), .c(new_n111), .out0(new_n117));
  nand42aa1n03x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nano22aa1n03x7               g023(.a(new_n113), .b(new_n118), .c(new_n114), .out0(new_n119));
  oai022aa1n12x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  nand43aa1n03x5               g025(.a(new_n119), .b(new_n112), .c(new_n120), .o1(new_n121));
  inv040aa1n02x5               g026(.a(new_n113), .o1(new_n122));
  oaoi03aa1n03x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  nanb02aa1n12x5               g028(.a(new_n123), .b(new_n121), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n03x5               g030(.a(new_n125), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n126));
  nor022aa1n16x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand02aa1d28x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n06x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  nona22aa1n09x5               g035(.a(new_n101), .b(new_n104), .c(new_n103), .out0(new_n131));
  nona22aa1n09x5               g036(.a(new_n131), .b(new_n102), .c(new_n106), .out0(new_n132));
  tech160nm_fixnrc02aa1n05x5   g037(.a(\b[5] ), .b(\a[6] ), .out0(new_n133));
  tech160nm_fixnrc02aa1n05x5   g038(.a(\b[4] ), .b(\a[5] ), .out0(new_n134));
  nona23aa1n03x5               g039(.a(new_n112), .b(new_n115), .c(new_n134), .d(new_n133), .out0(new_n135));
  aoi013aa1n06x4               g040(.a(new_n123), .b(new_n119), .c(new_n112), .d(new_n120), .o1(new_n136));
  aoai13aa1n12x5               g041(.a(new_n136), .b(new_n135), .c(new_n132), .d(new_n108), .o1(new_n137));
  aoai13aa1n03x5               g042(.a(new_n129), .b(new_n97), .c(new_n137), .d(new_n125), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n128), .o1(new_n139));
  oai022aa1n02x5               g044(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n140));
  oaib12aa1n06x5               g045(.a(new_n138), .b(new_n139), .c(new_n140), .out0(new_n141));
  nor042aa1n12x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand42aa1n20x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  aboi22aa1n03x5               g049(.a(new_n142), .b(new_n143), .c(new_n140), .d(new_n128), .out0(new_n145));
  aoi022aa1n02x5               g050(.a(new_n141), .b(new_n144), .c(new_n138), .d(new_n145), .o1(\s[11] ));
  nor002aa1n06x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand22aa1n09x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n03x5               g055(.a(new_n150), .b(new_n142), .c(new_n141), .d(new_n143), .o1(new_n151));
  aobi12aa1n03x5               g056(.a(new_n129), .b(new_n126), .c(new_n98), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n144), .b(new_n152), .c(new_n128), .d(new_n140), .o1(new_n153));
  nona22aa1n02x5               g058(.a(new_n153), .b(new_n150), .c(new_n142), .out0(new_n154));
  nanp02aa1n03x5               g059(.a(new_n151), .b(new_n154), .o1(\s[12] ));
  nano23aa1n06x5               g060(.a(new_n142), .b(new_n147), .c(new_n148), .d(new_n143), .out0(new_n156));
  nand23aa1d12x5               g061(.a(new_n156), .b(new_n125), .c(new_n129), .o1(new_n157));
  inv000aa1n02x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n159));
  nano22aa1n03x5               g064(.a(new_n147), .b(new_n143), .c(new_n148), .out0(new_n160));
  tech160nm_fioai012aa1n03p5x5 g065(.a(new_n128), .b(\b[10] ), .c(\a[11] ), .o1(new_n161));
  oab012aa1n06x5               g066(.a(new_n161), .b(new_n97), .c(new_n127), .out0(new_n162));
  nanp02aa1n02x5               g067(.a(new_n162), .b(new_n160), .o1(new_n163));
  tech160nm_fiaoi012aa1n02p5x5 g068(.a(new_n147), .b(new_n142), .c(new_n148), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(new_n163), .b(new_n164), .o1(new_n165));
  inv000aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  nor042aa1n09x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  nand42aa1d28x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n159), .c(new_n166), .out0(\s[13] ));
  nanp02aa1n02x5               g075(.a(new_n159), .b(new_n166), .o1(new_n171));
  aoi012aa1n02x5               g076(.a(new_n167), .b(new_n171), .c(new_n168), .o1(new_n172));
  xnrb03aa1n02x5               g077(.a(new_n172), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nand42aa1d28x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nano23aa1d15x5               g080(.a(new_n167), .b(new_n174), .c(new_n175), .d(new_n168), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  oai012aa1n18x5               g082(.a(new_n175), .b(new_n174), .c(new_n167), .o1(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n177), .c(new_n159), .d(new_n166), .o1(new_n179));
  xnrc02aa1n12x5               g084(.a(\b[14] ), .b(\a[15] ), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n178), .o1(new_n182));
  aoi112aa1n02x5               g087(.a(new_n181), .b(new_n182), .c(new_n171), .d(new_n176), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n183), .b(new_n179), .c(new_n181), .o1(\s[15] ));
  norp02aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  tech160nm_fixnrc02aa1n04x5   g090(.a(\b[15] ), .b(\a[16] ), .out0(new_n186));
  aoai13aa1n02x5               g091(.a(new_n186), .b(new_n185), .c(new_n179), .d(new_n181), .o1(new_n187));
  aoi112aa1n03x4               g092(.a(new_n185), .b(new_n186), .c(new_n179), .d(new_n181), .o1(new_n188));
  nanb02aa1n03x5               g093(.a(new_n188), .b(new_n187), .out0(\s[16] ));
  nor042aa1n06x5               g094(.a(new_n186), .b(new_n180), .o1(new_n190));
  nano22aa1d15x5               g095(.a(new_n157), .b(new_n190), .c(new_n176), .out0(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n192));
  inv020aa1n03x5               g097(.a(new_n164), .o1(new_n193));
  aoai13aa1n06x5               g098(.a(new_n176), .b(new_n193), .c(new_n162), .d(new_n160), .o1(new_n194));
  nand42aa1n02x5               g099(.a(new_n194), .b(new_n178), .o1(new_n195));
  nanp02aa1n03x5               g100(.a(new_n195), .b(new_n190), .o1(new_n196));
  orn002aa1n02x5               g101(.a(\a[15] ), .b(\b[14] ), .o(new_n197));
  oao003aa1n02x5               g102(.a(\a[16] ), .b(\b[15] ), .c(new_n197), .carry(new_n198));
  nand23aa1n06x5               g103(.a(new_n192), .b(new_n196), .c(new_n198), .o1(new_n199));
  nor002aa1d32x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  nand42aa1d28x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  nano22aa1n02x4               g107(.a(new_n202), .b(new_n196), .c(new_n198), .out0(new_n203));
  aoi022aa1n02x5               g108(.a(new_n203), .b(new_n192), .c(new_n199), .d(new_n202), .o1(\s[17] ));
  tech160nm_fiaoi012aa1n05x5   g109(.a(new_n200), .b(new_n199), .c(new_n202), .o1(new_n205));
  xnrb03aa1n03x5               g110(.a(new_n205), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv030aa1n02x5               g111(.a(new_n190), .o1(new_n207));
  aoai13aa1n04x5               g112(.a(new_n198), .b(new_n207), .c(new_n194), .d(new_n178), .o1(new_n208));
  nor002aa1d32x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nano23aa1d15x5               g115(.a(new_n200), .b(new_n209), .c(new_n210), .d(new_n201), .out0(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n208), .c(new_n137), .d(new_n191), .o1(new_n212));
  oa0012aa1n02x5               g117(.a(new_n210), .b(new_n209), .c(new_n200), .o(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nor042aa1d18x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand02aa1n10x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n06x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g124(.a(new_n212), .b(new_n214), .o1(new_n220));
  nor002aa1d32x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1d28x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanb02aa1n06x5               g127(.a(new_n221), .b(new_n222), .out0(new_n223));
  aoai13aa1n02x5               g128(.a(new_n223), .b(new_n215), .c(new_n220), .d(new_n216), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n217), .b(new_n213), .c(new_n199), .d(new_n211), .o1(new_n225));
  nona22aa1n03x5               g130(.a(new_n225), .b(new_n223), .c(new_n215), .out0(new_n226));
  nanp02aa1n03x5               g131(.a(new_n224), .b(new_n226), .o1(\s[20] ));
  nanb03aa1n09x5               g132(.a(new_n221), .b(new_n222), .c(new_n216), .out0(new_n228));
  oai122aa1n12x5               g133(.a(new_n210), .b(new_n209), .c(new_n200), .d(\b[18] ), .e(\a[19] ), .o1(new_n229));
  aoi012aa1n12x5               g134(.a(new_n221), .b(new_n215), .c(new_n222), .o1(new_n230));
  oai012aa1n18x5               g135(.a(new_n230), .b(new_n229), .c(new_n228), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aobi12aa1n02x5               g137(.a(new_n198), .b(new_n195), .c(new_n190), .out0(new_n233));
  nanb03aa1d18x5               g138(.a(new_n223), .b(new_n211), .c(new_n217), .out0(new_n234));
  aoai13aa1n02x7               g139(.a(new_n232), .b(new_n234), .c(new_n233), .d(new_n192), .o1(new_n235));
  nor002aa1d32x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nand42aa1d28x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n234), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n238), .b(new_n199), .c(new_n239), .o1(new_n240));
  aoi022aa1n02x5               g145(.a(new_n240), .b(new_n232), .c(new_n235), .d(new_n238), .o1(\s[21] ));
  nor002aa1d32x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  nand42aa1d28x5               g147(.a(\b[21] ), .b(\a[22] ), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n236), .c(new_n235), .d(new_n238), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n238), .b(new_n231), .c(new_n199), .d(new_n239), .o1(new_n246));
  nona22aa1n03x5               g151(.a(new_n246), .b(new_n244), .c(new_n236), .out0(new_n247));
  nanp02aa1n03x5               g152(.a(new_n245), .b(new_n247), .o1(\s[22] ));
  nano23aa1d15x5               g153(.a(new_n236), .b(new_n242), .c(new_n243), .d(new_n237), .out0(new_n249));
  nano32aa1n02x4               g154(.a(new_n223), .b(new_n249), .c(new_n211), .d(new_n217), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n208), .c(new_n137), .d(new_n191), .o1(new_n251));
  oa0012aa1n12x5               g156(.a(new_n243), .b(new_n242), .c(new_n236), .o(new_n252));
  aoi012aa1n02x5               g157(.a(new_n252), .b(new_n231), .c(new_n249), .o1(new_n253));
  nand02aa1n03x5               g158(.a(new_n251), .b(new_n253), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aoi112aa1n02x5               g160(.a(new_n255), .b(new_n252), .c(new_n231), .d(new_n249), .o1(new_n256));
  aoi022aa1n02x5               g161(.a(new_n254), .b(new_n255), .c(new_n251), .d(new_n256), .o1(\s[23] ));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[23] ), .b(\a[24] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n258), .c(new_n254), .d(new_n255), .o1(new_n260));
  inv000aa1n02x5               g165(.a(new_n253), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n255), .b(new_n261), .c(new_n199), .d(new_n250), .o1(new_n262));
  nona22aa1n03x5               g167(.a(new_n262), .b(new_n259), .c(new_n258), .out0(new_n263));
  nanp02aa1n03x5               g168(.a(new_n260), .b(new_n263), .o1(\s[24] ));
  norb02aa1n06x4               g169(.a(new_n255), .b(new_n259), .out0(new_n265));
  nano22aa1n03x7               g170(.a(new_n234), .b(new_n265), .c(new_n249), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n208), .c(new_n137), .d(new_n191), .o1(new_n267));
  nano22aa1n03x7               g172(.a(new_n221), .b(new_n216), .c(new_n222), .out0(new_n268));
  tech160nm_fioai012aa1n03p5x5 g173(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .o1(new_n269));
  oab012aa1n06x5               g174(.a(new_n269), .b(new_n200), .c(new_n209), .out0(new_n270));
  inv020aa1n03x5               g175(.a(new_n230), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n249), .b(new_n271), .c(new_n270), .d(new_n268), .o1(new_n272));
  inv030aa1n02x5               g177(.a(new_n252), .o1(new_n273));
  inv020aa1n04x5               g178(.a(new_n265), .o1(new_n274));
  oai022aa1n02x5               g179(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n275));
  aob012aa1n02x5               g180(.a(new_n275), .b(\b[23] ), .c(\a[24] ), .out0(new_n276));
  aoai13aa1n12x5               g181(.a(new_n276), .b(new_n274), .c(new_n272), .d(new_n273), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  tech160nm_finand02aa1n03p5x5 g183(.a(new_n267), .b(new_n278), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[25] ), .b(\b[24] ), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n265), .b(new_n252), .c(new_n231), .d(new_n249), .o1(new_n281));
  nano22aa1n02x4               g186(.a(new_n280), .b(new_n281), .c(new_n276), .out0(new_n282));
  aoi022aa1n02x5               g187(.a(new_n279), .b(new_n280), .c(new_n267), .d(new_n282), .o1(\s[25] ));
  norp02aa1n02x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  tech160nm_fixnrc02aa1n05x5   g189(.a(\b[25] ), .b(\a[26] ), .out0(new_n285));
  aoai13aa1n02x7               g190(.a(new_n285), .b(new_n284), .c(new_n279), .d(new_n280), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n280), .b(new_n277), .c(new_n199), .d(new_n266), .o1(new_n287));
  nona22aa1n03x5               g192(.a(new_n287), .b(new_n285), .c(new_n284), .out0(new_n288));
  nanp02aa1n03x5               g193(.a(new_n286), .b(new_n288), .o1(\s[26] ));
  norb02aa1n12x5               g194(.a(new_n280), .b(new_n285), .out0(new_n290));
  inv000aa1n02x5               g195(.a(new_n290), .o1(new_n291));
  nano23aa1d12x5               g196(.a(new_n291), .b(new_n234), .c(new_n265), .d(new_n249), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n208), .c(new_n137), .d(new_n191), .o1(new_n293));
  nanp02aa1n02x5               g198(.a(\b[25] ), .b(\a[26] ), .o1(new_n294));
  oai022aa1n02x5               g199(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n295));
  nanp02aa1n02x5               g200(.a(new_n295), .b(new_n294), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n296), .b(new_n291), .c(new_n281), .d(new_n276), .o1(new_n297));
  xorc02aa1n12x5               g202(.a(\a[27] ), .b(\b[26] ), .out0(new_n298));
  aoai13aa1n06x5               g203(.a(new_n298), .b(new_n297), .c(new_n199), .d(new_n292), .o1(new_n299));
  aoi122aa1n02x5               g204(.a(new_n298), .b(new_n294), .c(new_n295), .d(new_n277), .e(new_n290), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n299), .b(new_n300), .c(new_n293), .out0(\s[27] ));
  xnrc02aa1n02x5               g206(.a(\b[27] ), .b(\a[28] ), .out0(new_n302));
  aoi022aa1n12x5               g207(.a(new_n277), .b(new_n290), .c(new_n294), .d(new_n295), .o1(new_n303));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  inv000aa1n03x5               g209(.a(new_n304), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n298), .o1(new_n306));
  aoai13aa1n06x5               g211(.a(new_n305), .b(new_n306), .c(new_n293), .d(new_n303), .o1(new_n307));
  nanp02aa1n03x5               g212(.a(new_n307), .b(new_n302), .o1(new_n308));
  nona22aa1n02x5               g213(.a(new_n299), .b(new_n302), .c(new_n304), .out0(new_n309));
  nanp02aa1n03x5               g214(.a(new_n308), .b(new_n309), .o1(\s[28] ));
  norb02aa1n06x5               g215(.a(new_n298), .b(new_n302), .out0(new_n311));
  aoai13aa1n02x5               g216(.a(new_n311), .b(new_n297), .c(new_n199), .d(new_n292), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  oao003aa1n02x5               g218(.a(\a[28] ), .b(\b[27] ), .c(new_n305), .carry(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n313), .c(new_n293), .d(new_n303), .o1(new_n315));
  tech160nm_fixorc02aa1n02p5x5 g220(.a(\a[29] ), .b(\b[28] ), .out0(new_n316));
  norb02aa1n02x5               g221(.a(new_n314), .b(new_n316), .out0(new_n317));
  aoi022aa1n03x5               g222(.a(new_n315), .b(new_n316), .c(new_n312), .d(new_n317), .o1(\s[29] ));
  xorb03aa1n02x5               g223(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g224(.a(new_n302), .b(new_n298), .c(new_n316), .out0(new_n320));
  aoai13aa1n02x5               g225(.a(new_n320), .b(new_n297), .c(new_n199), .d(new_n292), .o1(new_n321));
  inv000aa1n02x5               g226(.a(new_n320), .o1(new_n322));
  oaoi03aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(new_n314), .o1(new_n323));
  inv000aa1n03x5               g228(.a(new_n323), .o1(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n322), .c(new_n293), .d(new_n303), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .out0(new_n326));
  norp02aa1n02x5               g231(.a(new_n323), .b(new_n326), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n325), .b(new_n326), .c(new_n321), .d(new_n327), .o1(\s[30] ));
  nano22aa1n03x7               g233(.a(new_n313), .b(new_n316), .c(new_n326), .out0(new_n329));
  aoai13aa1n02x5               g234(.a(new_n329), .b(new_n297), .c(new_n199), .d(new_n292), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  oao003aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .c(new_n324), .carry(new_n332));
  norb02aa1n02x5               g237(.a(new_n332), .b(new_n331), .out0(new_n333));
  inv000aa1d42x5               g238(.a(new_n329), .o1(new_n334));
  aoai13aa1n03x5               g239(.a(new_n332), .b(new_n334), .c(new_n293), .d(new_n303), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n335), .b(new_n331), .c(new_n330), .d(new_n333), .o1(\s[31] ));
  norp02aa1n02x5               g241(.a(new_n105), .b(new_n102), .o1(new_n337));
  aoi022aa1n02x5               g242(.a(new_n131), .b(new_n101), .c(new_n99), .d(new_n107), .o1(new_n338));
  norp02aa1n02x5               g243(.a(new_n338), .b(new_n337), .o1(\s[3] ));
  nano22aa1n02x4               g244(.a(new_n337), .b(new_n107), .c(new_n106), .out0(new_n340));
  oaoi13aa1n02x5               g245(.a(new_n340), .b(new_n109), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g246(.a(new_n111), .b(new_n132), .c(new_n108), .out0(\s[5] ));
  orn002aa1n02x5               g247(.a(\a[5] ), .b(\b[4] ), .o(new_n343));
  nanp02aa1n02x5               g248(.a(new_n109), .b(new_n111), .o1(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n110), .b(new_n344), .c(new_n343), .out0(\s[6] ));
  nona22aa1n02x4               g250(.a(new_n109), .b(new_n133), .c(new_n134), .out0(new_n346));
  aob012aa1n02x5               g251(.a(new_n346), .b(new_n120), .c(new_n118), .out0(new_n347));
  xorb03aa1n02x5               g252(.a(new_n347), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp02aa1n02x5               g253(.a(new_n347), .b(new_n115), .o1(new_n349));
  xnbna2aa1n03x5               g254(.a(new_n112), .b(new_n349), .c(new_n122), .out0(\s[8] ));
  aoi112aa1n02x5               g255(.a(new_n124), .b(new_n125), .c(new_n109), .d(new_n117), .o1(new_n351));
  aoi012aa1n02x5               g256(.a(new_n351), .b(new_n137), .c(new_n125), .o1(\s[9] ));
endmodule


