// Benchmark "adder" written by ABC on Wed Jul 17 18:15:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n321, new_n322, new_n323, new_n325,
    new_n327, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nand22aa1n12x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  norp02aa1n24x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nona23aa1d18x5               g005(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n101));
  inv040aa1n06x5               g006(.a(new_n101), .o1(new_n102));
  aoi112aa1n06x5               g007(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n103));
  oab012aa1n09x5               g008(.a(new_n103), .b(\a[6] ), .c(\b[5] ), .out0(new_n104));
  ao0012aa1n03x7               g009(.a(new_n97), .b(new_n99), .c(new_n98), .o(new_n105));
  oabi12aa1n18x5               g010(.a(new_n105), .b(new_n101), .c(new_n104), .out0(new_n106));
  oaih22aa1n04x5               g011(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n107));
  xnrc02aa1n12x5               g012(.a(\b[2] ), .b(\a[3] ), .out0(new_n108));
  nand42aa1n06x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  nor042aa1n09x5               g014(.a(\b[1] ), .b(\a[2] ), .o1(new_n110));
  nand02aa1d16x5               g015(.a(\b[0] ), .b(\a[1] ), .o1(new_n111));
  oai012aa1n18x5               g016(.a(new_n109), .b(new_n110), .c(new_n111), .o1(new_n112));
  oabi12aa1n18x5               g017(.a(new_n107), .b(new_n108), .c(new_n112), .out0(new_n113));
  tech160nm_fixnrc02aa1n04x5   g018(.a(\b[5] ), .b(\a[6] ), .out0(new_n114));
  orn002aa1n24x5               g019(.a(\a[5] ), .b(\b[4] ), .o(new_n115));
  nanp02aa1n04x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanp02aa1n09x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  nanp03aa1d12x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  nor042aa1n06x5               g023(.a(new_n118), .b(new_n114), .o1(new_n119));
  aoi013aa1n09x5               g024(.a(new_n106), .b(new_n113), .c(new_n102), .d(new_n119), .o1(new_n120));
  oaoi03aa1n09x5               g025(.a(\a[9] ), .b(\b[8] ), .c(new_n120), .o1(new_n121));
  xorb03aa1n02x5               g026(.a(new_n121), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n04x5               g027(.a(\b[9] ), .b(\a[10] ), .o1(new_n123));
  nand02aa1d12x5               g028(.a(\b[9] ), .b(\a[10] ), .o1(new_n124));
  norb02aa1n06x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  nor042aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(new_n126), .b(new_n124), .o1(new_n127));
  oai012aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .o1(new_n128));
  tech160nm_fixnrc02aa1n05x5   g033(.a(\b[10] ), .b(\a[11] ), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n128), .c(new_n121), .d(new_n125), .o1(new_n130));
  nanp02aa1n03x5               g035(.a(new_n121), .b(new_n125), .o1(new_n131));
  nor002aa1n03x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  and002aa1n24x5               g037(.a(\b[10] ), .b(\a[11] ), .o(new_n133));
  nona32aa1n03x5               g038(.a(new_n131), .b(new_n133), .c(new_n132), .d(new_n128), .out0(new_n134));
  nanp02aa1n02x5               g039(.a(new_n134), .b(new_n130), .o1(\s[11] ));
  nor022aa1n12x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  tech160nm_finand02aa1n05x5   g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  nona22aa1n02x4               g043(.a(new_n134), .b(new_n138), .c(new_n133), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n133), .o1(new_n140));
  aob012aa1n03x5               g045(.a(new_n138), .b(new_n134), .c(new_n140), .out0(new_n141));
  nanp02aa1n03x5               g046(.a(new_n141), .b(new_n139), .o1(\s[12] ));
  inv040aa1n06x5               g047(.a(new_n106), .o1(new_n143));
  nand23aa1n09x5               g048(.a(new_n113), .b(new_n102), .c(new_n119), .o1(new_n144));
  xnrc02aa1n12x5               g049(.a(\b[8] ), .b(\a[9] ), .out0(new_n145));
  inv000aa1n02x5               g050(.a(new_n125), .o1(new_n146));
  inv000aa1n02x5               g051(.a(new_n136), .o1(new_n147));
  nano22aa1n03x7               g052(.a(new_n129), .b(new_n147), .c(new_n137), .out0(new_n148));
  nona22aa1n06x5               g053(.a(new_n148), .b(new_n146), .c(new_n145), .out0(new_n149));
  nona22aa1n03x5               g054(.a(new_n127), .b(new_n132), .c(new_n123), .out0(new_n150));
  aoai13aa1n12x5               g055(.a(new_n137), .b(new_n136), .c(new_n150), .d(new_n140), .o1(new_n151));
  aoai13aa1n12x5               g056(.a(new_n151), .b(new_n149), .c(new_n144), .d(new_n143), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand02aa1d06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  tech160nm_fiaoi012aa1n05x5   g060(.a(new_n154), .b(new_n152), .c(new_n155), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand02aa1d16x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nona23aa1d18x5               g064(.a(new_n159), .b(new_n155), .c(new_n154), .d(new_n158), .out0(new_n160));
  inv040aa1n03x5               g065(.a(new_n160), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n158), .b(new_n154), .c(new_n159), .o1(new_n162));
  inv000aa1n02x5               g067(.a(new_n162), .o1(new_n163));
  nor002aa1d32x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand22aa1n12x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanb02aa1d36x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n163), .c(new_n152), .d(new_n161), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n167), .b(new_n163), .c(new_n152), .d(new_n161), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(\s[15] ));
  inv000aa1d42x5               g075(.a(new_n164), .o1(new_n171));
  xnrc02aa1n12x5               g076(.a(\b[15] ), .b(\a[16] ), .out0(new_n172));
  xobna2aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n171), .out0(\s[16] ));
  nand02aa1d10x5               g078(.a(new_n144), .b(new_n143), .o1(new_n174));
  nona22aa1n09x5               g079(.a(new_n161), .b(new_n172), .c(new_n166), .out0(new_n175));
  nor042aa1n06x5               g080(.a(new_n175), .b(new_n149), .o1(new_n176));
  nand02aa1d06x5               g081(.a(new_n174), .b(new_n176), .o1(new_n177));
  aoi112aa1n03x4               g082(.a(new_n123), .b(new_n132), .c(new_n126), .d(new_n124), .o1(new_n178));
  oai012aa1n03x5               g083(.a(new_n147), .b(new_n178), .c(new_n133), .o1(new_n179));
  nor043aa1n06x5               g084(.a(new_n160), .b(new_n166), .c(new_n172), .o1(new_n180));
  orn002aa1n02x5               g085(.a(\a[16] ), .b(\b[15] ), .o(new_n181));
  and002aa1n02x5               g086(.a(\b[15] ), .b(\a[16] ), .o(new_n182));
  aoai13aa1n04x5               g087(.a(new_n165), .b(new_n158), .c(new_n154), .d(new_n159), .o1(new_n183));
  aoai13aa1n06x5               g088(.a(new_n181), .b(new_n182), .c(new_n183), .d(new_n171), .o1(new_n184));
  aoi013aa1n06x4               g089(.a(new_n184), .b(new_n180), .c(new_n179), .d(new_n137), .o1(new_n185));
  tech160nm_fixorc02aa1n03p5x5 g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n177), .c(new_n185), .out0(\s[17] ));
  inv040aa1d32x5               g092(.a(\a[17] ), .o1(new_n188));
  inv040aa1d28x5               g093(.a(\b[16] ), .o1(new_n189));
  nanp02aa1n04x5               g094(.a(new_n189), .b(new_n188), .o1(new_n190));
  oabi12aa1n12x5               g095(.a(new_n184), .b(new_n151), .c(new_n175), .out0(new_n191));
  aoai13aa1n03x5               g096(.a(new_n186), .b(new_n191), .c(new_n174), .d(new_n176), .o1(new_n192));
  nor022aa1n08x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  nand02aa1d28x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  nanb02aa1d24x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  xobna2aa1n03x5               g100(.a(new_n195), .b(new_n192), .c(new_n190), .out0(\s[18] ));
  norb02aa1n02x5               g101(.a(new_n186), .b(new_n195), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n191), .c(new_n174), .d(new_n176), .o1(new_n198));
  aoi013aa1n09x5               g103(.a(new_n193), .b(new_n194), .c(new_n188), .d(new_n189), .o1(new_n199));
  nor002aa1d32x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand42aa1d28x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n198), .c(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n06x5               g109(.a(new_n198), .b(new_n199), .o1(new_n205));
  nor002aa1d32x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nand42aa1d28x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nanb02aa1n02x5               g112(.a(new_n206), .b(new_n207), .out0(new_n208));
  aoai13aa1n03x5               g113(.a(new_n208), .b(new_n200), .c(new_n205), .d(new_n202), .o1(new_n209));
  nona23aa1n06x5               g114(.a(new_n180), .b(new_n148), .c(new_n145), .d(new_n146), .out0(new_n210));
  oai012aa1n06x5               g115(.a(new_n185), .b(new_n120), .c(new_n210), .o1(new_n211));
  oaoi03aa1n09x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n190), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n202), .b(new_n212), .c(new_n211), .d(new_n197), .o1(new_n213));
  nona22aa1n02x4               g118(.a(new_n213), .b(new_n208), .c(new_n200), .out0(new_n214));
  nanp02aa1n03x5               g119(.a(new_n209), .b(new_n214), .o1(\s[20] ));
  nona23aa1d24x5               g120(.a(new_n207), .b(new_n201), .c(new_n200), .d(new_n206), .out0(new_n216));
  norb03aa1n12x5               g121(.a(new_n186), .b(new_n216), .c(new_n195), .out0(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n191), .c(new_n174), .d(new_n176), .o1(new_n218));
  oai012aa1n12x5               g123(.a(new_n207), .b(new_n206), .c(new_n200), .o1(new_n219));
  oai012aa1d24x5               g124(.a(new_n219), .b(new_n216), .c(new_n199), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  xorc02aa1n12x5               g126(.a(\a[21] ), .b(\b[20] ), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n218), .c(new_n221), .out0(\s[21] ));
  nand02aa1n03x5               g128(.a(new_n218), .b(new_n221), .o1(new_n224));
  nor042aa1d18x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n225), .c(new_n224), .d(new_n222), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n222), .b(new_n220), .c(new_n211), .d(new_n217), .o1(new_n228));
  nona22aa1n02x4               g133(.a(new_n228), .b(new_n226), .c(new_n225), .out0(new_n229));
  nanp02aa1n02x5               g134(.a(new_n227), .b(new_n229), .o1(\s[22] ));
  nano23aa1n09x5               g135(.a(new_n200), .b(new_n206), .c(new_n207), .d(new_n201), .out0(new_n231));
  norb02aa1n06x4               g136(.a(new_n222), .b(new_n226), .out0(new_n232));
  nand03aa1n02x5               g137(.a(new_n232), .b(new_n197), .c(new_n231), .o1(new_n233));
  nand02aa1d06x5               g138(.a(new_n231), .b(new_n212), .o1(new_n234));
  nanb02aa1n12x5               g139(.a(new_n226), .b(new_n222), .out0(new_n235));
  inv000aa1n09x5               g140(.a(\a[22] ), .o1(new_n236));
  inv040aa1d32x5               g141(.a(\b[21] ), .o1(new_n237));
  oao003aa1n03x5               g142(.a(new_n236), .b(new_n237), .c(new_n225), .carry(new_n238));
  inv040aa1n03x5               g143(.a(new_n238), .o1(new_n239));
  aoai13aa1n12x5               g144(.a(new_n239), .b(new_n235), .c(new_n234), .d(new_n219), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n233), .c(new_n177), .d(new_n185), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  tech160nm_fixorc02aa1n02p5x5 g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  xnrc02aa1n02x5               g150(.a(\b[23] ), .b(\a[24] ), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n244), .c(new_n242), .d(new_n245), .o1(new_n247));
  nanp02aa1n02x5               g152(.a(new_n242), .b(new_n245), .o1(new_n248));
  nona22aa1n02x4               g153(.a(new_n248), .b(new_n246), .c(new_n244), .out0(new_n249));
  nanp02aa1n03x5               g154(.a(new_n249), .b(new_n247), .o1(\s[24] ));
  norb02aa1n09x5               g155(.a(new_n245), .b(new_n246), .out0(new_n251));
  and003aa1n02x5               g156(.a(new_n217), .b(new_n251), .c(new_n232), .o(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n191), .c(new_n174), .d(new_n176), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n251), .b(new_n238), .c(new_n220), .d(new_n232), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\a[24] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(\b[23] ), .o1(new_n256));
  oao003aa1n02x5               g161(.a(new_n255), .b(new_n256), .c(new_n244), .carry(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  nand42aa1n02x5               g163(.a(new_n254), .b(new_n258), .o1(new_n259));
  nanb02aa1n06x5               g164(.a(new_n259), .b(new_n253), .out0(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  xorc02aa1n12x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  nor042aa1n06x5               g168(.a(\b[25] ), .b(\a[26] ), .o1(new_n264));
  nand42aa1d28x5               g169(.a(\b[25] ), .b(\a[26] ), .o1(new_n265));
  norb02aa1n12x5               g170(.a(new_n265), .b(new_n264), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n262), .c(new_n260), .d(new_n263), .o1(new_n268));
  aoai13aa1n02x5               g173(.a(new_n263), .b(new_n259), .c(new_n211), .d(new_n252), .o1(new_n269));
  nona22aa1n02x4               g174(.a(new_n269), .b(new_n267), .c(new_n262), .out0(new_n270));
  nanp02aa1n03x5               g175(.a(new_n268), .b(new_n270), .o1(\s[26] ));
  nand22aa1n12x5               g176(.a(new_n263), .b(new_n266), .o1(new_n272));
  nona23aa1n09x5               g177(.a(new_n217), .b(new_n251), .c(new_n235), .d(new_n272), .out0(new_n273));
  inv040aa1n03x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n191), .c(new_n174), .d(new_n176), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n272), .o1(new_n276));
  aoai13aa1n04x5               g181(.a(new_n276), .b(new_n257), .c(new_n240), .d(new_n251), .o1(new_n277));
  oai012aa1n02x5               g182(.a(new_n265), .b(new_n264), .c(new_n262), .o1(new_n278));
  nanp03aa1n03x5               g183(.a(new_n275), .b(new_n277), .c(new_n278), .o1(new_n279));
  xorb03aa1n02x5               g184(.a(new_n279), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g185(.a(\b[26] ), .b(\a[27] ), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n281), .c(new_n279), .d(new_n282), .o1(new_n284));
  oaoi13aa1n09x5               g189(.a(new_n273), .b(new_n185), .c(new_n120), .d(new_n210), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n278), .b(new_n272), .c(new_n254), .d(new_n258), .o1(new_n286));
  oaih12aa1n02x5               g191(.a(new_n282), .b(new_n286), .c(new_n285), .o1(new_n287));
  nona22aa1n02x5               g192(.a(new_n287), .b(new_n283), .c(new_n281), .out0(new_n288));
  nanp02aa1n03x5               g193(.a(new_n284), .b(new_n288), .o1(\s[28] ));
  norb02aa1n02x5               g194(.a(new_n282), .b(new_n283), .out0(new_n290));
  oaih12aa1n02x5               g195(.a(new_n290), .b(new_n286), .c(new_n285), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .out0(new_n292));
  inv000aa1d42x5               g197(.a(\a[28] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  aoi112aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n295));
  aoi112aa1n02x5               g200(.a(new_n292), .b(new_n295), .c(new_n293), .d(new_n294), .o1(new_n296));
  aoi012aa1n02x5               g201(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n297));
  nanp02aa1n03x5               g202(.a(new_n291), .b(new_n297), .o1(new_n298));
  aoi022aa1n02x7               g203(.a(new_n298), .b(new_n292), .c(new_n291), .d(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n111), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g205(.a(new_n283), .b(new_n292), .c(new_n282), .out0(new_n301));
  oabi12aa1n03x5               g206(.a(new_n301), .b(new_n286), .c(new_n285), .out0(new_n302));
  xorc02aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .o1(new_n304));
  aoi012aa1n02x5               g209(.a(new_n297), .b(\a[29] ), .c(\b[28] ), .o1(new_n305));
  norp03aa1n02x5               g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n307));
  nanp02aa1n03x5               g212(.a(new_n302), .b(new_n307), .o1(new_n308));
  aoi022aa1n02x7               g213(.a(new_n308), .b(new_n303), .c(new_n302), .d(new_n306), .o1(\s[30] ));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  norb02aa1n02x5               g215(.a(new_n303), .b(new_n301), .out0(new_n311));
  oaih12aa1n02x5               g216(.a(new_n311), .b(new_n286), .c(new_n285), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n313));
  aoi012aa1n03x5               g218(.a(new_n310), .b(new_n312), .c(new_n313), .o1(new_n314));
  inv000aa1n02x5               g219(.a(new_n311), .o1(new_n315));
  aoi013aa1n02x5               g220(.a(new_n315), .b(new_n275), .c(new_n277), .d(new_n278), .o1(new_n316));
  nano22aa1n02x4               g221(.a(new_n316), .b(new_n310), .c(new_n313), .out0(new_n317));
  norp02aa1n03x5               g222(.a(new_n314), .b(new_n317), .o1(\s[31] ));
  inv000aa1d42x5               g223(.a(\a[3] ), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n112), .b(\b[2] ), .c(new_n319), .out0(\s[3] ));
  norp02aa1n02x5               g225(.a(new_n108), .b(new_n112), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[4] ), .b(\b[3] ), .out0(new_n322));
  aoib12aa1n02x5               g227(.a(new_n322), .b(new_n319), .c(\b[2] ), .out0(new_n323));
  aboi22aa1n03x5               g228(.a(new_n321), .b(new_n323), .c(new_n113), .d(new_n322), .out0(\s[4] ));
  aoi022aa1n02x5               g229(.a(new_n113), .b(new_n117), .c(new_n115), .d(new_n116), .o1(new_n325));
  aoib12aa1n02x5               g230(.a(new_n325), .b(new_n113), .c(new_n118), .out0(\s[5] ));
  oaib12aa1n02x5               g231(.a(new_n115), .b(new_n118), .c(new_n113), .out0(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aob012aa1n02x5               g233(.a(new_n104), .b(new_n113), .c(new_n119), .out0(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g235(.a(new_n99), .b(new_n329), .c(new_n100), .o1(new_n331));
  xnrb03aa1n02x5               g236(.a(new_n331), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g237(.a(new_n145), .b(new_n144), .c(new_n143), .out0(\s[9] ));
endmodule


