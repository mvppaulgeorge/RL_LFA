// Benchmark "adder" written by ABC on Wed Jul 17 23:36:11 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n316, new_n317,
    new_n319, new_n320, new_n321, new_n323, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[8] ), .o1(new_n101));
  xnrc02aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .out0(new_n102));
  nanp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n03x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  tech160nm_fioai012aa1n05x5   g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\a[3] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[4] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[2] ), .o1(new_n109));
  aboi22aa1n03x5               g014(.a(\b[3] ), .b(new_n108), .c(new_n107), .d(new_n109), .out0(new_n110));
  tech160nm_fioai012aa1n05x5   g015(.a(new_n110), .b(new_n102), .c(new_n106), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  oai112aa1n02x5               g018(.a(new_n112), .b(new_n113), .c(\b[5] ), .d(\a[6] ), .o1(new_n114));
  nand22aa1n12x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\a[8] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[7] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  oai112aa1n02x5               g023(.a(new_n118), .b(new_n115), .c(\b[6] ), .d(\a[7] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[3] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  oai122aa1n02x7               g026(.a(new_n121), .b(new_n108), .c(new_n120), .d(\a[5] ), .e(\b[4] ), .o1(new_n122));
  nor043aa1n02x5               g027(.a(new_n119), .b(new_n122), .c(new_n114), .o1(new_n123));
  nand02aa1n04x5               g028(.a(new_n123), .b(new_n111), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\a[7] ), .o1(new_n125));
  inv000aa1d42x5               g030(.a(\b[6] ), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(new_n126), .b(new_n125), .o1(new_n127));
  oai022aa1n06x5               g032(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n128));
  nanp03aa1n03x5               g033(.a(new_n128), .b(new_n113), .c(new_n121), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(new_n129), .b(new_n127), .o1(new_n130));
  tech160nm_fioaoi03aa1n03p5x5 g035(.a(new_n116), .b(new_n117), .c(new_n130), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(new_n131), .b(new_n124), .o1(new_n132));
  tech160nm_fioaoi03aa1n03p5x5 g037(.a(new_n100), .b(new_n101), .c(new_n132), .o1(new_n133));
  oabi12aa1n02x5               g038(.a(new_n133), .b(new_n97), .c(new_n99), .out0(new_n134));
  nona22aa1n03x5               g039(.a(new_n133), .b(new_n99), .c(new_n97), .out0(new_n135));
  nanp02aa1n02x5               g040(.a(new_n134), .b(new_n135), .o1(\s[10] ));
  inv000aa1d42x5               g041(.a(\a[11] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(\b[10] ), .o1(new_n138));
  nand42aa1n02x5               g043(.a(new_n138), .b(new_n137), .o1(new_n139));
  nanp02aa1n04x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(new_n139), .b(new_n140), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n135), .c(new_n98), .out0(\s[11] ));
  nona22aa1n03x5               g047(.a(new_n135), .b(new_n141), .c(new_n99), .out0(new_n143));
  xnrc02aa1n02x5               g048(.a(\b[11] ), .b(\a[12] ), .out0(new_n144));
  tech160nm_fiaoi012aa1n02p5x5 g049(.a(new_n144), .b(new_n143), .c(new_n139), .o1(new_n145));
  nanp03aa1n02x5               g050(.a(new_n143), .b(new_n139), .c(new_n144), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(\s[12] ));
  norp02aa1n09x5               g052(.a(\b[8] ), .b(\a[9] ), .o1(new_n148));
  norb03aa1n02x5               g053(.a(new_n98), .b(new_n97), .c(new_n148), .out0(new_n149));
  oai112aa1n03x5               g054(.a(new_n139), .b(new_n140), .c(new_n101), .d(new_n100), .o1(new_n150));
  nona22aa1n03x5               g055(.a(new_n149), .b(new_n150), .c(new_n144), .out0(new_n151));
  oai112aa1n06x5               g056(.a(new_n140), .b(new_n98), .c(new_n148), .d(new_n97), .o1(new_n152));
  oa0022aa1n06x5               g057(.a(\a[12] ), .b(\b[11] ), .c(\a[11] ), .d(\b[10] ), .o(new_n153));
  aoi022aa1d18x5               g058(.a(new_n152), .b(new_n153), .c(\b[11] ), .d(\a[12] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n151), .c(new_n131), .d(new_n124), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv030aa1d32x5               g062(.a(\a[13] ), .o1(new_n158));
  inv000aa1n30x5               g063(.a(\b[12] ), .o1(new_n159));
  oaoi03aa1n02x5               g064(.a(new_n158), .b(new_n159), .c(new_n156), .o1(new_n160));
  xnrb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nor002aa1d32x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nand42aa1n08x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n162), .b(new_n164), .c(new_n165), .d(new_n163), .out0(new_n166));
  aoai13aa1n12x5               g071(.a(new_n165), .b(new_n164), .c(new_n158), .d(new_n159), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  orn002aa1n24x5               g073(.a(\a[15] ), .b(\b[14] ), .o(new_n169));
  nanp02aa1n06x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nanp02aa1n09x5               g075(.a(new_n169), .b(new_n170), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n156), .d(new_n166), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n172), .b(new_n168), .c(new_n156), .d(new_n166), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(\s[15] ));
  nor002aa1n20x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nanb02aa1n03x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  xobna2aa1n03x5               g083(.a(new_n178), .b(new_n173), .c(new_n169), .out0(\s[16] ));
  norb03aa1n02x5               g084(.a(new_n149), .b(new_n144), .c(new_n150), .out0(new_n180));
  nona23aa1n03x5               g085(.a(new_n165), .b(new_n163), .c(new_n162), .d(new_n164), .out0(new_n181));
  nor003aa1n06x5               g086(.a(new_n181), .b(new_n171), .c(new_n178), .o1(new_n182));
  nand02aa1n02x5               g087(.a(new_n180), .b(new_n182), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n176), .o1(new_n184));
  nand02aa1n02x5               g089(.a(new_n177), .b(new_n170), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n184), .b(new_n185), .c(new_n167), .d(new_n169), .o1(new_n186));
  aoi012aa1n12x5               g091(.a(new_n186), .b(new_n182), .c(new_n154), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n183), .c(new_n131), .d(new_n124), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g094(.a(\a[18] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\a[17] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[16] ), .o1(new_n192));
  oaoi03aa1n02x5               g097(.a(new_n191), .b(new_n192), .c(new_n188), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[17] ), .c(new_n190), .out0(\s[18] ));
  xroi22aa1d04x5               g099(.a(new_n191), .b(\b[16] ), .c(new_n190), .d(\b[17] ), .out0(new_n195));
  nor042aa1n02x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  aoi112aa1n06x5               g101(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n197));
  nor042aa1n06x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  nor002aa1n10x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand42aa1n02x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  norb02aa1n03x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n188), .d(new_n195), .o1(new_n203));
  aoi112aa1n02x5               g108(.a(new_n202), .b(new_n199), .c(new_n188), .d(new_n195), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g111(.a(new_n200), .o1(new_n207));
  nor042aa1n03x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nanp02aa1n04x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n03x4               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  xnbna2aa1n03x5               g115(.a(new_n210), .b(new_n203), .c(new_n207), .out0(\s[20] ));
  inv000aa1d42x5               g116(.a(new_n115), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n118), .b(new_n212), .c(new_n129), .d(new_n127), .o1(new_n213));
  nona22aa1n09x5               g118(.a(new_n166), .b(new_n171), .c(new_n178), .out0(new_n214));
  nor002aa1n02x5               g119(.a(new_n151), .b(new_n214), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n213), .c(new_n111), .d(new_n123), .o1(new_n216));
  nona23aa1d18x5               g121(.a(new_n209), .b(new_n201), .c(new_n200), .d(new_n208), .out0(new_n217));
  inv000aa1n06x5               g122(.a(new_n217), .o1(new_n218));
  nanp02aa1n06x5               g123(.a(new_n195), .b(new_n218), .o1(new_n219));
  tech160nm_fioai012aa1n04x5   g124(.a(new_n209), .b(new_n208), .c(new_n200), .o1(new_n220));
  oai012aa1n18x5               g125(.a(new_n220), .b(new_n217), .c(new_n198), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n222), .b(new_n219), .c(new_n216), .d(new_n187), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xorc02aa1n02x5               g130(.a(\a[21] ), .b(\b[20] ), .out0(new_n226));
  xorc02aa1n02x5               g131(.a(\a[22] ), .b(\b[21] ), .out0(new_n227));
  aoi112aa1n02x5               g132(.a(new_n225), .b(new_n227), .c(new_n223), .d(new_n226), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n227), .b(new_n225), .c(new_n223), .d(new_n226), .o1(new_n229));
  norb02aa1n02x7               g134(.a(new_n229), .b(new_n228), .out0(\s[22] ));
  nand02aa1d04x5               g135(.a(new_n227), .b(new_n226), .o1(new_n231));
  nano22aa1n02x4               g136(.a(new_n231), .b(new_n195), .c(new_n218), .out0(new_n232));
  oai112aa1n03x5               g137(.a(new_n202), .b(new_n210), .c(new_n197), .d(new_n196), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\a[22] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(\b[21] ), .o1(new_n235));
  oao003aa1n06x5               g140(.a(new_n234), .b(new_n235), .c(new_n225), .carry(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n237), .b(new_n231), .c(new_n233), .d(new_n220), .o1(new_n238));
  xorc02aa1n02x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n238), .c(new_n188), .d(new_n232), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(new_n239), .b(new_n238), .c(new_n188), .d(new_n232), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n240), .b(new_n241), .out0(\s[23] ));
  inv000aa1d42x5               g147(.a(\a[23] ), .o1(new_n243));
  nanb02aa1n12x5               g148(.a(\b[22] ), .b(new_n243), .out0(new_n244));
  xorc02aa1n02x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  xnbna2aa1n03x5               g150(.a(new_n245), .b(new_n240), .c(new_n244), .out0(\s[24] ));
  inv000aa1d42x5               g151(.a(\a[24] ), .o1(new_n247));
  xroi22aa1d04x5               g152(.a(new_n243), .b(\b[22] ), .c(new_n247), .d(\b[23] ), .out0(new_n248));
  nano32aa1n03x7               g153(.a(new_n219), .b(new_n248), .c(new_n226), .d(new_n227), .out0(new_n249));
  inv000aa1n02x5               g154(.a(new_n231), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n248), .b(new_n236), .c(new_n221), .d(new_n250), .o1(new_n251));
  oaoi03aa1n03x5               g156(.a(\a[24] ), .b(\b[23] ), .c(new_n244), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  nand42aa1n02x5               g158(.a(new_n251), .b(new_n253), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n188), .d(new_n249), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n254), .b(new_n255), .c(new_n188), .d(new_n249), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n256), .b(new_n257), .out0(\s[25] ));
  inv000aa1d42x5               g163(.a(\a[25] ), .o1(new_n259));
  nanb02aa1n02x5               g164(.a(\b[24] ), .b(new_n259), .out0(new_n260));
  xorc02aa1n02x5               g165(.a(\a[26] ), .b(\b[25] ), .out0(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n256), .c(new_n260), .out0(\s[26] ));
  inv000aa1d42x5               g167(.a(\a[26] ), .o1(new_n263));
  xroi22aa1d06x4               g168(.a(new_n259), .b(\b[24] ), .c(new_n263), .d(\b[25] ), .out0(new_n264));
  nano32aa1n03x5               g169(.a(new_n219), .b(new_n264), .c(new_n250), .d(new_n248), .out0(new_n265));
  nanp02aa1n09x5               g170(.a(new_n188), .b(new_n265), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n264), .b(new_n252), .c(new_n238), .d(new_n248), .o1(new_n267));
  oao003aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .c(new_n260), .carry(new_n268));
  norp02aa1n02x5               g173(.a(\b[26] ), .b(\a[27] ), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n270), .b(new_n269), .out0(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  aoi013aa1n06x4               g177(.a(new_n272), .b(new_n266), .c(new_n267), .d(new_n268), .o1(new_n273));
  nand02aa1n02x5               g178(.a(new_n249), .b(new_n264), .o1(new_n274));
  tech160nm_fiaoi012aa1n03p5x5 g179(.a(new_n274), .b(new_n216), .c(new_n187), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n264), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n268), .b(new_n276), .c(new_n251), .d(new_n253), .o1(new_n277));
  norp03aa1n02x5               g182(.a(new_n277), .b(new_n275), .c(new_n271), .o1(new_n278));
  norp02aa1n02x5               g183(.a(new_n273), .b(new_n278), .o1(\s[27] ));
  inv020aa1n02x5               g184(.a(new_n269), .o1(new_n280));
  tech160nm_fixnrc02aa1n05x5   g185(.a(\b[27] ), .b(\a[28] ), .out0(new_n281));
  nano22aa1n03x7               g186(.a(new_n273), .b(new_n280), .c(new_n281), .out0(new_n282));
  oai012aa1n02x5               g187(.a(new_n271), .b(new_n277), .c(new_n275), .o1(new_n283));
  aoi012aa1n03x5               g188(.a(new_n281), .b(new_n283), .c(new_n280), .o1(new_n284));
  norp02aa1n03x5               g189(.a(new_n284), .b(new_n282), .o1(\s[28] ));
  nano22aa1n06x5               g190(.a(new_n281), .b(new_n280), .c(new_n270), .out0(new_n286));
  oai012aa1n02x5               g191(.a(new_n286), .b(new_n277), .c(new_n275), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[28] ), .b(\a[29] ), .out0(new_n289));
  aoi012aa1n02x5               g194(.a(new_n289), .b(new_n287), .c(new_n288), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n286), .o1(new_n291));
  aoi013aa1n03x5               g196(.a(new_n291), .b(new_n266), .c(new_n267), .d(new_n268), .o1(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n288), .c(new_n289), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n290), .b(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g200(.a(new_n289), .b(new_n281), .c(new_n270), .d(new_n280), .out0(new_n296));
  oai012aa1n02x5               g201(.a(new_n296), .b(new_n277), .c(new_n275), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n288), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[29] ), .b(\a[30] ), .out0(new_n299));
  aoi012aa1n02x5               g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n296), .o1(new_n301));
  aoi013aa1n03x5               g206(.a(new_n301), .b(new_n266), .c(new_n267), .d(new_n268), .o1(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n298), .c(new_n299), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n300), .b(new_n303), .o1(\s[30] ));
  norb03aa1n02x5               g209(.a(new_n286), .b(new_n299), .c(new_n289), .out0(new_n305));
  inv000aa1n02x5               g210(.a(new_n305), .o1(new_n306));
  aoi013aa1n03x5               g211(.a(new_n306), .b(new_n266), .c(new_n267), .d(new_n268), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[30] ), .b(\a[31] ), .out0(new_n309));
  nano22aa1n03x5               g214(.a(new_n307), .b(new_n308), .c(new_n309), .out0(new_n310));
  oai012aa1n02x5               g215(.a(new_n305), .b(new_n277), .c(new_n275), .o1(new_n311));
  aoi012aa1n02x5               g216(.a(new_n309), .b(new_n311), .c(new_n308), .o1(new_n312));
  norp02aa1n03x5               g217(.a(new_n312), .b(new_n310), .o1(\s[31] ));
  xorb03aa1n02x5               g218(.a(new_n106), .b(\b[2] ), .c(new_n107), .out0(\s[3] ));
  norp02aa1n02x5               g219(.a(new_n102), .b(new_n106), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[4] ), .b(\b[3] ), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n316), .b(new_n107), .c(new_n109), .o1(new_n317));
  aboi22aa1n03x5               g222(.a(new_n315), .b(new_n317), .c(new_n111), .d(new_n316), .out0(\s[4] ));
  xorc02aa1n02x5               g223(.a(\a[5] ), .b(\b[4] ), .out0(new_n319));
  oaoi13aa1n02x5               g224(.a(new_n319), .b(new_n111), .c(new_n108), .d(new_n120), .o1(new_n320));
  oai112aa1n02x5               g225(.a(new_n111), .b(new_n319), .c(new_n120), .d(new_n108), .o1(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(\s[5] ));
  oa0012aa1n02x5               g227(.a(new_n321), .b(\b[4] ), .c(\a[5] ), .o(new_n323));
  xnrb03aa1n02x5               g228(.a(new_n323), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g229(.a(\a[6] ), .b(\b[5] ), .c(new_n323), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g231(.a(new_n125), .b(new_n126), .c(new_n325), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n327), .b(new_n115), .c(new_n118), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n132), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


