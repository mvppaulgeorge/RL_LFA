// Benchmark "adder" written by ABC on Wed Jul 17 15:27:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n319, new_n320, new_n323, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[2] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[1] ), .o1(new_n101));
  nand02aa1d08x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  tech160nm_fioaoi03aa1n02p5x5 g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nanp02aa1n09x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n16x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n104), .b(new_n107), .c(new_n106), .d(new_n105), .out0(new_n108));
  inv000aa1d42x5               g013(.a(\a[3] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  aoai13aa1n04x5               g015(.a(new_n104), .b(new_n105), .c(new_n110), .d(new_n109), .o1(new_n111));
  oai012aa1n06x5               g016(.a(new_n111), .b(new_n108), .c(new_n103), .o1(new_n112));
  nand02aa1d12x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand02aa1d06x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n113), .b(new_n116), .c(new_n115), .d(new_n114), .out0(new_n117));
  tech160nm_fixnrc02aa1n02p5x5 g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  tech160nm_fixnrc02aa1n02p5x5 g023(.a(\b[5] ), .b(\a[6] ), .out0(new_n119));
  nor003aa1n03x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n113), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n114), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n115), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\a[6] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[5] ), .o1(new_n125));
  oai022aa1d18x5               g030(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n126));
  oai112aa1n04x5               g031(.a(new_n126), .b(new_n116), .c(new_n125), .d(new_n124), .o1(new_n127));
  aoai13aa1n12x5               g032(.a(new_n122), .b(new_n121), .c(new_n127), .d(new_n123), .o1(new_n128));
  xorc02aa1n02x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n128), .c(new_n112), .d(new_n120), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n97), .b(new_n130), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g036(.a(new_n97), .o1(new_n132));
  aoi112aa1n09x5               g037(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n133));
  oab012aa1n12x5               g038(.a(new_n133), .b(\a[10] ), .c(\b[9] ), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n134), .b(new_n132), .c(new_n130), .d(new_n99), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanp02aa1n12x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nor002aa1d32x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand02aa1d06x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n137), .c(new_n135), .d(new_n138), .o1(new_n142));
  aoi112aa1n02x5               g047(.a(new_n137), .b(new_n141), .c(new_n135), .d(new_n138), .o1(new_n143));
  nanb02aa1n03x5               g048(.a(new_n143), .b(new_n142), .out0(\s[12] ));
  nona23aa1d18x5               g049(.a(new_n140), .b(new_n138), .c(new_n137), .d(new_n139), .out0(new_n145));
  nano22aa1n02x4               g050(.a(new_n145), .b(new_n97), .c(new_n129), .out0(new_n146));
  aoai13aa1n02x5               g051(.a(new_n146), .b(new_n128), .c(new_n112), .d(new_n120), .o1(new_n147));
  oa0012aa1n03x5               g052(.a(new_n140), .b(new_n139), .c(new_n137), .o(new_n148));
  oabi12aa1n18x5               g053(.a(new_n148), .b(new_n134), .c(new_n145), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nor042aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1n16x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n147), .c(new_n150), .out0(\s[13] ));
  orn002aa1n02x5               g059(.a(\a[13] ), .b(\b[12] ), .o(new_n155));
  oao003aa1n02x5               g060(.a(new_n100), .b(new_n101), .c(new_n102), .carry(new_n156));
  nano23aa1n03x5               g061(.a(new_n106), .b(new_n105), .c(new_n107), .d(new_n104), .out0(new_n157));
  aobi12aa1n02x5               g062(.a(new_n111), .b(new_n157), .c(new_n156), .out0(new_n158));
  nor042aa1n02x5               g063(.a(new_n119), .b(new_n118), .o1(new_n159));
  nanb02aa1n02x5               g064(.a(new_n117), .b(new_n159), .out0(new_n160));
  oabi12aa1n02x7               g065(.a(new_n128), .b(new_n158), .c(new_n160), .out0(new_n161));
  aoai13aa1n02x5               g066(.a(new_n153), .b(new_n149), .c(new_n161), .d(new_n146), .o1(new_n162));
  nor042aa1n04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n12x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  xobna2aa1n03x5               g070(.a(new_n165), .b(new_n162), .c(new_n155), .out0(\s[14] ));
  nano23aa1d15x5               g071(.a(new_n151), .b(new_n163), .c(new_n164), .d(new_n152), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoi012aa1n06x5               g073(.a(new_n163), .b(new_n151), .c(new_n164), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n168), .c(new_n147), .d(new_n150), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n03x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nor042aa1n06x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n177));
  aoi112aa1n02x5               g082(.a(new_n172), .b(new_n176), .c(new_n170), .d(new_n173), .o1(new_n178));
  nanb02aa1n03x5               g083(.a(new_n178), .b(new_n177), .out0(\s[16] ));
  nano23aa1n03x7               g084(.a(new_n137), .b(new_n139), .c(new_n140), .d(new_n138), .out0(new_n180));
  nano23aa1n03x5               g085(.a(new_n172), .b(new_n174), .c(new_n175), .d(new_n173), .out0(new_n181));
  nand02aa1d04x5               g086(.a(new_n181), .b(new_n167), .o1(new_n182));
  nano32aa1n03x7               g087(.a(new_n182), .b(new_n180), .c(new_n129), .d(new_n97), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n128), .c(new_n112), .d(new_n120), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n174), .o1(new_n185));
  tech160nm_fioaoi03aa1n03p5x5 g090(.a(\a[15] ), .b(\b[14] ), .c(new_n169), .o1(new_n186));
  nand42aa1n02x5               g091(.a(new_n186), .b(new_n175), .o1(new_n187));
  nanp02aa1n02x5               g092(.a(new_n187), .b(new_n185), .o1(new_n188));
  aoib12aa1n09x5               g093(.a(new_n188), .b(new_n149), .c(new_n182), .out0(new_n189));
  nanp02aa1n06x5               g094(.a(new_n189), .b(new_n184), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[18] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[16] ), .o1(new_n194));
  oaoi03aa1n03x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d06x4               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  nand22aa1n12x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nona22aa1n02x4               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(new_n199));
  oaib12aa1n09x5               g104(.a(new_n199), .b(\b[17] ), .c(new_n192), .out0(new_n200));
  nor042aa1n06x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nand02aa1n08x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n200), .c(new_n190), .d(new_n197), .o1(new_n204));
  aoi112aa1n02x5               g109(.a(new_n203), .b(new_n200), .c(new_n190), .d(new_n197), .o1(new_n205));
  norb02aa1n03x4               g110(.a(new_n204), .b(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1d08x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  tech160nm_fioai012aa1n03p5x5 g115(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .o1(new_n211));
  nanp02aa1n03x5               g116(.a(new_n211), .b(new_n210), .o1(new_n212));
  nona22aa1n02x5               g117(.a(new_n204), .b(new_n210), .c(new_n201), .out0(new_n213));
  nanp02aa1n03x5               g118(.a(new_n212), .b(new_n213), .o1(\s[20] ));
  nano23aa1n09x5               g119(.a(new_n201), .b(new_n208), .c(new_n209), .d(new_n202), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n197), .b(new_n215), .o1(new_n216));
  norp02aa1n02x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  aoi013aa1n06x5               g122(.a(new_n217), .b(new_n198), .c(new_n193), .d(new_n194), .o1(new_n218));
  nona23aa1n09x5               g123(.a(new_n209), .b(new_n202), .c(new_n201), .d(new_n208), .out0(new_n219));
  tech160nm_fioai012aa1n04x5   g124(.a(new_n209), .b(new_n208), .c(new_n201), .o1(new_n220));
  oai012aa1n12x5               g125(.a(new_n220), .b(new_n219), .c(new_n218), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n222), .b(new_n216), .c(new_n189), .d(new_n184), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  tech160nm_fixnrc02aa1n04x5   g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  aoai13aa1n02x5               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n229));
  aoi112aa1n03x4               g134(.a(new_n225), .b(new_n228), .c(new_n223), .d(new_n227), .o1(new_n230));
  nanb02aa1n03x5               g135(.a(new_n230), .b(new_n229), .out0(\s[22] ));
  nor042aa1n06x5               g136(.a(new_n228), .b(new_n226), .o1(new_n232));
  nand03aa1n02x5               g137(.a(new_n197), .b(new_n232), .c(new_n215), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\a[22] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(\b[21] ), .o1(new_n235));
  oaoi03aa1n12x5               g140(.a(new_n234), .b(new_n235), .c(new_n225), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi012aa1n02x5               g142(.a(new_n237), .b(new_n221), .c(new_n232), .o1(new_n238));
  aoai13aa1n04x5               g143(.a(new_n238), .b(new_n233), .c(new_n189), .d(new_n184), .o1(new_n239));
  xorb03aa1n02x5               g144(.a(new_n239), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  xorc02aa1n12x5               g146(.a(\a[23] ), .b(\b[22] ), .out0(new_n242));
  nor022aa1n12x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  nand42aa1n03x5               g148(.a(\b[23] ), .b(\a[24] ), .o1(new_n244));
  nanb02aa1n06x5               g149(.a(new_n243), .b(new_n244), .out0(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n241), .c(new_n239), .d(new_n242), .o1(new_n246));
  aoi112aa1n03x4               g151(.a(new_n241), .b(new_n245), .c(new_n239), .d(new_n242), .o1(new_n247));
  nanb02aa1n03x5               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  aoi012aa1n02x5               g153(.a(new_n174), .b(new_n186), .c(new_n175), .o1(new_n249));
  oaib12aa1n02x5               g154(.a(new_n249), .b(new_n182), .c(new_n149), .out0(new_n250));
  norb02aa1n02x7               g155(.a(new_n242), .b(new_n245), .out0(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  nano32aa1n02x4               g157(.a(new_n252), .b(new_n197), .c(new_n232), .d(new_n215), .out0(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n250), .c(new_n161), .d(new_n183), .o1(new_n254));
  inv000aa1n03x5               g159(.a(new_n220), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n232), .b(new_n255), .c(new_n215), .d(new_n200), .o1(new_n256));
  tech160nm_fioai012aa1n03p5x5 g161(.a(new_n244), .b(new_n243), .c(new_n241), .o1(new_n257));
  aoai13aa1n12x5               g162(.a(new_n257), .b(new_n252), .c(new_n256), .d(new_n236), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xorc02aa1n12x5               g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n254), .c(new_n259), .out0(\s[25] ));
  nand42aa1n02x5               g166(.a(new_n254), .b(new_n259), .o1(new_n262));
  norp02aa1n02x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  nor042aa1n04x5               g168(.a(\b[25] ), .b(\a[26] ), .o1(new_n264));
  nand02aa1d16x5               g169(.a(\b[25] ), .b(\a[26] ), .o1(new_n265));
  norb02aa1n09x5               g170(.a(new_n265), .b(new_n264), .out0(new_n266));
  inv000aa1n06x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n263), .c(new_n262), .d(new_n260), .o1(new_n268));
  aoai13aa1n02x5               g173(.a(new_n260), .b(new_n258), .c(new_n190), .d(new_n253), .o1(new_n269));
  nona22aa1n02x4               g174(.a(new_n269), .b(new_n267), .c(new_n263), .out0(new_n270));
  nanp02aa1n03x5               g175(.a(new_n268), .b(new_n270), .o1(\s[26] ));
  norb02aa1n12x5               g176(.a(new_n260), .b(new_n267), .out0(new_n272));
  nano22aa1n02x5               g177(.a(new_n233), .b(new_n272), .c(new_n251), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n250), .c(new_n161), .d(new_n183), .o1(new_n274));
  oai012aa1n02x5               g179(.a(new_n265), .b(new_n264), .c(new_n263), .o1(new_n275));
  aobi12aa1n12x5               g180(.a(new_n275), .b(new_n258), .c(new_n272), .out0(new_n276));
  xorc02aa1n02x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n276), .c(new_n274), .out0(\s[27] ));
  nand22aa1n03x5               g183(.a(new_n276), .b(new_n274), .o1(new_n279));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(\b[27] ), .b(\a[28] ), .o1(new_n281));
  nand42aa1n03x5               g186(.a(\b[27] ), .b(\a[28] ), .o1(new_n282));
  norb02aa1n03x5               g187(.a(new_n282), .b(new_n281), .out0(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n280), .c(new_n279), .d(new_n277), .o1(new_n285));
  aobi12aa1n06x5               g190(.a(new_n273), .b(new_n189), .c(new_n184), .out0(new_n286));
  aoai13aa1n04x5               g191(.a(new_n251), .b(new_n237), .c(new_n221), .d(new_n232), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n272), .o1(new_n288));
  aoai13aa1n04x5               g193(.a(new_n275), .b(new_n288), .c(new_n287), .d(new_n257), .o1(new_n289));
  oai012aa1n02x5               g194(.a(new_n277), .b(new_n289), .c(new_n286), .o1(new_n290));
  nona22aa1n02x4               g195(.a(new_n290), .b(new_n284), .c(new_n280), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n285), .b(new_n291), .o1(\s[28] ));
  norb02aa1n02x5               g197(.a(new_n277), .b(new_n284), .out0(new_n293));
  oai012aa1n02x5               g198(.a(new_n293), .b(new_n289), .c(new_n286), .o1(new_n294));
  aoi012aa1n02x5               g199(.a(new_n281), .b(new_n280), .c(new_n282), .o1(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[28] ), .b(\a[29] ), .out0(new_n296));
  tech160nm_fiaoi012aa1n02p5x5 g201(.a(new_n296), .b(new_n294), .c(new_n295), .o1(new_n297));
  aobi12aa1n06x5               g202(.a(new_n293), .b(new_n276), .c(new_n274), .out0(new_n298));
  nano22aa1n03x7               g203(.a(new_n298), .b(new_n295), .c(new_n296), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g206(.a(new_n296), .b(new_n277), .c(new_n283), .out0(new_n302));
  oai012aa1n02x5               g207(.a(new_n302), .b(new_n289), .c(new_n286), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[29] ), .b(\a[30] ), .out0(new_n305));
  tech160nm_fiaoi012aa1n02p5x5 g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  aobi12aa1n06x5               g211(.a(new_n302), .b(new_n276), .c(new_n274), .out0(new_n307));
  nano22aa1n03x7               g212(.a(new_n307), .b(new_n304), .c(new_n305), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n306), .b(new_n308), .o1(\s[30] ));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  nano23aa1n02x4               g215(.a(new_n305), .b(new_n296), .c(new_n277), .d(new_n283), .out0(new_n311));
  oai012aa1n02x5               g216(.a(new_n311), .b(new_n289), .c(new_n286), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .c(new_n304), .carry(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n310), .b(new_n312), .c(new_n313), .o1(new_n314));
  aobi12aa1n06x5               g219(.a(new_n311), .b(new_n276), .c(new_n274), .out0(new_n315));
  nano22aa1n03x7               g220(.a(new_n315), .b(new_n310), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[31] ));
  xorb03aa1n02x5               g222(.a(new_n103), .b(\b[2] ), .c(new_n109), .out0(\s[3] ));
  nanb03aa1n02x5               g223(.a(new_n106), .b(new_n156), .c(new_n107), .out0(new_n319));
  aboi22aa1n03x5               g224(.a(new_n105), .b(new_n104), .c(new_n110), .d(new_n109), .out0(new_n320));
  aboi22aa1n03x5               g225(.a(new_n105), .b(new_n112), .c(new_n319), .d(new_n320), .out0(\s[4] ));
  xorb03aa1n02x5               g226(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g227(.a(\a[5] ), .b(\b[4] ), .c(new_n158), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g229(.a(new_n124), .b(new_n125), .c(new_n323), .o1(new_n325));
  xnbna2aa1n03x5               g230(.a(new_n325), .b(new_n123), .c(new_n116), .out0(\s[7] ));
  oaoi03aa1n02x5               g231(.a(\a[7] ), .b(\b[6] ), .c(new_n325), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n161), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


