// Benchmark "adder" written by ABC on Thu Jul 18 07:09:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n306, new_n309, new_n311, new_n313, new_n315;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  xnrc02aa1n12x5               g006(.a(\b[7] ), .b(\a[8] ), .out0(new_n102));
  nor002aa1n10x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nanb02aa1n03x5               g009(.a(new_n103), .b(new_n104), .out0(new_n105));
  aoi112aa1n09x5               g010(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n106));
  oab012aa1n04x5               g011(.a(new_n106), .b(\a[6] ), .c(\b[5] ), .out0(new_n107));
  aoi112aa1n02x5               g012(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n108));
  oab012aa1n02x5               g013(.a(new_n108), .b(\a[8] ), .c(\b[7] ), .out0(new_n109));
  oai013aa1n06x5               g014(.a(new_n109), .b(new_n107), .c(new_n102), .d(new_n105), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  nand02aa1d04x5               g016(.a(\b[0] ), .b(\a[1] ), .o1(new_n112));
  nor042aa1n02x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  oai012aa1n09x5               g018(.a(new_n111), .b(new_n113), .c(new_n112), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  nor022aa1n16x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nor022aa1n08x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  tech160nm_finand02aa1n03p5x5 g022(.a(\b[3] ), .b(\a[4] ), .o1(new_n118));
  nona23aa1n09x5               g023(.a(new_n115), .b(new_n118), .c(new_n117), .d(new_n116), .out0(new_n119));
  tech160nm_fioai012aa1n03p5x5 g024(.a(new_n118), .b(new_n117), .c(new_n116), .o1(new_n120));
  oaih12aa1n12x5               g025(.a(new_n120), .b(new_n119), .c(new_n114), .o1(new_n121));
  nor022aa1n16x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  nand42aa1n03x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  nona23aa1n09x5               g028(.a(new_n123), .b(new_n104), .c(new_n103), .d(new_n122), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[5] ), .b(\a[6] ), .out0(new_n125));
  nor043aa1n06x5               g030(.a(new_n124), .b(new_n125), .c(new_n102), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n110), .c(new_n121), .d(new_n126), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n99), .b(new_n128), .c(new_n101), .out0(\s[10] ));
  inv000aa1d42x5               g034(.a(new_n97), .o1(new_n130));
  inv000aa1n02x5               g035(.a(new_n98), .o1(new_n131));
  aoai13aa1n03x5               g036(.a(new_n130), .b(new_n131), .c(new_n128), .d(new_n101), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n134), .o1(new_n135));
  nand02aa1d28x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nor002aa1n16x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand02aa1d20x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  aoi012aa1n02x5               g043(.a(new_n137), .b(new_n132), .c(new_n138), .o1(new_n139));
  nano22aa1n02x4               g044(.a(new_n139), .b(new_n135), .c(new_n136), .out0(new_n140));
  aoi122aa1n02x5               g045(.a(new_n137), .b(new_n135), .c(new_n136), .d(new_n132), .e(new_n138), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n140), .b(new_n141), .o1(\s[12] ));
  nona32aa1n09x5               g047(.a(new_n127), .b(new_n131), .c(new_n137), .d(new_n97), .out0(new_n143));
  nanb03aa1d24x5               g048(.a(new_n134), .b(new_n136), .c(new_n138), .out0(new_n144));
  norp02aa1n02x5               g049(.a(new_n143), .b(new_n144), .o1(new_n145));
  aoai13aa1n03x5               g050(.a(new_n145), .b(new_n110), .c(new_n121), .d(new_n126), .o1(new_n146));
  aoi012aa1d18x5               g051(.a(new_n97), .b(new_n100), .c(new_n98), .o1(new_n147));
  aoi012aa1n06x5               g052(.a(new_n134), .b(new_n137), .c(new_n136), .o1(new_n148));
  oai013aa1d12x5               g053(.a(new_n148), .b(new_n144), .c(new_n147), .d(new_n137), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nor042aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1d28x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  norb02aa1n06x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n146), .c(new_n150), .out0(\s[13] ));
  nanp02aa1n02x5               g059(.a(new_n146), .b(new_n150), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n151), .b(new_n155), .c(new_n152), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand22aa1n06x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nona23aa1n03x5               g064(.a(new_n159), .b(new_n152), .c(new_n151), .d(new_n158), .out0(new_n160));
  aoi012aa1n02x7               g065(.a(new_n158), .b(new_n151), .c(new_n159), .o1(new_n161));
  aoai13aa1n03x5               g066(.a(new_n161), .b(new_n160), .c(new_n146), .d(new_n150), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n06x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand02aa1d24x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nor042aa1d18x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand02aa1n12x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n164), .b(new_n168), .c(new_n162), .d(new_n165), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nano22aa1n02x4               g076(.a(new_n134), .b(new_n138), .c(new_n136), .out0(new_n172));
  nona23aa1n09x5               g077(.a(new_n153), .b(new_n159), .c(new_n164), .d(new_n158), .out0(new_n173));
  nanb03aa1d24x5               g078(.a(new_n166), .b(new_n167), .c(new_n165), .out0(new_n174));
  inv040aa1n03x5               g079(.a(new_n174), .o1(new_n175));
  nano23aa1n06x5               g080(.a(new_n143), .b(new_n173), .c(new_n175), .d(new_n172), .out0(new_n176));
  aoai13aa1n12x5               g081(.a(new_n176), .b(new_n110), .c(new_n126), .d(new_n121), .o1(new_n177));
  nor043aa1n03x5               g082(.a(new_n160), .b(new_n164), .c(new_n174), .o1(new_n178));
  norp03aa1n04x5               g083(.a(new_n174), .b(new_n161), .c(new_n164), .o1(new_n179));
  ao0012aa1n06x5               g084(.a(new_n166), .b(new_n164), .c(new_n167), .o(new_n180));
  aoi112aa1n09x5               g085(.a(new_n180), .b(new_n179), .c(new_n149), .d(new_n178), .o1(new_n181));
  nand02aa1d08x5               g086(.a(new_n177), .b(new_n181), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g088(.a(\a[18] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\a[17] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\b[16] ), .o1(new_n186));
  oaoi03aa1n02x5               g091(.a(new_n185), .b(new_n186), .c(new_n182), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[17] ), .c(new_n184), .out0(\s[18] ));
  xroi22aa1d06x4               g093(.a(new_n185), .b(\b[16] ), .c(new_n184), .d(\b[17] ), .out0(new_n189));
  oai022aa1d24x5               g094(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n190));
  oaib12aa1n18x5               g095(.a(new_n190), .b(new_n184), .c(\b[17] ), .out0(new_n191));
  inv000aa1n06x5               g096(.a(new_n191), .o1(new_n192));
  nor002aa1n20x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nand02aa1d28x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  aoai13aa1n06x5               g100(.a(new_n195), .b(new_n192), .c(new_n182), .d(new_n189), .o1(new_n196));
  aoi112aa1n02x5               g101(.a(new_n195), .b(new_n192), .c(new_n182), .d(new_n189), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n196), .b(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g103(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g104(.a(new_n193), .o1(new_n200));
  nor042aa1n06x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand02aa1d28x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n06x4               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  inv040aa1n03x5               g108(.a(new_n203), .o1(new_n204));
  tech160nm_fiaoi012aa1n03p5x5 g109(.a(new_n204), .b(new_n196), .c(new_n200), .o1(new_n205));
  nona22aa1n02x5               g110(.a(new_n196), .b(new_n203), .c(new_n193), .out0(new_n206));
  norb02aa1n03x4               g111(.a(new_n206), .b(new_n205), .out0(\s[20] ));
  nona23aa1n06x5               g112(.a(new_n189), .b(new_n194), .c(new_n204), .d(new_n193), .out0(new_n208));
  aoi012aa1n12x5               g113(.a(new_n201), .b(new_n193), .c(new_n202), .o1(new_n209));
  nona23aa1d18x5               g114(.a(new_n202), .b(new_n194), .c(new_n193), .d(new_n201), .out0(new_n210));
  oai012aa1d24x5               g115(.a(new_n209), .b(new_n210), .c(new_n191), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n04x5               g117(.a(new_n212), .b(new_n208), .c(new_n177), .d(new_n181), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n04x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  xorc02aa1n02x5               g121(.a(\a[22] ), .b(\b[21] ), .out0(new_n217));
  aoai13aa1n04x5               g122(.a(new_n217), .b(new_n215), .c(new_n213), .d(new_n216), .o1(new_n218));
  aoi112aa1n03x5               g123(.a(new_n215), .b(new_n217), .c(new_n213), .d(new_n216), .o1(new_n219));
  norb02aa1n02x7               g124(.a(new_n218), .b(new_n219), .out0(\s[22] ));
  inv000aa1d42x5               g125(.a(\a[21] ), .o1(new_n221));
  inv040aa1d32x5               g126(.a(\a[22] ), .o1(new_n222));
  xroi22aa1d06x4               g127(.a(new_n221), .b(\b[20] ), .c(new_n222), .d(\b[21] ), .out0(new_n223));
  nanb02aa1n02x5               g128(.a(new_n208), .b(new_n223), .out0(new_n224));
  inv000aa1d42x5               g129(.a(\b[21] ), .o1(new_n225));
  oaoi03aa1n12x5               g130(.a(new_n222), .b(new_n225), .c(new_n215), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoi012aa1n02x5               g132(.a(new_n227), .b(new_n211), .c(new_n223), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n224), .c(new_n177), .d(new_n181), .o1(new_n229));
  xorb03aa1n02x5               g134(.a(new_n229), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g135(.a(\b[22] ), .b(\a[23] ), .o1(new_n231));
  xorc02aa1n02x5               g136(.a(\a[23] ), .b(\b[22] ), .out0(new_n232));
  xorc02aa1n02x5               g137(.a(\a[24] ), .b(\b[23] ), .out0(new_n233));
  aoai13aa1n02x5               g138(.a(new_n233), .b(new_n231), .c(new_n229), .d(new_n232), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n231), .b(new_n233), .c(new_n229), .d(new_n232), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n234), .b(new_n235), .out0(\s[24] ));
  inv040aa1n03x5               g141(.a(new_n209), .o1(new_n237));
  nano23aa1n02x5               g142(.a(new_n193), .b(new_n201), .c(new_n202), .d(new_n194), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n223), .b(new_n237), .c(new_n238), .d(new_n192), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\a[23] ), .o1(new_n240));
  inv040aa1d32x5               g145(.a(\a[24] ), .o1(new_n241));
  xroi22aa1d04x5               g146(.a(new_n240), .b(\b[22] ), .c(new_n241), .d(\b[23] ), .out0(new_n242));
  inv000aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n244));
  aoib12aa1n02x5               g149(.a(new_n244), .b(new_n241), .c(\b[23] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n243), .c(new_n239), .d(new_n226), .o1(new_n246));
  nano22aa1n02x5               g151(.a(new_n208), .b(new_n223), .c(new_n242), .out0(new_n247));
  xorc02aa1n02x5               g152(.a(\a[25] ), .b(\b[24] ), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n246), .c(new_n182), .d(new_n247), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(new_n246), .b(new_n248), .c(new_n182), .d(new_n247), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n249), .b(new_n250), .out0(\s[25] ));
  nor042aa1n03x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  inv000aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  xorc02aa1n02x5               g158(.a(\a[26] ), .b(\b[25] ), .out0(new_n254));
  aobi12aa1n06x5               g159(.a(new_n254), .b(new_n249), .c(new_n253), .out0(new_n255));
  nona22aa1n02x5               g160(.a(new_n249), .b(new_n254), .c(new_n252), .out0(new_n256));
  norb02aa1n03x4               g161(.a(new_n256), .b(new_n255), .out0(\s[26] ));
  inv040aa1d30x5               g162(.a(\a[25] ), .o1(new_n258));
  inv040aa1d32x5               g163(.a(\a[26] ), .o1(new_n259));
  xroi22aa1d06x4               g164(.a(new_n258), .b(\b[24] ), .c(new_n259), .d(\b[25] ), .out0(new_n260));
  nano32aa1n03x7               g165(.a(new_n208), .b(new_n260), .c(new_n223), .d(new_n242), .out0(new_n261));
  nand02aa1d06x5               g166(.a(new_n182), .b(new_n261), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[26] ), .b(\b[25] ), .c(new_n253), .carry(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  tech160nm_fiaoi012aa1n05x5   g169(.a(new_n264), .b(new_n246), .c(new_n260), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[27] ), .b(\b[26] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n265), .c(new_n262), .out0(\s[27] ));
  norp02aa1n02x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  inv040aa1n03x5               g173(.a(new_n268), .o1(new_n269));
  aobi12aa1n06x5               g174(.a(new_n261), .b(new_n177), .c(new_n181), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n242), .b(new_n227), .c(new_n211), .d(new_n223), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n260), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n263), .b(new_n272), .c(new_n271), .d(new_n245), .o1(new_n273));
  oaih12aa1n02x5               g178(.a(new_n266), .b(new_n273), .c(new_n270), .o1(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[27] ), .b(\a[28] ), .out0(new_n275));
  tech160nm_fiaoi012aa1n02p5x5 g180(.a(new_n275), .b(new_n274), .c(new_n269), .o1(new_n276));
  aobi12aa1n06x5               g181(.a(new_n266), .b(new_n265), .c(new_n262), .out0(new_n277));
  nano22aa1n03x5               g182(.a(new_n277), .b(new_n269), .c(new_n275), .out0(new_n278));
  norp02aa1n03x5               g183(.a(new_n276), .b(new_n278), .o1(\s[28] ));
  xnrc02aa1n02x5               g184(.a(\b[28] ), .b(\a[29] ), .out0(new_n280));
  norb02aa1n02x5               g185(.a(new_n266), .b(new_n275), .out0(new_n281));
  oaih12aa1n02x5               g186(.a(new_n281), .b(new_n273), .c(new_n270), .o1(new_n282));
  oao003aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n269), .carry(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n280), .b(new_n282), .c(new_n283), .o1(new_n284));
  aobi12aa1n06x5               g189(.a(new_n281), .b(new_n265), .c(new_n262), .out0(new_n285));
  nano22aa1n03x5               g190(.a(new_n285), .b(new_n280), .c(new_n283), .out0(new_n286));
  norp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n112), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g193(.a(\b[29] ), .b(\a[30] ), .out0(new_n289));
  norb03aa1n02x5               g194(.a(new_n266), .b(new_n280), .c(new_n275), .out0(new_n290));
  oaih12aa1n02x5               g195(.a(new_n290), .b(new_n273), .c(new_n270), .o1(new_n291));
  oao003aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .c(new_n283), .carry(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n289), .b(new_n291), .c(new_n292), .o1(new_n293));
  aobi12aa1n06x5               g198(.a(new_n290), .b(new_n265), .c(new_n262), .out0(new_n294));
  nano22aa1n03x5               g199(.a(new_n294), .b(new_n289), .c(new_n292), .out0(new_n295));
  norp02aa1n03x5               g200(.a(new_n293), .b(new_n295), .o1(\s[30] ));
  norb02aa1n02x5               g201(.a(new_n290), .b(new_n289), .out0(new_n297));
  oaih12aa1n02x5               g202(.a(new_n297), .b(new_n273), .c(new_n270), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n292), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n298), .c(new_n299), .o1(new_n301));
  aobi12aa1n06x5               g206(.a(new_n297), .b(new_n265), .c(new_n262), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n299), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[31] ));
  xnrb03aa1n02x5               g209(.a(new_n114), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g210(.a(\a[3] ), .b(\b[2] ), .c(new_n114), .o1(new_n306));
  xorb03aa1n02x5               g211(.a(new_n306), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g212(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g213(.a(new_n122), .b(new_n121), .c(new_n123), .o1(new_n309));
  xnrb03aa1n02x5               g214(.a(new_n309), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oai012aa1n02x5               g215(.a(new_n107), .b(new_n309), .c(new_n125), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g217(.a(new_n103), .b(new_n311), .c(new_n104), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  aoi112aa1n02x5               g219(.a(new_n110), .b(new_n127), .c(new_n121), .d(new_n126), .o1(new_n315));
  norb02aa1n02x5               g220(.a(new_n128), .b(new_n315), .out0(\s[9] ));
endmodule


