// Benchmark "adder" written by ABC on Wed Jul 17 17:39:23 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n331, new_n332, new_n333,
    new_n335, new_n336, new_n337, new_n339, new_n340;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1d28x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  nor002aa1n16x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  and002aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o(new_n101));
  inv040aa1d32x5               g006(.a(\a[3] ), .o1(new_n102));
  inv030aa1d32x5               g007(.a(\b[2] ), .o1(new_n103));
  nand02aa1n03x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1n02x5               g010(.a(new_n104), .b(new_n105), .o1(new_n106));
  nor042aa1n04x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nand02aa1d08x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nand02aa1n08x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  aoi012aa1d18x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  oa0022aa1n02x5               g015(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n111));
  oaih12aa1n02x5               g016(.a(new_n111), .b(new_n110), .c(new_n106), .o1(new_n112));
  nor042aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor022aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n03x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nor042aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nand42aa1n10x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor042aa1n04x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nand42aa1n06x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nano23aa1n06x5               g026(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n122));
  nona23aa1n09x5               g027(.a(new_n112), .b(new_n122), .c(new_n117), .d(new_n101), .out0(new_n123));
  aoi012aa1n02x5               g028(.a(new_n118), .b(new_n120), .c(new_n119), .o1(new_n124));
  ao0012aa1n03x5               g029(.a(new_n113), .b(new_n115), .c(new_n114), .o(new_n125));
  oab012aa1n06x5               g030(.a(new_n125), .b(new_n117), .c(new_n124), .out0(new_n126));
  nand22aa1n03x5               g031(.a(new_n123), .b(new_n126), .o1(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoi012aa1n02x5               g033(.a(new_n100), .b(new_n127), .c(new_n128), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n98), .c(new_n99), .out0(\s[10] ));
  nanp02aa1n09x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nano23aa1d15x5               g036(.a(new_n97), .b(new_n100), .c(new_n131), .d(new_n99), .out0(new_n132));
  aoi012aa1d24x5               g037(.a(new_n97), .b(new_n100), .c(new_n99), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand42aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n12x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  aoai13aa1n06x5               g042(.a(new_n137), .b(new_n134), .c(new_n127), .d(new_n132), .o1(new_n138));
  aoi112aa1n02x5               g043(.a(new_n137), .b(new_n134), .c(new_n127), .d(new_n132), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n138), .b(new_n139), .out0(\s[11] ));
  inv000aa1d42x5               g045(.a(new_n135), .o1(new_n141));
  nor002aa1d32x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d08x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n09x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n138), .c(new_n141), .out0(\s[12] ));
  nona23aa1d18x5               g050(.a(new_n143), .b(new_n136), .c(new_n135), .d(new_n142), .out0(new_n146));
  aoi012aa1d18x5               g051(.a(new_n142), .b(new_n135), .c(new_n143), .o1(new_n147));
  oai012aa1d24x5               g052(.a(new_n147), .b(new_n146), .c(new_n133), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nand23aa1d12x5               g054(.a(new_n132), .b(new_n137), .c(new_n144), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n149), .b(new_n150), .c(new_n123), .d(new_n126), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n16x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  tech160nm_finand02aa1n05x5   g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n03x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  oaoi13aa1n12x5               g061(.a(new_n101), .b(new_n111), .c(new_n110), .d(new_n106), .o1(new_n157));
  norb02aa1n02x7               g062(.a(new_n122), .b(new_n117), .out0(new_n158));
  oabi12aa1n03x5               g063(.a(new_n125), .b(new_n117), .c(new_n124), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n150), .o1(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n159), .c(new_n157), .d(new_n158), .o1(new_n161));
  nor002aa1d32x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand02aa1d16x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  aoi012aa1d18x5               g068(.a(new_n162), .b(new_n153), .c(new_n163), .o1(new_n164));
  nona23aa1n03x5               g069(.a(new_n163), .b(new_n154), .c(new_n153), .d(new_n162), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n164), .b(new_n165), .c(new_n161), .d(new_n149), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  norb02aa1n02x7               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  nor042aa1n06x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nanp02aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n12x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(new_n173), .b(new_n168), .c(new_n166), .d(new_n170), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n168), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n164), .o1(new_n176));
  nano23aa1d12x5               g081(.a(new_n153), .b(new_n162), .c(new_n163), .d(new_n154), .out0(new_n177));
  aoai13aa1n02x5               g082(.a(new_n170), .b(new_n176), .c(new_n151), .d(new_n177), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n173), .o1(new_n179));
  tech160nm_fiaoi012aa1n02p5x5 g084(.a(new_n179), .b(new_n178), .c(new_n175), .o1(new_n180));
  norp02aa1n02x5               g085(.a(new_n180), .b(new_n174), .o1(\s[16] ));
  nona23aa1n09x5               g086(.a(new_n172), .b(new_n169), .c(new_n168), .d(new_n171), .out0(new_n182));
  nona23aa1d18x5               g087(.a(new_n132), .b(new_n177), .c(new_n182), .d(new_n146), .out0(new_n183));
  nor002aa1n03x5               g088(.a(new_n182), .b(new_n165), .o1(new_n184));
  aoi012aa1n02x7               g089(.a(new_n171), .b(new_n168), .c(new_n172), .o1(new_n185));
  tech160nm_fioai012aa1n04x5   g090(.a(new_n185), .b(new_n182), .c(new_n164), .o1(new_n186));
  aoi012aa1d24x5               g091(.a(new_n186), .b(new_n148), .c(new_n184), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n183), .c(new_n123), .d(new_n126), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1n06x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nanp02aa1n04x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  tech160nm_fiaoi012aa1n05x5   g096(.a(new_n190), .b(new_n188), .c(new_n191), .o1(new_n192));
  xnrb03aa1n03x5               g097(.a(new_n192), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nano32aa1n03x7               g098(.a(new_n150), .b(new_n173), .c(new_n170), .d(new_n177), .out0(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n159), .c(new_n157), .d(new_n158), .o1(new_n195));
  norp02aa1n09x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nand02aa1d10x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nano23aa1n06x5               g102(.a(new_n190), .b(new_n196), .c(new_n197), .d(new_n191), .out0(new_n198));
  inv040aa1n08x5               g103(.a(new_n198), .o1(new_n199));
  aoi012aa1d18x5               g104(.a(new_n196), .b(new_n190), .c(new_n197), .o1(new_n200));
  aoai13aa1n02x7               g105(.a(new_n200), .b(new_n199), .c(new_n195), .d(new_n187), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  xorc02aa1n12x5               g109(.a(\a[19] ), .b(\b[18] ), .out0(new_n205));
  nor042aa1n04x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nand02aa1d16x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  norb02aa1n03x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  aoi112aa1n03x4               g113(.a(new_n204), .b(new_n208), .c(new_n201), .d(new_n205), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n204), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n200), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n205), .b(new_n211), .c(new_n188), .d(new_n198), .o1(new_n212));
  nanb02aa1n06x5               g117(.a(new_n206), .b(new_n207), .out0(new_n213));
  aoi012aa1n03x5               g118(.a(new_n213), .b(new_n212), .c(new_n210), .o1(new_n214));
  norp02aa1n03x5               g119(.a(new_n214), .b(new_n209), .o1(\s[20] ));
  nano22aa1n12x5               g120(.a(new_n199), .b(new_n205), .c(new_n208), .out0(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  tech160nm_fixnrc02aa1n04x5   g122(.a(\b[18] ), .b(\a[19] ), .out0(new_n218));
  aoi012aa1n09x5               g123(.a(new_n206), .b(new_n204), .c(new_n207), .o1(new_n219));
  oai013aa1d12x5               g124(.a(new_n219), .b(new_n218), .c(new_n200), .d(new_n213), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n04x5               g126(.a(new_n221), .b(new_n217), .c(new_n195), .d(new_n187), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  nand02aa1d06x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  norb02aa1n02x5               g130(.a(new_n225), .b(new_n224), .out0(new_n226));
  nor042aa1n04x5               g131(.a(\b[21] ), .b(\a[22] ), .o1(new_n227));
  nand22aa1n04x5               g132(.a(\b[21] ), .b(\a[22] ), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  aoi112aa1n02x5               g134(.a(new_n224), .b(new_n229), .c(new_n222), .d(new_n226), .o1(new_n230));
  inv040aa1n12x5               g135(.a(new_n224), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n226), .b(new_n220), .c(new_n188), .d(new_n216), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n229), .o1(new_n233));
  aoi012aa1n03x5               g138(.a(new_n233), .b(new_n232), .c(new_n231), .o1(new_n234));
  norp02aa1n03x5               g139(.a(new_n234), .b(new_n230), .o1(\s[22] ));
  nano23aa1d15x5               g140(.a(new_n224), .b(new_n227), .c(new_n228), .d(new_n225), .out0(new_n236));
  nano32aa1n02x4               g141(.a(new_n199), .b(new_n236), .c(new_n205), .d(new_n208), .out0(new_n237));
  inv000aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  oaoi03aa1n12x5               g143(.a(\a[22] ), .b(\b[21] ), .c(new_n231), .o1(new_n239));
  aoi012aa1d24x5               g144(.a(new_n239), .b(new_n220), .c(new_n236), .o1(new_n240));
  aoai13aa1n04x5               g145(.a(new_n240), .b(new_n238), .c(new_n195), .d(new_n187), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1d32x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  nand42aa1n06x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  nor022aa1n08x5               g150(.a(\b[23] ), .b(\a[24] ), .o1(new_n246));
  nand42aa1n04x5               g151(.a(\b[23] ), .b(\a[24] ), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  aoi112aa1n02x5               g153(.a(new_n243), .b(new_n248), .c(new_n241), .d(new_n245), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n243), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n240), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n245), .b(new_n251), .c(new_n188), .d(new_n237), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n248), .o1(new_n253));
  aoi012aa1n03x5               g158(.a(new_n253), .b(new_n252), .c(new_n250), .o1(new_n254));
  norp02aa1n03x5               g159(.a(new_n254), .b(new_n249), .o1(\s[24] ));
  nona23aa1n03x5               g160(.a(new_n228), .b(new_n225), .c(new_n224), .d(new_n227), .out0(new_n256));
  nona23aa1n02x4               g161(.a(new_n247), .b(new_n244), .c(new_n243), .d(new_n246), .out0(new_n257));
  nona22aa1d18x5               g162(.a(new_n216), .b(new_n256), .c(new_n257), .out0(new_n258));
  aoi112aa1n03x5               g163(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n259));
  oai112aa1n04x5               g164(.a(new_n205), .b(new_n208), .c(new_n259), .d(new_n196), .o1(new_n260));
  nano23aa1n09x5               g165(.a(new_n243), .b(new_n246), .c(new_n247), .d(new_n244), .out0(new_n261));
  nand22aa1n03x5               g166(.a(new_n261), .b(new_n236), .o1(new_n262));
  oaoi03aa1n09x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n250), .o1(new_n263));
  aoi012aa1n12x5               g168(.a(new_n263), .b(new_n261), .c(new_n239), .o1(new_n264));
  aoai13aa1n12x5               g169(.a(new_n264), .b(new_n262), .c(new_n260), .d(new_n219), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  aoai13aa1n02x7               g171(.a(new_n266), .b(new_n258), .c(new_n195), .d(new_n187), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xorc02aa1n12x5               g175(.a(\a[26] ), .b(\b[25] ), .out0(new_n271));
  aoi112aa1n03x4               g176(.a(new_n269), .b(new_n271), .c(new_n267), .d(new_n270), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n269), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n258), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n270), .b(new_n265), .c(new_n188), .d(new_n274), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n271), .o1(new_n276));
  aoi012aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n273), .o1(new_n277));
  nor002aa1n02x5               g182(.a(new_n277), .b(new_n272), .o1(\s[26] ));
  nand02aa1d06x5               g183(.a(new_n271), .b(new_n270), .o1(new_n279));
  nona32aa1n02x4               g184(.a(new_n216), .b(new_n279), .c(new_n257), .d(new_n256), .out0(new_n280));
  inv000aa1d42x5               g185(.a(new_n279), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[26] ), .b(\b[25] ), .c(new_n273), .carry(new_n282));
  aobi12aa1n06x5               g187(.a(new_n282), .b(new_n265), .c(new_n281), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n280), .c(new_n195), .d(new_n187), .o1(new_n284));
  xorb03aa1n03x5               g189(.a(new_n284), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  inv000aa1n03x5               g191(.a(new_n286), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .out0(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  inv040aa1n03x5               g194(.a(new_n280), .o1(new_n290));
  nor002aa1n02x5               g195(.a(new_n257), .b(new_n256), .o1(new_n291));
  nand22aa1n03x5               g196(.a(new_n220), .b(new_n291), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n282), .b(new_n279), .c(new_n292), .d(new_n264), .o1(new_n293));
  nanp02aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  aoai13aa1n02x7               g199(.a(new_n294), .b(new_n293), .c(new_n188), .d(new_n290), .o1(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n289), .b(new_n295), .c(new_n287), .o1(new_n296));
  aoi112aa1n03x4               g201(.a(new_n286), .b(new_n288), .c(new_n284), .d(new_n294), .o1(new_n297));
  norp02aa1n03x5               g202(.a(new_n296), .b(new_n297), .o1(\s[28] ));
  nano22aa1n02x4               g203(.a(new_n289), .b(new_n287), .c(new_n294), .out0(new_n299));
  aoai13aa1n02x7               g204(.a(new_n299), .b(new_n293), .c(new_n188), .d(new_n290), .o1(new_n300));
  oaoi03aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .o1(new_n301));
  inv000aa1n03x5               g206(.a(new_n301), .o1(new_n302));
  xorc02aa1n12x5               g207(.a(\a[29] ), .b(\b[28] ), .out0(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  tech160nm_fiaoi012aa1n02p5x5 g209(.a(new_n304), .b(new_n300), .c(new_n302), .o1(new_n305));
  aoi112aa1n03x4               g210(.a(new_n303), .b(new_n301), .c(new_n284), .d(new_n299), .o1(new_n306));
  norp02aa1n03x5               g211(.a(new_n305), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g213(.a(new_n304), .b(new_n288), .c(new_n294), .d(new_n287), .out0(new_n309));
  aoai13aa1n02x7               g214(.a(new_n309), .b(new_n293), .c(new_n188), .d(new_n290), .o1(new_n310));
  oao003aa1n09x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n302), .carry(new_n311));
  tech160nm_fixorc02aa1n03p5x5 g216(.a(\a[30] ), .b(\b[29] ), .out0(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n313), .b(new_n310), .c(new_n311), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n311), .o1(new_n315));
  aoi112aa1n03x4               g220(.a(new_n312), .b(new_n315), .c(new_n284), .d(new_n309), .o1(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[30] ));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  inv000aa1d42x5               g223(.a(new_n318), .o1(new_n319));
  and003aa1n02x5               g224(.a(new_n299), .b(new_n312), .c(new_n303), .o(new_n320));
  tech160nm_fioaoi03aa1n03p5x5 g225(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .o1(new_n321));
  aoi112aa1n02x7               g226(.a(new_n319), .b(new_n321), .c(new_n284), .d(new_n320), .o1(new_n322));
  aoai13aa1n02x7               g227(.a(new_n320), .b(new_n293), .c(new_n188), .d(new_n290), .o1(new_n323));
  inv000aa1n02x5               g228(.a(new_n321), .o1(new_n324));
  aoi012aa1n03x5               g229(.a(new_n318), .b(new_n323), .c(new_n324), .o1(new_n325));
  nor002aa1n02x5               g230(.a(new_n325), .b(new_n322), .o1(\s[31] ));
  xnbna2aa1n03x5               g231(.a(new_n110), .b(new_n104), .c(new_n105), .out0(\s[3] ));
  oaoi03aa1n02x5               g232(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g234(.a(new_n157), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g235(.a(new_n119), .b(new_n118), .out0(new_n331));
  oai112aa1n06x5               g236(.a(new_n121), .b(new_n331), .c(new_n157), .d(new_n120), .o1(new_n332));
  oaoi13aa1n02x5               g237(.a(new_n331), .b(new_n121), .c(new_n157), .d(new_n120), .o1(new_n333));
  norb02aa1n02x5               g238(.a(new_n332), .b(new_n333), .out0(\s[6] ));
  nanb02aa1n02x5               g239(.a(new_n115), .b(new_n116), .out0(new_n335));
  oaoi13aa1n04x5               g240(.a(new_n335), .b(new_n332), .c(\a[6] ), .d(\b[5] ), .o1(new_n336));
  oai112aa1n02x5               g241(.a(new_n332), .b(new_n335), .c(\b[5] ), .d(\a[6] ), .o1(new_n337));
  norb02aa1n02x5               g242(.a(new_n337), .b(new_n336), .out0(\s[7] ));
  orn002aa1n02x5               g243(.a(\a[8] ), .b(\b[7] ), .o(new_n339));
  nor042aa1n03x5               g244(.a(new_n336), .b(new_n115), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n340), .b(new_n339), .c(new_n114), .out0(\s[8] ));
  xnbna2aa1n03x5               g246(.a(new_n128), .b(new_n123), .c(new_n126), .out0(\s[9] ));
endmodule


