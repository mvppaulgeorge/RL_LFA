// Benchmark "adder" written by ABC on Wed Jul 17 17:04:51 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n317,
    new_n320, new_n321, new_n323, new_n325, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[8] ), .o1(new_n97));
  nanb02aa1d36x5               g002(.a(\a[9] ), .b(new_n97), .out0(new_n98));
  nor002aa1d32x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand02aa1d06x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  aoi012aa1n02x5               g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  oaih22aa1n04x5               g007(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n103));
  and002aa1n12x5               g008(.a(\b[5] ), .b(\a[6] ), .o(new_n104));
  nand02aa1d06x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  inv000aa1n02x5               g010(.a(new_n105), .o1(new_n106));
  norb03aa1n03x5               g011(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n107));
  nona23aa1n03x5               g012(.a(new_n107), .b(new_n103), .c(new_n104), .d(new_n106), .out0(new_n108));
  nand22aa1n03x5               g013(.a(new_n108), .b(new_n102), .o1(new_n109));
  norp02aa1n03x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nor022aa1n16x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  aoi012aa1n02x7               g017(.a(new_n110), .b(new_n112), .c(new_n111), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[0] ), .b(\a[1] ), .o1(new_n115));
  nor002aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  tech160nm_fioai012aa1n04x5   g021(.a(new_n114), .b(new_n116), .c(new_n115), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[2] ), .b(\a[3] ), .o1(new_n118));
  nona23aa1n06x5               g023(.a(new_n118), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n119));
  oai012aa1n12x5               g024(.a(new_n113), .b(new_n119), .c(new_n117), .o1(new_n120));
  nona23aa1d18x5               g025(.a(new_n105), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n121));
  xnrc02aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .out0(new_n122));
  xnrc02aa1n02x5               g027(.a(\b[5] ), .b(\a[6] ), .out0(new_n123));
  nor043aa1n06x5               g028(.a(new_n121), .b(new_n122), .c(new_n123), .o1(new_n124));
  nand22aa1n09x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nand22aa1n12x5               g030(.a(new_n98), .b(new_n125), .o1(new_n126));
  inv000aa1d42x5               g031(.a(new_n126), .o1(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n109), .c(new_n120), .d(new_n124), .o1(new_n128));
  nor002aa1d32x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1n06x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1d24x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  aoi112aa1n09x5               g038(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n134));
  norp02aa1n02x5               g039(.a(new_n134), .b(new_n129), .o1(new_n135));
  aoai13aa1n06x5               g040(.a(new_n135), .b(new_n128), .c(\a[10] ), .d(\b[9] ), .o1(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nand02aa1d28x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nor002aa1n12x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nor042aa1d18x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n06x4               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  aoi112aa1n02x5               g047(.a(new_n142), .b(new_n139), .c(new_n136), .d(new_n138), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n142), .b(new_n139), .c(new_n136), .d(new_n138), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(\s[12] ));
  inv000aa1d42x5               g050(.a(new_n104), .o1(new_n146));
  nano22aa1n02x4               g051(.a(new_n121), .b(new_n103), .c(new_n146), .out0(new_n147));
  norb02aa1n03x5               g052(.a(new_n102), .b(new_n147), .out0(new_n148));
  nanp02aa1n03x5               g053(.a(new_n120), .b(new_n124), .o1(new_n149));
  nano23aa1d15x5               g054(.a(new_n140), .b(new_n139), .c(new_n141), .d(new_n138), .out0(new_n150));
  nona22aa1d36x5               g055(.a(new_n150), .b(new_n131), .c(new_n126), .out0(new_n151));
  aoi112aa1n02x7               g056(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n152));
  norb02aa1n06x4               g057(.a(new_n138), .b(new_n139), .out0(new_n153));
  oai112aa1n06x5               g058(.a(new_n142), .b(new_n153), .c(new_n134), .d(new_n129), .o1(new_n154));
  nona22aa1d24x5               g059(.a(new_n154), .b(new_n152), .c(new_n140), .out0(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n151), .c(new_n149), .d(new_n148), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nand42aa1n03x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nor002aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n160), .b(new_n157), .c(new_n159), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g067(.a(new_n151), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n109), .c(new_n120), .d(new_n124), .o1(new_n164));
  nor022aa1n04x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand22aa1n04x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n165), .b(new_n160), .c(new_n166), .o1(new_n167));
  nona23aa1n03x5               g072(.a(new_n159), .b(new_n166), .c(new_n165), .d(new_n160), .out0(new_n168));
  aoai13aa1n06x5               g073(.a(new_n167), .b(new_n168), .c(new_n164), .d(new_n156), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand42aa1n08x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nor002aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norp02aa1n12x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand02aa1d12x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanb02aa1n18x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  aoi112aa1n02x5               g081(.a(new_n176), .b(new_n172), .c(new_n169), .d(new_n171), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n176), .b(new_n172), .c(new_n169), .d(new_n171), .o1(new_n178));
  norb02aa1n03x4               g083(.a(new_n178), .b(new_n177), .out0(\s[16] ));
  xorc02aa1n12x5               g084(.a(\a[17] ), .b(\b[16] ), .out0(new_n180));
  nano23aa1n03x5               g085(.a(new_n165), .b(new_n160), .c(new_n166), .d(new_n159), .out0(new_n181));
  nano23aa1n02x4               g086(.a(new_n173), .b(new_n172), .c(new_n174), .d(new_n171), .out0(new_n182));
  nanp02aa1n03x5               g087(.a(new_n182), .b(new_n181), .o1(new_n183));
  nor042aa1n12x5               g088(.a(new_n151), .b(new_n183), .o1(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n109), .c(new_n120), .d(new_n124), .o1(new_n185));
  nanb02aa1n02x5               g090(.a(new_n172), .b(new_n171), .out0(new_n186));
  nor043aa1n02x5               g091(.a(new_n168), .b(new_n175), .c(new_n186), .o1(new_n187));
  nor003aa1n03x5               g092(.a(new_n167), .b(new_n175), .c(new_n186), .o1(new_n188));
  tech160nm_fiao0012aa1n02p5x5 g093(.a(new_n173), .b(new_n172), .c(new_n174), .o(new_n189));
  aoi112aa1n09x5               g094(.a(new_n189), .b(new_n188), .c(new_n155), .d(new_n187), .o1(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n180), .b(new_n190), .c(new_n185), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[18] ), .o1(new_n192));
  norp02aa1n02x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  nand02aa1d06x5               g098(.a(new_n190), .b(new_n185), .o1(new_n194));
  tech160nm_fiaoi012aa1n05x5   g099(.a(new_n193), .b(new_n194), .c(new_n180), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xorc02aa1n02x5               g101(.a(\a[18] ), .b(\b[17] ), .out0(new_n197));
  and002aa1n02x5               g102(.a(new_n197), .b(new_n180), .o(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\b[17] ), .o1(new_n200));
  oao003aa1n02x5               g105(.a(new_n192), .b(new_n200), .c(new_n193), .carry(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n185), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n09x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nor042aa1n03x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1n08x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n06x4               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi112aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n203), .d(new_n206), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n210), .b(new_n207), .c(new_n203), .d(new_n206), .o1(new_n212));
  norb02aa1n03x4               g117(.a(new_n212), .b(new_n211), .out0(\s[20] ));
  nano23aa1n02x4               g118(.a(new_n208), .b(new_n207), .c(new_n209), .d(new_n206), .out0(new_n214));
  nanp03aa1n02x5               g119(.a(new_n214), .b(new_n180), .c(new_n197), .o1(new_n215));
  aoi112aa1n02x5               g120(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n216));
  norp02aa1n02x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  aoi112aa1n03x5               g122(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n218));
  norb02aa1n03x4               g123(.a(new_n206), .b(new_n207), .out0(new_n219));
  oai112aa1n06x5               g124(.a(new_n219), .b(new_n210), .c(new_n218), .d(new_n217), .o1(new_n220));
  nona22aa1d18x5               g125(.a(new_n220), .b(new_n216), .c(new_n208), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n215), .c(new_n190), .d(new_n185), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoi112aa1n03x5               g134(.a(new_n225), .b(new_n229), .c(new_n223), .d(new_n227), .o1(new_n230));
  aoai13aa1n03x5               g135(.a(new_n229), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n231));
  norb02aa1n03x4               g136(.a(new_n231), .b(new_n230), .out0(\s[22] ));
  nor042aa1n02x5               g137(.a(new_n228), .b(new_n226), .o1(new_n233));
  nand03aa1n02x5               g138(.a(new_n198), .b(new_n214), .c(new_n233), .o1(new_n234));
  inv000aa1n02x5               g139(.a(new_n225), .o1(new_n235));
  oaoi03aa1n02x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n221), .c(new_n233), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n234), .c(new_n190), .d(new_n185), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n04x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  nand22aa1n03x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  nor002aa1n06x5               g146(.a(\b[23] ), .b(\a[24] ), .o1(new_n242));
  nanp02aa1n02x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n243), .b(new_n242), .out0(new_n244));
  aoi112aa1n03x5               g149(.a(new_n240), .b(new_n244), .c(new_n238), .d(new_n241), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n244), .b(new_n240), .c(new_n238), .d(new_n241), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n246), .b(new_n245), .out0(\s[24] ));
  nona23aa1n03x5               g152(.a(new_n243), .b(new_n241), .c(new_n240), .d(new_n242), .out0(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  nano22aa1n02x4               g154(.a(new_n215), .b(new_n249), .c(new_n233), .out0(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  nona32aa1n09x5               g156(.a(new_n221), .b(new_n248), .c(new_n228), .d(new_n226), .out0(new_n252));
  aoi112aa1n02x5               g157(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n253));
  aoi112aa1n03x5               g158(.a(new_n253), .b(new_n242), .c(new_n249), .d(new_n236), .o1(new_n254));
  nanp02aa1n06x5               g159(.a(new_n252), .b(new_n254), .o1(new_n255));
  inv040aa1n06x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n251), .c(new_n190), .d(new_n185), .o1(new_n257));
  xorb03aa1n02x5               g162(.a(new_n257), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  tech160nm_fixorc02aa1n04x5   g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  tech160nm_fixorc02aa1n04x5   g165(.a(\a[26] ), .b(\b[25] ), .out0(new_n261));
  aoi112aa1n02x7               g166(.a(new_n259), .b(new_n261), .c(new_n257), .d(new_n260), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n261), .b(new_n259), .c(new_n257), .d(new_n260), .o1(new_n263));
  norb02aa1n02x7               g168(.a(new_n263), .b(new_n262), .out0(\s[26] ));
  nanp02aa1n03x5               g169(.a(new_n149), .b(new_n148), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(new_n155), .b(new_n187), .o1(new_n266));
  nona22aa1n02x4               g171(.a(new_n266), .b(new_n189), .c(new_n188), .out0(new_n267));
  and002aa1n12x5               g172(.a(new_n261), .b(new_n260), .o(new_n268));
  nano32aa1n03x7               g173(.a(new_n215), .b(new_n268), .c(new_n233), .d(new_n249), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n267), .c(new_n265), .d(new_n184), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n259), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  aoi012aa1n12x5               g178(.a(new_n273), .b(new_n255), .c(new_n268), .o1(new_n274));
  xorc02aa1n12x5               g179(.a(\a[27] ), .b(\b[26] ), .out0(new_n275));
  xnbna2aa1n03x5               g180(.a(new_n275), .b(new_n270), .c(new_n274), .out0(\s[27] ));
  norp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  inv040aa1n03x5               g182(.a(new_n277), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n275), .o1(new_n279));
  tech160nm_fiaoi012aa1n02p5x5 g184(.a(new_n279), .b(new_n270), .c(new_n274), .o1(new_n280));
  xnrc02aa1n12x5               g185(.a(\b[27] ), .b(\a[28] ), .out0(new_n281));
  nano22aa1n03x5               g186(.a(new_n280), .b(new_n278), .c(new_n281), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n268), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n272), .b(new_n283), .c(new_n252), .d(new_n254), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n275), .b(new_n284), .c(new_n194), .d(new_n269), .o1(new_n285));
  tech160nm_fiaoi012aa1n02p5x5 g190(.a(new_n281), .b(new_n285), .c(new_n278), .o1(new_n286));
  norp02aa1n03x5               g191(.a(new_n286), .b(new_n282), .o1(\s[28] ));
  norb02aa1d21x5               g192(.a(new_n275), .b(new_n281), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n284), .c(new_n194), .d(new_n269), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n278), .carry(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  aoi012aa1n02x7               g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n288), .o1(new_n293));
  aoi012aa1n02x7               g198(.a(new_n293), .b(new_n270), .c(new_n274), .o1(new_n294));
  nano22aa1n03x5               g199(.a(new_n294), .b(new_n290), .c(new_n291), .out0(new_n295));
  norp02aa1n03x5               g200(.a(new_n292), .b(new_n295), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n115), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g202(.a(new_n275), .b(new_n291), .c(new_n281), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n284), .c(new_n194), .d(new_n269), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[29] ), .b(\a[30] ), .out0(new_n301));
  tech160nm_fiaoi012aa1n02p5x5 g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n298), .o1(new_n303));
  tech160nm_fiaoi012aa1n03p5x5 g208(.a(new_n303), .b(new_n270), .c(new_n274), .o1(new_n304));
  nano22aa1n03x7               g209(.a(new_n304), .b(new_n300), .c(new_n301), .out0(new_n305));
  norp02aa1n03x5               g210(.a(new_n302), .b(new_n305), .o1(\s[30] ));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  norb02aa1n03x4               g212(.a(new_n298), .b(new_n301), .out0(new_n308));
  inv020aa1n02x5               g213(.a(new_n308), .o1(new_n309));
  aoi012aa1n06x5               g214(.a(new_n309), .b(new_n270), .c(new_n274), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n311));
  nano22aa1n03x5               g216(.a(new_n310), .b(new_n307), .c(new_n311), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n308), .b(new_n284), .c(new_n194), .d(new_n269), .o1(new_n313));
  aoi012aa1n03x5               g218(.a(new_n307), .b(new_n313), .c(new_n311), .o1(new_n314));
  nor002aa1n02x5               g219(.a(new_n314), .b(new_n312), .o1(\s[31] ));
  xnrb03aa1n02x5               g220(.a(new_n117), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g221(.a(\a[3] ), .b(\b[2] ), .c(new_n117), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g223(.a(new_n120), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanp02aa1n02x5               g224(.a(\b[4] ), .b(\a[5] ), .o1(new_n320));
  tech160nm_fioai012aa1n05x5   g225(.a(new_n320), .b(new_n120), .c(new_n122), .o1(new_n321));
  xnrb03aa1n02x5               g226(.a(new_n321), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g227(.a(\a[6] ), .b(\b[5] ), .c(new_n321), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  inv000aa1d42x5               g229(.a(new_n99), .o1(new_n325));
  tech160nm_fiaoi012aa1n05x5   g230(.a(new_n101), .b(new_n323), .c(new_n105), .o1(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n326), .b(new_n325), .c(new_n100), .out0(\s[8] ));
  xnbna2aa1n03x5               g232(.a(new_n127), .b(new_n149), .c(new_n148), .out0(\s[9] ));
endmodule


