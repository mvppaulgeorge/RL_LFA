// Benchmark "adder" written by ABC on Thu Jul 18 03:31:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n323,
    new_n325, new_n326, new_n329, new_n331, new_n333;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nand02aa1d24x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n09x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor042aa1n09x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  norb03aa1n02x5               g007(.a(new_n101), .b(new_n100), .c(new_n102), .out0(new_n103));
  nor002aa1n20x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb03aa1n02x5               g010(.a(new_n104), .b(new_n105), .c(new_n101), .out0(new_n106));
  oab012aa1n03x5               g011(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .out0(new_n107));
  oai012aa1n02x5               g012(.a(new_n107), .b(new_n103), .c(new_n106), .o1(new_n108));
  nor042aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nanp02aa1n12x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nor042aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n08x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nona23aa1n02x4               g017(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[5] ), .b(\a[6] ), .out0(new_n114));
  tech160nm_fixnrc02aa1n02p5x5 g019(.a(\b[4] ), .b(\a[5] ), .out0(new_n115));
  nor043aa1n03x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nand23aa1n03x5               g021(.a(new_n116), .b(new_n108), .c(new_n99), .o1(new_n117));
  nano23aa1n09x5               g022(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n118));
  oa0012aa1n03x5               g023(.a(new_n110), .b(new_n111), .c(new_n109), .o(new_n119));
  inv000aa1d42x5               g024(.a(\a[5] ), .o1(new_n120));
  nanb02aa1n12x5               g025(.a(\b[4] ), .b(new_n120), .out0(new_n121));
  oaoi03aa1n06x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  aoi012aa1n12x5               g027(.a(new_n119), .b(new_n118), .c(new_n122), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nanb02aa1n02x5               g029(.a(new_n97), .b(new_n124), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n98), .b(new_n125), .c(new_n117), .d(new_n123), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1n04x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanb02aa1n09x5               g034(.a(new_n128), .b(new_n129), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  nona22aa1n02x5               g036(.a(new_n101), .b(new_n102), .c(new_n100), .out0(new_n132));
  nano22aa1n03x7               g037(.a(new_n104), .b(new_n101), .c(new_n105), .out0(new_n133));
  inv030aa1n02x5               g038(.a(new_n107), .o1(new_n134));
  aoai13aa1n12x5               g039(.a(new_n99), .b(new_n134), .c(new_n133), .d(new_n132), .o1(new_n135));
  nona22aa1n02x4               g040(.a(new_n118), .b(new_n114), .c(new_n115), .out0(new_n136));
  oai012aa1n02x5               g041(.a(new_n123), .b(new_n135), .c(new_n136), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n131), .b(new_n97), .c(new_n137), .d(new_n124), .o1(new_n138));
  tech160nm_fioai012aa1n05x5   g043(.a(new_n129), .b(new_n97), .c(new_n128), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nand22aa1n06x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n139), .out0(\s[11] ));
  inv000aa1d42x5               g048(.a(new_n140), .o1(new_n144));
  inv030aa1n02x5               g049(.a(new_n139), .o1(new_n145));
  aoai13aa1n02x5               g050(.a(new_n142), .b(new_n145), .c(new_n126), .d(new_n131), .o1(new_n146));
  nor022aa1n16x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  tech160nm_finand02aa1n05x5   g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  aobi12aa1n06x5               g054(.a(new_n149), .b(new_n146), .c(new_n144), .out0(new_n150));
  nona22aa1n02x4               g055(.a(new_n146), .b(new_n149), .c(new_n140), .out0(new_n151));
  norb02aa1n03x4               g056(.a(new_n151), .b(new_n150), .out0(\s[12] ));
  nano23aa1n03x7               g057(.a(new_n140), .b(new_n147), .c(new_n148), .d(new_n141), .out0(new_n153));
  nona22aa1n03x5               g058(.a(new_n153), .b(new_n130), .c(new_n125), .out0(new_n154));
  nona23aa1d18x5               g059(.a(new_n148), .b(new_n141), .c(new_n140), .d(new_n147), .out0(new_n155));
  oaoi03aa1n06x5               g060(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n156));
  oabi12aa1n12x5               g061(.a(new_n156), .b(new_n155), .c(new_n139), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n154), .c(new_n117), .d(new_n123), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nand42aa1n06x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  aoi012aa1n02x5               g067(.a(new_n161), .b(new_n159), .c(new_n162), .o1(new_n163));
  xnrb03aa1n02x5               g068(.a(new_n163), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand42aa1n06x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nano23aa1d15x5               g071(.a(new_n161), .b(new_n165), .c(new_n166), .d(new_n162), .out0(new_n167));
  oai012aa1n12x5               g072(.a(new_n166), .b(new_n165), .c(new_n161), .o1(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand42aa1d28x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  aoai13aa1n04x5               g078(.a(new_n173), .b(new_n169), .c(new_n159), .d(new_n167), .o1(new_n174));
  aoi112aa1n02x5               g079(.a(new_n173), .b(new_n169), .c(new_n159), .d(new_n167), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n174), .b(new_n175), .out0(\s[15] ));
  nor002aa1n03x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand42aa1n20x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  oaoi13aa1n06x5               g084(.a(new_n179), .b(new_n174), .c(\a[15] ), .d(\b[14] ), .o1(new_n180));
  oai112aa1n02x5               g085(.a(new_n174), .b(new_n179), .c(\b[14] ), .d(\a[15] ), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n181), .b(new_n180), .out0(\s[16] ));
  nona23aa1n02x5               g087(.a(new_n124), .b(new_n129), .c(new_n128), .d(new_n97), .out0(new_n183));
  nano23aa1d12x5               g088(.a(new_n170), .b(new_n177), .c(new_n178), .d(new_n171), .out0(new_n184));
  nona23aa1n09x5               g089(.a(new_n167), .b(new_n184), .c(new_n183), .d(new_n155), .out0(new_n185));
  oaoi13aa1n12x5               g090(.a(new_n185), .b(new_n123), .c(new_n135), .d(new_n136), .o1(new_n186));
  inv040aa1n03x5               g091(.a(new_n184), .o1(new_n187));
  aoai13aa1n04x5               g092(.a(new_n167), .b(new_n156), .c(new_n153), .d(new_n145), .o1(new_n188));
  aoi012aa1n02x5               g093(.a(new_n177), .b(new_n170), .c(new_n178), .o1(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n187), .c(new_n188), .d(new_n168), .o1(new_n190));
  nor042aa1n06x5               g095(.a(new_n190), .b(new_n186), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[16] ), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(new_n193), .b(new_n192), .o1(new_n194));
  nanp02aa1n02x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n191), .b(new_n195), .c(new_n194), .out0(\s[17] ));
  norp02aa1n12x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nanp02aa1n09x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nanb02aa1n06x5               g103(.a(new_n197), .b(new_n198), .out0(new_n199));
  tech160nm_fioaoi03aa1n03p5x5 g104(.a(\a[17] ), .b(\b[16] ), .c(new_n191), .o1(new_n200));
  xnrc02aa1n03x5               g105(.a(new_n200), .b(new_n199), .out0(\s[18] ));
  nano22aa1n03x7               g106(.a(new_n199), .b(new_n194), .c(new_n195), .out0(new_n202));
  tech160nm_fioai012aa1n03p5x5 g107(.a(new_n202), .b(new_n190), .c(new_n186), .o1(new_n203));
  aoai13aa1n12x5               g108(.a(new_n198), .b(new_n197), .c(new_n192), .d(new_n193), .o1(new_n204));
  nor042aa1d18x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand02aa1d04x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  xobna2aa1n03x5               g112(.a(new_n207), .b(new_n203), .c(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n03x5               g114(.a(new_n204), .o1(new_n210));
  oaoi13aa1n03x5               g115(.a(new_n210), .b(new_n202), .c(new_n190), .d(new_n186), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n205), .o1(new_n212));
  nor042aa1n04x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d04x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  oaoi13aa1n02x7               g120(.a(new_n215), .b(new_n212), .c(new_n211), .d(new_n207), .o1(new_n216));
  tech160nm_fiaoi012aa1n02p5x5 g121(.a(new_n207), .b(new_n203), .c(new_n204), .o1(new_n217));
  nano22aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n215), .out0(new_n218));
  norp02aa1n03x5               g123(.a(new_n216), .b(new_n218), .o1(\s[20] ));
  nano23aa1n06x5               g124(.a(new_n205), .b(new_n213), .c(new_n214), .d(new_n206), .out0(new_n220));
  nanp02aa1n06x5               g125(.a(new_n202), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  nona23aa1n09x5               g127(.a(new_n214), .b(new_n206), .c(new_n205), .d(new_n213), .out0(new_n223));
  tech160nm_fiaoi012aa1n05x5   g128(.a(new_n213), .b(new_n205), .c(new_n214), .o1(new_n224));
  oai012aa1n12x5               g129(.a(new_n224), .b(new_n223), .c(new_n204), .o1(new_n225));
  oaoi13aa1n06x5               g130(.a(new_n225), .b(new_n222), .c(new_n190), .d(new_n186), .o1(new_n226));
  xnrb03aa1n03x5               g131(.a(new_n226), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  tech160nm_fixnrc02aa1n04x5   g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  tech160nm_fixnrc02aa1n05x5   g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  oaoi13aa1n02x7               g136(.a(new_n231), .b(new_n229), .c(new_n226), .d(new_n230), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n225), .o1(new_n233));
  oaoi13aa1n09x5               g138(.a(new_n230), .b(new_n233), .c(new_n191), .d(new_n221), .o1(new_n234));
  nano22aa1n03x5               g139(.a(new_n234), .b(new_n229), .c(new_n231), .out0(new_n235));
  norp02aa1n03x5               g140(.a(new_n232), .b(new_n235), .o1(\s[22] ));
  nor042aa1n03x5               g141(.a(new_n231), .b(new_n230), .o1(new_n237));
  norb02aa1n03x5               g142(.a(new_n237), .b(new_n221), .out0(new_n238));
  oao003aa1n06x5               g143(.a(\a[22] ), .b(\b[21] ), .c(new_n229), .carry(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  tech160nm_fiaoi012aa1n02p5x5 g145(.a(new_n240), .b(new_n225), .c(new_n237), .o1(new_n241));
  inv020aa1n03x5               g146(.a(new_n241), .o1(new_n242));
  oaoi13aa1n06x5               g147(.a(new_n242), .b(new_n238), .c(new_n190), .d(new_n186), .o1(new_n243));
  xnrb03aa1n03x5               g148(.a(new_n243), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[22] ), .b(\a[23] ), .out0(new_n247));
  tech160nm_fixnrc02aa1n05x5   g152(.a(\b[23] ), .b(\a[24] ), .out0(new_n248));
  oaoi13aa1n02x7               g153(.a(new_n248), .b(new_n246), .c(new_n243), .d(new_n247), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n238), .o1(new_n250));
  oaoi13aa1n06x5               g155(.a(new_n247), .b(new_n241), .c(new_n191), .d(new_n250), .o1(new_n251));
  nano22aa1n03x5               g156(.a(new_n251), .b(new_n246), .c(new_n248), .out0(new_n252));
  norp02aa1n03x5               g157(.a(new_n249), .b(new_n252), .o1(\s[24] ));
  norp02aa1n02x5               g158(.a(new_n248), .b(new_n247), .o1(new_n254));
  nano22aa1n06x5               g159(.a(new_n221), .b(new_n237), .c(new_n254), .out0(new_n255));
  oai012aa1n06x5               g160(.a(new_n255), .b(new_n190), .c(new_n186), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n224), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n237), .b(new_n257), .c(new_n220), .d(new_n210), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n254), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .c(new_n246), .carry(new_n260));
  aoai13aa1n12x5               g165(.a(new_n260), .b(new_n259), .c(new_n258), .d(new_n239), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[24] ), .b(\a[25] ), .out0(new_n263));
  xobna2aa1n03x5               g168(.a(new_n263), .b(new_n256), .c(new_n262), .out0(\s[25] ));
  oaoi13aa1n03x5               g169(.a(new_n261), .b(new_n255), .c(new_n190), .d(new_n186), .o1(new_n265));
  nor042aa1n03x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnrc02aa1n06x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  oaoi13aa1n02x7               g173(.a(new_n268), .b(new_n267), .c(new_n265), .d(new_n263), .o1(new_n269));
  aoi012aa1n02x7               g174(.a(new_n263), .b(new_n256), .c(new_n262), .o1(new_n270));
  nano22aa1n03x5               g175(.a(new_n270), .b(new_n267), .c(new_n268), .out0(new_n271));
  norp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[26] ));
  nor042aa1n02x5               g177(.a(new_n268), .b(new_n263), .o1(new_n273));
  nano32aa1n03x7               g178(.a(new_n221), .b(new_n273), .c(new_n237), .d(new_n254), .out0(new_n274));
  oai012aa1n06x5               g179(.a(new_n274), .b(new_n190), .c(new_n186), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .c(new_n267), .carry(new_n276));
  aobi12aa1n06x5               g181(.a(new_n276), .b(new_n261), .c(new_n273), .out0(new_n277));
  xorc02aa1n02x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n277), .c(new_n275), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv040aa1n03x5               g185(.a(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n99), .o1(new_n282));
  oaoi13aa1n02x5               g187(.a(new_n282), .b(new_n107), .c(new_n103), .d(new_n106), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n123), .o1(new_n284));
  nano22aa1n03x7               g189(.a(new_n154), .b(new_n167), .c(new_n184), .out0(new_n285));
  aoai13aa1n02x5               g190(.a(new_n285), .b(new_n284), .c(new_n283), .d(new_n116), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n184), .b(new_n169), .c(new_n157), .d(new_n167), .o1(new_n287));
  nanp03aa1n03x5               g192(.a(new_n286), .b(new_n287), .c(new_n189), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n254), .b(new_n240), .c(new_n225), .d(new_n237), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n273), .o1(new_n290));
  aoai13aa1n04x5               g195(.a(new_n276), .b(new_n290), .c(new_n289), .d(new_n260), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n278), .b(new_n291), .c(new_n288), .d(new_n274), .o1(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .out0(new_n293));
  aoi012aa1n02x5               g198(.a(new_n293), .b(new_n292), .c(new_n281), .o1(new_n294));
  aobi12aa1n03x5               g199(.a(new_n278), .b(new_n277), .c(new_n275), .out0(new_n295));
  nano22aa1n03x5               g200(.a(new_n295), .b(new_n281), .c(new_n293), .out0(new_n296));
  norp02aa1n03x5               g201(.a(new_n294), .b(new_n296), .o1(\s[28] ));
  norb02aa1n02x5               g202(.a(new_n278), .b(new_n293), .out0(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n291), .c(new_n288), .d(new_n274), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .c(new_n281), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[28] ), .b(\a[29] ), .out0(new_n301));
  aoi012aa1n02x5               g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  aobi12aa1n03x5               g207(.a(new_n298), .b(new_n277), .c(new_n275), .out0(new_n303));
  nano22aa1n03x5               g208(.a(new_n303), .b(new_n300), .c(new_n301), .out0(new_n304));
  norp02aa1n03x5               g209(.a(new_n302), .b(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g211(.a(new_n278), .b(new_n301), .c(new_n293), .out0(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n291), .c(new_n288), .d(new_n274), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[29] ), .b(\a[30] ), .out0(new_n310));
  aoi012aa1n02x5               g215(.a(new_n310), .b(new_n308), .c(new_n309), .o1(new_n311));
  aobi12aa1n03x5               g216(.a(new_n307), .b(new_n277), .c(new_n275), .out0(new_n312));
  nano22aa1n03x5               g217(.a(new_n312), .b(new_n309), .c(new_n310), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[30] ));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  norb02aa1n02x5               g220(.a(new_n307), .b(new_n310), .out0(new_n316));
  aoai13aa1n02x5               g221(.a(new_n316), .b(new_n291), .c(new_n288), .d(new_n274), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .carry(new_n318));
  aoi012aa1n02x5               g223(.a(new_n315), .b(new_n317), .c(new_n318), .o1(new_n319));
  aobi12aa1n03x5               g224(.a(new_n316), .b(new_n277), .c(new_n275), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n320), .b(new_n315), .c(new_n318), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[31] ));
  nanb02aa1n02x5               g227(.a(new_n104), .b(new_n105), .out0(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n323), .b(new_n132), .c(new_n101), .out0(\s[3] ));
  xorc02aa1n02x5               g229(.a(\a[4] ), .b(\b[3] ), .out0(new_n325));
  aoi112aa1n02x5               g230(.a(new_n325), .b(new_n104), .c(new_n133), .d(new_n132), .o1(new_n326));
  oaoi13aa1n02x5               g231(.a(new_n326), .b(new_n283), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g232(.a(new_n135), .b(\b[4] ), .c(new_n120), .out0(\s[5] ));
  oao003aa1n02x5               g233(.a(\a[5] ), .b(\b[4] ), .c(new_n135), .carry(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g235(.a(\a[6] ), .b(\b[5] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g237(.a(new_n111), .b(new_n331), .c(new_n112), .o1(new_n333));
  xnrb03aa1n02x5               g238(.a(new_n333), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g239(.a(new_n125), .b(new_n117), .c(new_n123), .out0(\s[9] ));
endmodule


