// Benchmark "adder" written by ABC on Thu Jul 18 01:32:26 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n339, new_n340, new_n342, new_n344, new_n346, new_n348, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  tech160nm_fiaoi012aa1n05x5   g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  norp02aa1n04x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n03x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  tech160nm_fiaoi012aa1n03p5x5 g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  oaih12aa1n06x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  nor042aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nand22aa1n03x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  norp02aa1n04x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nona23aa1n02x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  xorc02aa1n12x5               g017(.a(\a[8] ), .b(\b[7] ), .out0(new_n113));
  nor042aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  and002aa1n12x5               g019(.a(\b[6] ), .b(\a[7] ), .o(new_n115));
  norp02aa1n06x5               g020(.a(new_n115), .b(new_n114), .o1(new_n116));
  nano22aa1n03x7               g021(.a(new_n112), .b(new_n113), .c(new_n116), .out0(new_n117));
  aoi012aa1n02x5               g022(.a(new_n108), .b(new_n110), .c(new_n109), .o1(new_n118));
  nanb03aa1n06x5               g023(.a(new_n118), .b(new_n113), .c(new_n116), .out0(new_n119));
  inv000aa1d42x5               g024(.a(new_n114), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  nanb02aa1n06x5               g026(.a(new_n121), .b(new_n119), .out0(new_n122));
  tech160nm_fiaoi012aa1n04x5   g027(.a(new_n122), .b(new_n107), .c(new_n117), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .c(new_n123), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  orn002aa1n02x5               g030(.a(\a[10] ), .b(\b[9] ), .o(new_n126));
  nand42aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  xnrc02aa1n03x5               g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  nano22aa1n02x4               g033(.a(new_n128), .b(new_n126), .c(new_n127), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n122), .c(new_n107), .d(new_n117), .o1(new_n130));
  oai022aa1d18x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(new_n131), .b(new_n127), .o1(new_n132));
  nor042aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n130), .c(new_n132), .out0(\s[11] ));
  nor042aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  nanp02aa1n09x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n130), .b(new_n132), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n133), .b(new_n140), .c(new_n134), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n138), .c(new_n139), .out0(\s[12] ));
  norb02aa1n02x5               g047(.a(new_n102), .b(new_n101), .out0(new_n143));
  norb02aa1n02x5               g048(.a(new_n104), .b(new_n103), .out0(new_n144));
  nanb03aa1n03x5               g049(.a(new_n100), .b(new_n144), .c(new_n143), .out0(new_n145));
  nano23aa1n02x4               g050(.a(new_n108), .b(new_n110), .c(new_n111), .d(new_n109), .out0(new_n146));
  nanp03aa1n02x5               g051(.a(new_n146), .b(new_n113), .c(new_n116), .o1(new_n147));
  tech160nm_fiao0012aa1n02p5x5 g052(.a(new_n108), .b(new_n110), .c(new_n109), .o(new_n148));
  aoi013aa1n06x4               g053(.a(new_n121), .b(new_n148), .c(new_n113), .d(new_n116), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n147), .c(new_n145), .d(new_n106), .o1(new_n150));
  nano23aa1n02x5               g055(.a(new_n133), .b(new_n137), .c(new_n139), .d(new_n134), .out0(new_n151));
  nanp02aa1n02x5               g056(.a(new_n129), .b(new_n151), .o1(new_n152));
  nanb02aa1n02x5               g057(.a(new_n152), .b(new_n150), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n133), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n139), .o1(new_n155));
  nanp03aa1n06x5               g060(.a(new_n131), .b(new_n127), .c(new_n134), .o1(new_n156));
  aoai13aa1n12x5               g061(.a(new_n138), .b(new_n155), .c(new_n156), .d(new_n154), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nor042aa1n06x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n153), .c(new_n158), .out0(\s[13] ));
  nanp02aa1n02x5               g067(.a(new_n107), .b(new_n117), .o1(new_n163));
  aoai13aa1n06x5               g068(.a(new_n158), .b(new_n152), .c(new_n163), .d(new_n149), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n159), .b(new_n164), .c(new_n160), .o1(new_n165));
  xnrb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand42aa1n04x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nano23aa1d15x5               g073(.a(new_n159), .b(new_n167), .c(new_n168), .d(new_n160), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  oa0012aa1n02x5               g075(.a(new_n168), .b(new_n167), .c(new_n159), .o(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n04x5               g077(.a(new_n172), .b(new_n170), .c(new_n153), .d(new_n158), .o1(new_n173));
  nor042aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nanp02aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  norb02aa1n06x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  aoi112aa1n02x5               g081(.a(new_n176), .b(new_n171), .c(new_n164), .d(new_n169), .o1(new_n177));
  aoi012aa1n02x5               g082(.a(new_n177), .b(new_n173), .c(new_n176), .o1(\s[15] ));
  xorc02aa1n12x5               g083(.a(\a[16] ), .b(\b[15] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n174), .c(new_n173), .d(new_n175), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n176), .b(new_n171), .c(new_n164), .d(new_n169), .o1(new_n182));
  nona22aa1n02x5               g087(.a(new_n182), .b(new_n180), .c(new_n174), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n181), .b(new_n183), .o1(\s[16] ));
  nand23aa1d12x5               g089(.a(new_n169), .b(new_n176), .c(new_n179), .o1(new_n185));
  nano22aa1n09x5               g090(.a(new_n185), .b(new_n129), .c(new_n151), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n122), .c(new_n107), .d(new_n117), .o1(new_n187));
  inv040aa1n03x5               g092(.a(new_n185), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\a[16] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[15] ), .o1(new_n190));
  oai112aa1n04x5               g095(.a(new_n168), .b(new_n175), .c(new_n167), .d(new_n159), .o1(new_n191));
  tech160nm_fioai012aa1n03p5x5 g096(.a(new_n191), .b(\b[14] ), .c(\a[15] ), .o1(new_n192));
  oaoi03aa1n09x5               g097(.a(new_n189), .b(new_n190), .c(new_n192), .o1(new_n193));
  inv000aa1n02x5               g098(.a(new_n193), .o1(new_n194));
  aoi012aa1d18x5               g099(.a(new_n194), .b(new_n157), .c(new_n188), .o1(new_n195));
  oaib12aa1n12x5               g100(.a(new_n195), .b(new_n123), .c(new_n186), .out0(new_n196));
  nor002aa1n16x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nand42aa1n03x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  aoi112aa1n02x5               g104(.a(new_n194), .b(new_n199), .c(new_n157), .d(new_n188), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n196), .b(new_n199), .c(new_n187), .d(new_n200), .o1(\s[17] ));
  inv000aa1d42x5               g106(.a(\a[18] ), .o1(new_n202));
  tech160nm_fiaoi012aa1n05x5   g107(.a(new_n197), .b(new_n196), .c(new_n199), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[17] ), .c(new_n202), .out0(\s[18] ));
  nanp02aa1n02x5               g109(.a(new_n156), .b(new_n154), .o1(new_n205));
  nanp02aa1n02x5               g110(.a(new_n205), .b(new_n139), .o1(new_n206));
  aoai13aa1n09x5               g111(.a(new_n193), .b(new_n185), .c(new_n206), .d(new_n138), .o1(new_n207));
  nor042aa1n09x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand22aa1n09x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nano23aa1d15x5               g114(.a(new_n197), .b(new_n208), .c(new_n209), .d(new_n198), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n207), .c(new_n150), .d(new_n186), .o1(new_n211));
  oa0012aa1n02x5               g116(.a(new_n209), .b(new_n208), .c(new_n197), .o(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  nor042aa1n04x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nanp02aa1n04x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norb02aa1n06x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n211), .c(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g123(.a(new_n211), .b(new_n213), .o1(new_n219));
  nor042aa1n04x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nand02aa1n08x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nanb02aa1n02x5               g126(.a(new_n220), .b(new_n221), .out0(new_n222));
  aoai13aa1n02x5               g127(.a(new_n222), .b(new_n214), .c(new_n219), .d(new_n215), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n216), .b(new_n212), .c(new_n196), .d(new_n210), .o1(new_n224));
  nona22aa1n03x5               g129(.a(new_n224), .b(new_n222), .c(new_n214), .out0(new_n225));
  nanp02aa1n03x5               g130(.a(new_n223), .b(new_n225), .o1(\s[20] ));
  nanb03aa1d18x5               g131(.a(new_n222), .b(new_n210), .c(new_n216), .out0(new_n227));
  nanb03aa1n06x5               g132(.a(new_n220), .b(new_n221), .c(new_n215), .out0(new_n228));
  orn002aa1n03x5               g133(.a(\a[19] ), .b(\b[18] ), .o(new_n229));
  oai112aa1n06x5               g134(.a(new_n229), .b(new_n209), .c(new_n208), .d(new_n197), .o1(new_n230));
  aoi012aa1n12x5               g135(.a(new_n220), .b(new_n214), .c(new_n221), .o1(new_n231));
  oai012aa1n18x5               g136(.a(new_n231), .b(new_n230), .c(new_n228), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n04x5               g138(.a(new_n233), .b(new_n227), .c(new_n195), .d(new_n187), .o1(new_n234));
  nor042aa1n04x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  tech160nm_finand02aa1n03p5x5 g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n227), .o1(new_n238));
  aoi112aa1n02x5               g143(.a(new_n237), .b(new_n232), .c(new_n196), .d(new_n238), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n234), .c(new_n237), .o1(\s[21] ));
  nor042aa1n04x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  nand02aa1n08x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n242), .b(new_n241), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n235), .c(new_n234), .d(new_n237), .o1(new_n245));
  nanp02aa1n02x5               g150(.a(new_n234), .b(new_n237), .o1(new_n246));
  nona22aa1n02x5               g151(.a(new_n246), .b(new_n244), .c(new_n235), .out0(new_n247));
  nanp02aa1n03x5               g152(.a(new_n247), .b(new_n245), .o1(\s[22] ));
  nano23aa1n09x5               g153(.a(new_n235), .b(new_n241), .c(new_n242), .d(new_n236), .out0(new_n249));
  nanb02aa1n02x5               g154(.a(new_n227), .b(new_n249), .out0(new_n250));
  aoi012aa1n02x5               g155(.a(new_n250), .b(new_n195), .c(new_n187), .o1(new_n251));
  aoi012aa1d18x5               g156(.a(new_n241), .b(new_n235), .c(new_n242), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  aoi012aa1n02x5               g158(.a(new_n253), .b(new_n232), .c(new_n249), .o1(new_n254));
  aoai13aa1n04x5               g159(.a(new_n254), .b(new_n250), .c(new_n195), .d(new_n187), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  aoi112aa1n02x5               g161(.a(new_n256), .b(new_n253), .c(new_n232), .d(new_n249), .o1(new_n257));
  aboi22aa1n03x5               g162(.a(new_n251), .b(new_n257), .c(new_n255), .d(new_n256), .out0(\s[23] ));
  norp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  tech160nm_fixnrc02aa1n05x5   g164(.a(\b[23] ), .b(\a[24] ), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n259), .c(new_n255), .d(new_n256), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(new_n255), .b(new_n256), .o1(new_n262));
  nona22aa1n02x4               g167(.a(new_n262), .b(new_n260), .c(new_n259), .out0(new_n263));
  nanp02aa1n03x5               g168(.a(new_n263), .b(new_n261), .o1(\s[24] ));
  norb02aa1n12x5               g169(.a(new_n256), .b(new_n260), .out0(new_n265));
  nano22aa1n03x7               g170(.a(new_n227), .b(new_n265), .c(new_n249), .out0(new_n266));
  aoai13aa1n02x5               g171(.a(new_n266), .b(new_n207), .c(new_n150), .d(new_n186), .o1(new_n267));
  nano22aa1n03x5               g172(.a(new_n220), .b(new_n215), .c(new_n221), .out0(new_n268));
  oai012aa1n02x5               g173(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .o1(new_n269));
  oab012aa1n02x5               g174(.a(new_n269), .b(new_n197), .c(new_n208), .out0(new_n270));
  inv020aa1n02x5               g175(.a(new_n231), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n249), .b(new_n271), .c(new_n270), .d(new_n268), .o1(new_n272));
  inv000aa1n02x5               g177(.a(new_n265), .o1(new_n273));
  orn002aa1n02x5               g178(.a(\a[23] ), .b(\b[22] ), .o(new_n274));
  oao003aa1n02x5               g179(.a(\a[24] ), .b(\b[23] ), .c(new_n274), .carry(new_n275));
  aoai13aa1n12x5               g180(.a(new_n275), .b(new_n273), .c(new_n272), .d(new_n252), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  nand42aa1n03x5               g182(.a(new_n267), .b(new_n277), .o1(new_n278));
  tech160nm_fixorc02aa1n05x5   g183(.a(\a[25] ), .b(\b[24] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n265), .b(new_n253), .c(new_n232), .d(new_n249), .o1(new_n280));
  nano22aa1n02x4               g185(.a(new_n279), .b(new_n280), .c(new_n275), .out0(new_n281));
  aoi022aa1n02x5               g186(.a(new_n278), .b(new_n279), .c(new_n267), .d(new_n281), .o1(\s[25] ));
  norp02aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  xorc02aa1n12x5               g188(.a(\a[26] ), .b(\b[25] ), .out0(new_n284));
  inv000aa1d42x5               g189(.a(new_n284), .o1(new_n285));
  aoai13aa1n02x5               g190(.a(new_n285), .b(new_n283), .c(new_n278), .d(new_n279), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n279), .b(new_n276), .c(new_n196), .d(new_n266), .o1(new_n287));
  nona22aa1n03x5               g192(.a(new_n287), .b(new_n285), .c(new_n283), .out0(new_n288));
  nanp02aa1n03x5               g193(.a(new_n286), .b(new_n288), .o1(\s[26] ));
  and002aa1n24x5               g194(.a(new_n284), .b(new_n279), .o(new_n290));
  nano32aa1d15x5               g195(.a(new_n227), .b(new_n290), .c(new_n249), .d(new_n265), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n207), .c(new_n150), .d(new_n186), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\a[26] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[25] ), .o1(new_n294));
  oaoi03aa1n09x5               g199(.a(new_n293), .b(new_n294), .c(new_n283), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoi012aa1n09x5               g201(.a(new_n296), .b(new_n276), .c(new_n290), .o1(new_n297));
  nanp02aa1n06x5               g202(.a(new_n297), .b(new_n292), .o1(new_n298));
  xorc02aa1n12x5               g203(.a(\a[27] ), .b(\b[26] ), .out0(new_n299));
  aoi112aa1n02x5               g204(.a(new_n299), .b(new_n296), .c(new_n276), .d(new_n290), .o1(new_n300));
  aoi022aa1n02x5               g205(.a(new_n298), .b(new_n299), .c(new_n292), .d(new_n300), .o1(\s[27] ));
  norp02aa1n02x5               g206(.a(\b[26] ), .b(\a[27] ), .o1(new_n302));
  norp02aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .o1(new_n303));
  nanp02aa1n02x5               g208(.a(\b[27] ), .b(\a[28] ), .o1(new_n304));
  nanb02aa1n06x5               g209(.a(new_n303), .b(new_n304), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n302), .c(new_n298), .d(new_n299), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n290), .o1(new_n307));
  aoai13aa1n06x5               g212(.a(new_n295), .b(new_n307), .c(new_n280), .d(new_n275), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n299), .b(new_n308), .c(new_n196), .d(new_n291), .o1(new_n309));
  nona22aa1n02x5               g214(.a(new_n309), .b(new_n305), .c(new_n302), .out0(new_n310));
  nanp02aa1n03x5               g215(.a(new_n306), .b(new_n310), .o1(\s[28] ));
  norb02aa1n03x5               g216(.a(new_n299), .b(new_n305), .out0(new_n312));
  aoai13aa1n06x5               g217(.a(new_n312), .b(new_n308), .c(new_n196), .d(new_n291), .o1(new_n313));
  tech160nm_fixorc02aa1n05x5   g218(.a(\a[29] ), .b(\b[28] ), .out0(new_n314));
  oai012aa1n02x5               g219(.a(new_n304), .b(new_n303), .c(new_n302), .o1(new_n315));
  norb02aa1n02x5               g220(.a(new_n315), .b(new_n314), .out0(new_n316));
  inv000aa1d42x5               g221(.a(new_n312), .o1(new_n317));
  aoai13aa1n02x5               g222(.a(new_n315), .b(new_n317), .c(new_n297), .d(new_n292), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n313), .d(new_n316), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g225(.a(new_n305), .b(new_n299), .c(new_n314), .out0(new_n321));
  aoai13aa1n06x5               g226(.a(new_n321), .b(new_n308), .c(new_n196), .d(new_n291), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[29] ), .b(\b[28] ), .c(new_n315), .carry(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(new_n325));
  inv000aa1n02x5               g230(.a(new_n321), .o1(new_n326));
  aoai13aa1n03x5               g231(.a(new_n324), .b(new_n326), .c(new_n297), .d(new_n292), .o1(new_n327));
  aoi022aa1n02x7               g232(.a(new_n327), .b(new_n323), .c(new_n322), .d(new_n325), .o1(\s[30] ));
  nand03aa1n02x5               g233(.a(new_n312), .b(new_n314), .c(new_n323), .o1(new_n329));
  nanb02aa1n02x5               g234(.a(new_n329), .b(new_n298), .out0(new_n330));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  and002aa1n02x5               g236(.a(\b[29] ), .b(\a[30] ), .o(new_n332));
  oabi12aa1n02x5               g237(.a(new_n331), .b(\a[30] ), .c(\b[29] ), .out0(new_n333));
  oab012aa1n02x4               g238(.a(new_n333), .b(new_n324), .c(new_n332), .out0(new_n334));
  oao003aa1n02x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n324), .carry(new_n335));
  aoai13aa1n02x7               g240(.a(new_n335), .b(new_n329), .c(new_n297), .d(new_n292), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n330), .b(new_n334), .c(new_n336), .d(new_n331), .o1(\s[31] ));
  xnrb03aa1n02x5               g242(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoai13aa1n02x5               g243(.a(new_n144), .b(new_n97), .c(new_n99), .d(new_n98), .o1(new_n339));
  aoib12aa1n02x5               g244(.a(new_n103), .b(new_n102), .c(new_n101), .out0(new_n340));
  aboi22aa1n03x5               g245(.a(new_n101), .b(new_n107), .c(new_n339), .d(new_n340), .out0(\s[4] ));
  norb02aa1n02x5               g246(.a(new_n111), .b(new_n110), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n342), .b(new_n145), .c(new_n106), .out0(\s[5] ));
  tech160nm_fiao0012aa1n02p5x5 g248(.a(new_n110), .b(new_n107), .c(new_n111), .o(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi012aa1n03x5               g250(.a(new_n108), .b(new_n344), .c(new_n109), .o1(new_n346));
  xnrc02aa1n02x5               g251(.a(new_n346), .b(new_n116), .out0(\s[7] ));
  aoi112aa1n03x4               g252(.a(new_n115), .b(new_n113), .c(new_n346), .d(new_n120), .o1(new_n348));
  aoai13aa1n02x5               g253(.a(new_n113), .b(new_n115), .c(new_n346), .d(new_n120), .o1(new_n349));
  nanb02aa1n03x5               g254(.a(new_n348), .b(new_n349), .out0(\s[8] ));
  xobna2aa1n03x5               g255(.a(new_n128), .b(new_n163), .c(new_n149), .out0(\s[9] ));
endmodule


