// Benchmark "adder" written by ABC on Wed Jul 17 19:23:18 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n179, new_n180, new_n181,
    new_n182, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n328, new_n331, new_n332, new_n333,
    new_n334, new_n336, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  xnrc02aa1n12x5               g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  orn002aa1n24x5               g004(.a(\a[2] ), .b(\b[1] ), .o(new_n100));
  nand42aa1n04x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n12x5               g006(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(new_n102));
  norp02aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1d28x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb03aa1n03x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n106));
  aoai13aa1n12x5               g011(.a(new_n106), .b(new_n99), .c(new_n102), .d(new_n100), .o1(new_n107));
  nand42aa1n16x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  aoi022aa1d24x5               g013(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n109));
  oai112aa1n06x5               g014(.a(new_n109), .b(new_n108), .c(\b[7] ), .d(\a[8] ), .o1(new_n110));
  tech160nm_fixnrc02aa1n04x5   g015(.a(\b[4] ), .b(\a[5] ), .out0(new_n111));
  oai122aa1n06x5               g016(.a(new_n104), .b(\a[7] ), .c(\b[6] ), .d(\a[6] ), .e(\b[5] ), .o1(new_n112));
  nor043aa1d12x5               g017(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n113));
  nand02aa1n03x5               g018(.a(new_n109), .b(new_n108), .o1(new_n114));
  oai022aa1d18x5               g019(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n115));
  inv000aa1n06x5               g020(.a(new_n115), .o1(new_n116));
  tech160nm_fiaoi012aa1n04x5   g021(.a(new_n116), .b(\a[8] ), .c(\b[7] ), .o1(new_n117));
  inv020aa1n04x5               g022(.a(new_n117), .o1(new_n118));
  norp02aa1n04x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nor042aa1n02x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  norb03aa1n09x5               g025(.a(new_n108), .b(new_n120), .c(new_n119), .out0(new_n121));
  oai013aa1n06x5               g026(.a(new_n118), .b(new_n121), .c(new_n114), .d(new_n115), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  norb02aa1n02x5               g028(.a(new_n123), .b(new_n97), .out0(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n122), .c(new_n107), .d(new_n113), .o1(new_n125));
  xnrc02aa1n12x5               g030(.a(\b[9] ), .b(\a[10] ), .out0(new_n126));
  xobna2aa1n03x5               g031(.a(new_n126), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  nor042aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  and002aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o(new_n129));
  oabi12aa1n02x5               g034(.a(new_n129), .b(new_n97), .c(new_n128), .out0(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n126), .c(new_n125), .d(new_n98), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand22aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norp02aa1n12x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nand22aa1n09x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  aoai13aa1n02x5               g042(.a(new_n137), .b(new_n133), .c(new_n131), .d(new_n134), .o1(new_n138));
  aoi112aa1n02x5               g043(.a(new_n133), .b(new_n137), .c(new_n131), .d(new_n134), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n138), .b(new_n139), .out0(\s[12] ));
  nona23aa1n03x5               g045(.a(new_n136), .b(new_n134), .c(new_n133), .d(new_n135), .out0(new_n141));
  nano23aa1n03x7               g046(.a(new_n141), .b(new_n126), .c(new_n123), .d(new_n98), .out0(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n122), .c(new_n107), .d(new_n113), .o1(new_n143));
  oab012aa1n03x5               g048(.a(new_n129), .b(new_n97), .c(new_n128), .out0(new_n144));
  nano23aa1n06x5               g049(.a(new_n133), .b(new_n135), .c(new_n136), .d(new_n134), .out0(new_n145));
  tech160nm_fiao0012aa1n05x5   g050(.a(new_n135), .b(new_n133), .c(new_n136), .o(new_n146));
  aoi012aa1n06x5               g051(.a(new_n146), .b(new_n145), .c(new_n144), .o1(new_n147));
  xnrc02aa1n12x5               g052(.a(\b[12] ), .b(\a[13] ), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  xnbna2aa1n03x5               g054(.a(new_n149), .b(new_n143), .c(new_n147), .out0(\s[13] ));
  orn002aa1n02x5               g055(.a(\a[13] ), .b(\b[12] ), .o(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n148), .c(new_n143), .d(new_n147), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xnrc02aa1n12x5               g058(.a(\b[13] ), .b(\a[14] ), .out0(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n155), .b(new_n149), .o1(new_n156));
  oaih22aa1d12x5               g061(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n157));
  aob012aa1n12x5               g062(.a(new_n157), .b(\b[13] ), .c(\a[14] ), .out0(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n156), .c(new_n143), .d(new_n147), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor022aa1n08x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nor002aa1n12x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nanp02aa1n04x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  aoai13aa1n03x5               g070(.a(new_n165), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n161), .b(new_n165), .c(new_n159), .d(new_n162), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(\s[16] ));
  tech160nm_fiaoi012aa1n05x5   g073(.a(new_n122), .b(new_n107), .c(new_n113), .o1(new_n169));
  nona23aa1n03x5               g074(.a(new_n164), .b(new_n162), .c(new_n161), .d(new_n163), .out0(new_n170));
  nor043aa1n03x5               g075(.a(new_n170), .b(new_n154), .c(new_n148), .o1(new_n171));
  nand42aa1n02x5               g076(.a(new_n142), .b(new_n171), .o1(new_n172));
  oabi12aa1n03x5               g077(.a(new_n146), .b(new_n141), .c(new_n130), .out0(new_n173));
  aoi112aa1n09x5               g078(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n174));
  oai022aa1n02x7               g079(.a(new_n170), .b(new_n158), .c(\b[15] ), .d(\a[16] ), .o1(new_n175));
  aoi112aa1n06x5               g080(.a(new_n175), .b(new_n174), .c(new_n173), .d(new_n171), .o1(new_n176));
  oai012aa1n12x5               g081(.a(new_n176), .b(new_n169), .c(new_n172), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g083(.a(\a[18] ), .o1(new_n179));
  inv000aa1d42x5               g084(.a(\a[17] ), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\b[16] ), .o1(new_n181));
  oaoi03aa1n02x5               g086(.a(new_n180), .b(new_n181), .c(new_n177), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[17] ), .c(new_n179), .out0(\s[18] ));
  nanp02aa1n06x5               g088(.a(new_n107), .b(new_n113), .o1(new_n184));
  nor003aa1n03x5               g089(.a(new_n121), .b(new_n114), .c(new_n115), .o1(new_n185));
  nor022aa1n04x5               g090(.a(new_n185), .b(new_n117), .o1(new_n186));
  nand02aa1d06x5               g091(.a(new_n184), .b(new_n186), .o1(new_n187));
  nano22aa1n02x4               g092(.a(new_n126), .b(new_n98), .c(new_n123), .out0(new_n188));
  nano23aa1n09x5               g093(.a(new_n161), .b(new_n163), .c(new_n164), .d(new_n162), .out0(new_n189));
  nona22aa1n09x5               g094(.a(new_n189), .b(new_n154), .c(new_n148), .out0(new_n190));
  nano22aa1n06x5               g095(.a(new_n190), .b(new_n188), .c(new_n145), .out0(new_n191));
  inv000aa1d42x5               g096(.a(new_n158), .o1(new_n192));
  aoi112aa1n06x5               g097(.a(new_n163), .b(new_n174), .c(new_n192), .d(new_n189), .o1(new_n193));
  oai012aa1n09x5               g098(.a(new_n193), .b(new_n147), .c(new_n190), .o1(new_n194));
  xroi22aa1d06x4               g099(.a(new_n180), .b(\b[16] ), .c(new_n179), .d(\b[17] ), .out0(new_n195));
  aoai13aa1n03x5               g100(.a(new_n195), .b(new_n194), .c(new_n187), .d(new_n191), .o1(new_n196));
  oai022aa1d24x5               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oaib12aa1n18x5               g102(.a(new_n197), .b(new_n179), .c(\b[17] ), .out0(new_n198));
  nor002aa1n20x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nand02aa1n06x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nanb02aa1d24x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n196), .c(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g109(.a(new_n199), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n198), .o1(new_n206));
  aoai13aa1n02x7               g111(.a(new_n202), .b(new_n206), .c(new_n177), .d(new_n195), .o1(new_n207));
  inv040aa1d32x5               g112(.a(\a[20] ), .o1(new_n208));
  inv040aa1d28x5               g113(.a(\b[19] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(new_n209), .b(new_n208), .o1(new_n210));
  nanp02aa1n06x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nand42aa1n10x5               g116(.a(new_n210), .b(new_n211), .o1(new_n212));
  tech160nm_fiaoi012aa1n02p5x5 g117(.a(new_n212), .b(new_n207), .c(new_n205), .o1(new_n213));
  aoi012aa1n03x5               g118(.a(new_n201), .b(new_n196), .c(new_n198), .o1(new_n214));
  nano22aa1n03x5               g119(.a(new_n214), .b(new_n205), .c(new_n212), .out0(new_n215));
  norp02aa1n03x5               g120(.a(new_n213), .b(new_n215), .o1(\s[20] ));
  nano22aa1n03x7               g121(.a(new_n212), .b(new_n205), .c(new_n200), .out0(new_n217));
  nand22aa1n06x5               g122(.a(new_n195), .b(new_n217), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n06x5               g124(.a(new_n219), .b(new_n194), .c(new_n187), .d(new_n191), .o1(new_n220));
  aoi112aa1n03x5               g125(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n221));
  inv000aa1n02x5               g126(.a(new_n221), .o1(new_n222));
  nor043aa1d12x5               g127(.a(new_n198), .b(new_n201), .c(new_n212), .o1(new_n223));
  nano22aa1d15x5               g128(.a(new_n223), .b(new_n210), .c(new_n222), .out0(new_n224));
  xorc02aa1n12x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n220), .c(new_n224), .out0(\s[21] ));
  norp02aa1n02x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n224), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n225), .b(new_n229), .c(new_n177), .d(new_n219), .o1(new_n230));
  xorc02aa1n12x5               g135(.a(\a[22] ), .b(\b[21] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoi012aa1n03x5               g137(.a(new_n232), .b(new_n230), .c(new_n228), .o1(new_n233));
  aobi12aa1n03x5               g138(.a(new_n225), .b(new_n220), .c(new_n224), .out0(new_n234));
  nano22aa1n03x5               g139(.a(new_n234), .b(new_n228), .c(new_n232), .out0(new_n235));
  norp02aa1n03x5               g140(.a(new_n233), .b(new_n235), .o1(\s[22] ));
  nand02aa1d04x5               g141(.a(new_n231), .b(new_n225), .o1(new_n237));
  nano22aa1n02x4               g142(.a(new_n237), .b(new_n195), .c(new_n217), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n194), .c(new_n187), .d(new_n191), .o1(new_n239));
  inv040aa1d32x5               g144(.a(\a[22] ), .o1(new_n240));
  oai022aa1d18x5               g145(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n241));
  oaib12aa1n06x5               g146(.a(new_n241), .b(new_n240), .c(\b[21] ), .out0(new_n242));
  oa0012aa1n06x5               g147(.a(new_n242), .b(new_n224), .c(new_n237), .o(new_n243));
  tech160nm_fixorc02aa1n03p5x5 g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  xnbna2aa1n03x5               g149(.a(new_n244), .b(new_n239), .c(new_n243), .out0(\s[23] ));
  nor042aa1n04x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  inv040aa1n06x5               g152(.a(new_n243), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n244), .b(new_n248), .c(new_n177), .d(new_n238), .o1(new_n249));
  nor002aa1d32x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  nand02aa1n10x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nanb02aa1d24x5               g156(.a(new_n250), .b(new_n251), .out0(new_n252));
  aoi012aa1n03x5               g157(.a(new_n252), .b(new_n249), .c(new_n247), .o1(new_n253));
  xnrc02aa1n12x5               g158(.a(\b[22] ), .b(\a[23] ), .out0(new_n254));
  tech160nm_fiaoi012aa1n05x5   g159(.a(new_n254), .b(new_n239), .c(new_n243), .o1(new_n255));
  nano22aa1n03x7               g160(.a(new_n255), .b(new_n247), .c(new_n252), .out0(new_n256));
  nor002aa1n02x5               g161(.a(new_n253), .b(new_n256), .o1(\s[24] ));
  inv000aa1d42x5               g162(.a(\a[21] ), .o1(new_n258));
  xroi22aa1d06x4               g163(.a(new_n258), .b(\b[20] ), .c(new_n240), .d(\b[21] ), .out0(new_n259));
  nor002aa1n03x5               g164(.a(new_n254), .b(new_n252), .o1(new_n260));
  nano22aa1n03x7               g165(.a(new_n218), .b(new_n259), .c(new_n260), .out0(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n194), .c(new_n187), .d(new_n191), .o1(new_n262));
  nanp02aa1n03x5               g167(.a(new_n259), .b(new_n260), .o1(new_n263));
  norp03aa1n03x5               g168(.a(new_n254), .b(new_n242), .c(new_n252), .o1(new_n264));
  aoi112aa1n06x5               g169(.a(new_n264), .b(new_n250), .c(new_n251), .d(new_n246), .o1(new_n265));
  oai012aa1d24x5               g170(.a(new_n265), .b(new_n224), .c(new_n263), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnrc02aa1n12x5               g172(.a(\b[24] ), .b(\a[25] ), .out0(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  xnbna2aa1n03x5               g174(.a(new_n269), .b(new_n262), .c(new_n267), .out0(\s[25] ));
  nor042aa1n03x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n269), .b(new_n266), .c(new_n177), .d(new_n261), .o1(new_n273));
  tech160nm_fixnrc02aa1n05x5   g178(.a(\b[25] ), .b(\a[26] ), .out0(new_n274));
  aoi012aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n272), .o1(new_n275));
  aoi012aa1n03x5               g180(.a(new_n268), .b(new_n262), .c(new_n267), .o1(new_n276));
  nano22aa1n03x5               g181(.a(new_n276), .b(new_n272), .c(new_n274), .out0(new_n277));
  norp02aa1n03x5               g182(.a(new_n275), .b(new_n277), .o1(\s[26] ));
  nor042aa1d18x5               g183(.a(new_n274), .b(new_n268), .o1(new_n279));
  nano32aa1n03x7               g184(.a(new_n218), .b(new_n279), .c(new_n259), .d(new_n260), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n194), .c(new_n187), .d(new_n191), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[26] ), .b(\b[25] ), .c(new_n272), .carry(new_n282));
  aobi12aa1n18x5               g187(.a(new_n282), .b(new_n266), .c(new_n279), .out0(new_n283));
  xorc02aa1n12x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  xnbna2aa1n03x5               g189(.a(new_n284), .b(new_n283), .c(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  inv040aa1n03x5               g191(.a(new_n286), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n210), .o1(new_n288));
  norb02aa1n02x5               g193(.a(new_n251), .b(new_n250), .out0(new_n289));
  nano22aa1n02x4               g194(.a(new_n237), .b(new_n244), .c(new_n289), .out0(new_n290));
  oai013aa1n03x5               g195(.a(new_n290), .b(new_n223), .c(new_n288), .d(new_n221), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n279), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n282), .b(new_n292), .c(new_n291), .d(new_n265), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n284), .b(new_n293), .c(new_n177), .d(new_n280), .o1(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  aoi012aa1n02x5               g200(.a(new_n295), .b(new_n294), .c(new_n287), .o1(new_n296));
  aobi12aa1n03x5               g201(.a(new_n284), .b(new_n283), .c(new_n281), .out0(new_n297));
  nano22aa1n03x5               g202(.a(new_n297), .b(new_n287), .c(new_n295), .out0(new_n298));
  norp02aa1n03x5               g203(.a(new_n296), .b(new_n298), .o1(\s[28] ));
  norb02aa1n02x5               g204(.a(new_n284), .b(new_n295), .out0(new_n300));
  aoai13aa1n02x7               g205(.a(new_n300), .b(new_n293), .c(new_n177), .d(new_n280), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[28] ), .b(\a[29] ), .out0(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n301), .c(new_n302), .o1(new_n304));
  aobi12aa1n06x5               g209(.a(new_n300), .b(new_n283), .c(new_n281), .out0(new_n305));
  nano22aa1n03x7               g210(.a(new_n305), .b(new_n302), .c(new_n303), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n304), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g213(.a(new_n284), .b(new_n303), .c(new_n295), .out0(new_n309));
  aoai13aa1n02x5               g214(.a(new_n309), .b(new_n293), .c(new_n177), .d(new_n280), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n302), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .out0(new_n312));
  aoi012aa1n02x5               g217(.a(new_n312), .b(new_n310), .c(new_n311), .o1(new_n313));
  aobi12aa1n03x5               g218(.a(new_n309), .b(new_n283), .c(new_n281), .out0(new_n314));
  nano22aa1n03x5               g219(.a(new_n314), .b(new_n311), .c(new_n312), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n313), .b(new_n315), .o1(\s[30] ));
  norb02aa1n03x4               g221(.a(new_n309), .b(new_n312), .out0(new_n317));
  aobi12aa1n03x5               g222(.a(new_n317), .b(new_n283), .c(new_n281), .out0(new_n318));
  oao003aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n319));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n320), .out0(new_n321));
  aoai13aa1n02x5               g226(.a(new_n317), .b(new_n293), .c(new_n177), .d(new_n280), .o1(new_n322));
  aoi012aa1n02x5               g227(.a(new_n320), .b(new_n322), .c(new_n319), .o1(new_n323));
  norp02aa1n03x5               g228(.a(new_n323), .b(new_n321), .o1(\s[31] ));
  xobna2aa1n03x5               g229(.a(new_n99), .b(new_n102), .c(new_n100), .out0(\s[3] ));
  norb02aa1n02x5               g230(.a(new_n104), .b(new_n105), .out0(new_n326));
  nanp02aa1n02x5               g231(.a(new_n102), .b(new_n100), .o1(new_n327));
  aoib12aa1n02x5               g232(.a(new_n103), .b(new_n327), .c(new_n99), .out0(new_n328));
  oai012aa1n02x5               g233(.a(new_n107), .b(new_n328), .c(new_n326), .o1(\s[4] ));
  xnbna2aa1n03x5               g234(.a(new_n111), .b(new_n107), .c(new_n104), .out0(\s[5] ));
  orn002aa1n02x5               g235(.a(\a[6] ), .b(\b[5] ), .o(new_n331));
  nanb03aa1n02x5               g236(.a(new_n111), .b(new_n107), .c(new_n104), .out0(new_n332));
  norb02aa1n02x5               g237(.a(new_n332), .b(new_n119), .out0(new_n333));
  nanp02aa1n02x5               g238(.a(new_n332), .b(new_n121), .o1(new_n334));
  aoai13aa1n02x5               g239(.a(new_n334), .b(new_n333), .c(new_n108), .d(new_n331), .o1(\s[6] ));
  nanp02aa1n02x5               g240(.a(new_n334), .b(new_n108), .o1(new_n336));
  xnrb03aa1n02x5               g241(.a(new_n336), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g242(.a(\a[7] ), .b(\b[6] ), .c(new_n336), .o1(new_n338));
  xorb03aa1n02x5               g243(.a(new_n338), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g244(.a(new_n124), .b(new_n184), .c(new_n186), .out0(\s[9] ));
endmodule


