// Benchmark "adder" written by ABC on Thu Jul 18 05:26:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n336, new_n338,
    new_n340, new_n342, new_n343, new_n345, new_n346, new_n347, new_n348,
    new_n350, new_n352, new_n353, new_n354;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nand42aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  orn002aa1n02x7               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n03x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  nor042aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n03x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor042aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  tech160nm_finand02aa1n05x5   g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n06x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nand23aa1n04x5               g013(.a(new_n102), .b(new_n105), .c(new_n108), .o1(new_n109));
  tech160nm_fioai012aa1n04x5   g014(.a(new_n104), .b(new_n106), .c(new_n103), .o1(new_n110));
  norp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor042aa1n06x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nand42aa1n06x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nano23aa1n03x7               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  nor042aa1n04x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  tech160nm_finand02aa1n05x5   g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor022aa1n06x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  tech160nm_finand02aa1n05x5   g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano23aa1n09x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nand42aa1n02x5               g025(.a(new_n120), .b(new_n115), .o1(new_n121));
  inv040aa1n02x5               g026(.a(new_n113), .o1(new_n122));
  oaoi03aa1n09x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  oa0012aa1n02x5               g028(.a(new_n117), .b(new_n118), .c(new_n116), .o(new_n124));
  tech160nm_fiaoi012aa1n05x5   g029(.a(new_n124), .b(new_n120), .c(new_n123), .o1(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n126));
  xorc02aa1n02x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n97), .c(new_n126), .d(new_n98), .o1(new_n128));
  aoi112aa1n02x5               g033(.a(new_n127), .b(new_n97), .c(new_n126), .d(new_n98), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n128), .b(new_n129), .out0(\s[10] ));
  nor002aa1n02x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  oai012aa1n02x5               g037(.a(new_n132), .b(new_n131), .c(new_n97), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  tech160nm_finand02aa1n05x5   g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n06x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n128), .c(new_n133), .out0(\s[11] ));
  nor042aa1n03x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n128), .b(new_n133), .o1(new_n139));
  nand02aa1d06x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n138), .b(new_n140), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n134), .c(new_n139), .d(new_n135), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n136), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n140), .b(new_n143), .c(new_n128), .d(new_n133), .o1(new_n144));
  oai013aa1n02x4               g049(.a(new_n142), .b(new_n144), .c(new_n134), .d(new_n138), .o1(\s[12] ));
  norb02aa1n06x5               g050(.a(new_n98), .b(new_n97), .out0(new_n146));
  nano32aa1n03x7               g051(.a(new_n141), .b(new_n127), .c(new_n146), .d(new_n136), .out0(new_n147));
  nano22aa1n03x7               g052(.a(new_n138), .b(new_n135), .c(new_n140), .out0(new_n148));
  tech160nm_fiaoi012aa1n04x5   g053(.a(new_n134), .b(\a[10] ), .c(\b[9] ), .o1(new_n149));
  oai112aa1n06x5               g054(.a(new_n148), .b(new_n149), .c(new_n131), .d(new_n97), .o1(new_n150));
  aoi012aa1n06x5               g055(.a(new_n138), .b(new_n134), .c(new_n140), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n150), .b(new_n151), .o1(new_n152));
  aoi012aa1n02x5               g057(.a(new_n152), .b(new_n126), .c(new_n147), .o1(new_n153));
  nor042aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand02aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n154), .b(new_n155), .out0(new_n156));
  and003aa1n02x5               g061(.a(new_n150), .b(new_n156), .c(new_n151), .o(new_n157));
  aobi12aa1n02x5               g062(.a(new_n157), .b(new_n126), .c(new_n147), .out0(new_n158));
  oab012aa1n02x4               g063(.a(new_n158), .b(new_n153), .c(new_n156), .out0(\s[13] ));
  nor002aa1n20x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  nand22aa1n09x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norp02aa1n02x5               g067(.a(new_n153), .b(new_n156), .o1(new_n163));
  aoi112aa1n02x5               g068(.a(new_n163), .b(new_n154), .c(new_n161), .d(new_n162), .o1(new_n164));
  oaoi03aa1n02x5               g069(.a(\a[13] ), .b(\b[12] ), .c(new_n153), .o1(new_n165));
  aoi013aa1n02x4               g070(.a(new_n164), .b(new_n165), .c(new_n161), .d(new_n162), .o1(\s[14] ));
  nano23aa1n06x5               g071(.a(new_n154), .b(new_n160), .c(new_n162), .d(new_n155), .out0(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n152), .c(new_n126), .d(new_n147), .o1(new_n168));
  aoi012aa1n06x5               g073(.a(new_n160), .b(new_n154), .c(new_n162), .o1(new_n169));
  nor042aa1n06x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand02aa1n03x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n169), .out0(\s[15] ));
  nor042aa1n04x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand42aa1n02x5               g079(.a(new_n168), .b(new_n169), .o1(new_n175));
  nand02aa1d08x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n174), .b(new_n176), .out0(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n170), .c(new_n175), .d(new_n172), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n172), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n176), .b(new_n179), .c(new_n168), .d(new_n169), .o1(new_n180));
  oai013aa1n02x4               g085(.a(new_n178), .b(new_n180), .c(new_n170), .d(new_n174), .o1(\s[16] ));
  aoi012aa1n12x5               g086(.a(new_n174), .b(new_n170), .c(new_n176), .o1(new_n182));
  xnrc02aa1n03x5               g087(.a(\b[16] ), .b(\a[17] ), .out0(new_n183));
  nano23aa1n02x4               g088(.a(new_n97), .b(new_n138), .c(new_n140), .d(new_n98), .out0(new_n184));
  nano23aa1n09x5               g089(.a(new_n170), .b(new_n174), .c(new_n176), .d(new_n171), .out0(new_n185));
  nanp02aa1n03x5               g090(.a(new_n185), .b(new_n167), .o1(new_n186));
  nano32aa1n03x7               g091(.a(new_n186), .b(new_n184), .c(new_n136), .d(new_n127), .out0(new_n187));
  nanp02aa1n02x5               g092(.a(new_n126), .b(new_n187), .o1(new_n188));
  inv020aa1n03x5               g093(.a(new_n169), .o1(new_n189));
  aobi12aa1n06x5               g094(.a(new_n182), .b(new_n185), .c(new_n189), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n186), .c(new_n150), .d(new_n151), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  tech160nm_fiaoi012aa1n05x5   g097(.a(new_n183), .b(new_n188), .c(new_n192), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(new_n175), .b(new_n185), .o1(new_n194));
  aoi013aa1n02x4               g099(.a(new_n193), .b(new_n194), .c(new_n182), .d(new_n183), .o1(\s[17] ));
  nor002aa1n03x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nor042aa1n06x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  inv030aa1n02x5               g102(.a(new_n197), .o1(new_n198));
  nand22aa1n03x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  aoi112aa1n02x5               g104(.a(new_n193), .b(new_n196), .c(new_n198), .d(new_n199), .o1(new_n200));
  oai112aa1n02x5               g105(.a(new_n198), .b(new_n199), .c(new_n193), .d(new_n196), .o1(new_n201));
  norb02aa1n03x4               g106(.a(new_n201), .b(new_n200), .out0(\s[18] ));
  nano22aa1n02x5               g107(.a(new_n183), .b(new_n198), .c(new_n199), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n191), .c(new_n126), .d(new_n187), .o1(new_n204));
  tech160nm_fiaoi012aa1n05x5   g109(.a(new_n197), .b(new_n196), .c(new_n199), .o1(new_n205));
  nor042aa1d18x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nanp02aa1n09x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  norb02aa1n12x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n204), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n208), .o1(new_n212));
  aoi012aa1n03x5               g117(.a(new_n212), .b(new_n204), .c(new_n205), .o1(new_n213));
  nand42aa1n08x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1n06x4               g119(.a(new_n214), .b(new_n211), .out0(new_n215));
  oabi12aa1n03x5               g120(.a(new_n215), .b(new_n213), .c(new_n206), .out0(new_n216));
  aoai13aa1n02x5               g121(.a(new_n214), .b(new_n212), .c(new_n204), .d(new_n205), .o1(new_n217));
  oai013aa1n02x4               g122(.a(new_n216), .b(new_n217), .c(new_n206), .d(new_n211), .o1(\s[20] ));
  nano23aa1d15x5               g123(.a(new_n206), .b(new_n211), .c(new_n214), .d(new_n207), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  norb02aa1n02x5               g125(.a(new_n203), .b(new_n220), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n191), .c(new_n126), .d(new_n187), .o1(new_n222));
  aoi112aa1n09x5               g127(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n223));
  oai112aa1n06x5               g128(.a(new_n208), .b(new_n215), .c(new_n223), .d(new_n197), .o1(new_n224));
  aoi012aa1n12x5               g129(.a(new_n211), .b(new_n206), .c(new_n214), .o1(new_n225));
  nanp02aa1n02x5               g130(.a(new_n224), .b(new_n225), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nanp02aa1n03x5               g132(.a(new_n222), .b(new_n227), .o1(new_n228));
  tech160nm_fixorc02aa1n02p5x5 g133(.a(\a[21] ), .b(\b[20] ), .out0(new_n229));
  inv040aa1n03x5               g134(.a(new_n205), .o1(new_n230));
  inv000aa1n02x5               g135(.a(new_n225), .o1(new_n231));
  aoi112aa1n02x5               g136(.a(new_n231), .b(new_n229), .c(new_n219), .d(new_n230), .o1(new_n232));
  aoi022aa1n02x5               g137(.a(new_n228), .b(new_n229), .c(new_n222), .d(new_n232), .o1(\s[21] ));
  norp02aa1n02x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  nor042aa1n04x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  nanp02aa1n04x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  nanb02aa1n03x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n234), .c(new_n228), .d(new_n229), .o1(new_n238));
  xnrc02aa1n02x5               g143(.a(\b[20] ), .b(\a[21] ), .out0(new_n239));
  aoai13aa1n02x5               g144(.a(new_n236), .b(new_n239), .c(new_n222), .d(new_n227), .o1(new_n240));
  oai013aa1n02x4               g145(.a(new_n238), .b(new_n240), .c(new_n234), .d(new_n235), .o1(\s[22] ));
  nor042aa1n02x5               g146(.a(new_n239), .b(new_n237), .o1(new_n242));
  and003aa1n02x5               g147(.a(new_n203), .b(new_n242), .c(new_n219), .o(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n191), .c(new_n126), .d(new_n187), .o1(new_n244));
  nanb02aa1n06x5               g149(.a(new_n237), .b(new_n229), .out0(new_n245));
  aoi012aa1n09x5               g150(.a(new_n235), .b(new_n234), .c(new_n236), .o1(new_n246));
  aoai13aa1n12x5               g151(.a(new_n246), .b(new_n245), .c(new_n224), .d(new_n225), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  nanp02aa1n03x5               g153(.a(new_n244), .b(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  aoai13aa1n09x5               g155(.a(new_n242), .b(new_n231), .c(new_n219), .d(new_n230), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n250), .o1(new_n252));
  and003aa1n02x5               g157(.a(new_n251), .b(new_n252), .c(new_n246), .o(new_n253));
  aoi022aa1n02x5               g158(.a(new_n249), .b(new_n250), .c(new_n244), .d(new_n253), .o1(\s[23] ));
  norp02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  nor042aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nanp02aa1n02x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  nanb02aa1n02x5               g162(.a(new_n256), .b(new_n257), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n255), .c(new_n249), .d(new_n250), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n257), .b(new_n252), .c(new_n244), .d(new_n248), .o1(new_n260));
  oai013aa1n02x4               g165(.a(new_n259), .b(new_n260), .c(new_n255), .d(new_n256), .o1(\s[24] ));
  norb02aa1n03x5               g166(.a(new_n250), .b(new_n258), .out0(new_n262));
  inv030aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  nano32aa1n02x4               g168(.a(new_n263), .b(new_n203), .c(new_n242), .d(new_n219), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n191), .c(new_n126), .d(new_n187), .o1(new_n265));
  aoi012aa1n12x5               g170(.a(new_n256), .b(new_n255), .c(new_n257), .o1(new_n266));
  aoai13aa1n12x5               g171(.a(new_n266), .b(new_n263), .c(new_n251), .d(new_n246), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  nanp02aa1n03x5               g173(.a(new_n265), .b(new_n268), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  inv000aa1d42x5               g175(.a(new_n266), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(new_n270), .b(new_n271), .c(new_n247), .d(new_n262), .o1(new_n272));
  aoi022aa1n02x5               g177(.a(new_n269), .b(new_n270), .c(new_n265), .d(new_n272), .o1(\s[25] ));
  nor002aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  norp02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .o1(new_n275));
  nanp02aa1n02x5               g180(.a(\b[25] ), .b(\a[26] ), .o1(new_n276));
  nanb02aa1n02x5               g181(.a(new_n275), .b(new_n276), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n274), .c(new_n269), .d(new_n270), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n270), .o1(new_n279));
  aoai13aa1n02x5               g184(.a(new_n276), .b(new_n279), .c(new_n265), .d(new_n268), .o1(new_n280));
  oai013aa1n02x4               g185(.a(new_n278), .b(new_n280), .c(new_n274), .d(new_n275), .o1(\s[26] ));
  norb02aa1n03x5               g186(.a(new_n270), .b(new_n277), .out0(new_n282));
  nona23aa1n02x4               g187(.a(new_n250), .b(new_n229), .c(new_n258), .d(new_n237), .out0(new_n283));
  nano32aa1n02x5               g188(.a(new_n283), .b(new_n282), .c(new_n219), .d(new_n203), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n191), .c(new_n126), .d(new_n187), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n282), .b(new_n271), .c(new_n247), .d(new_n262), .o1(new_n286));
  aoi012aa1n02x5               g191(.a(new_n275), .b(new_n274), .c(new_n276), .o1(new_n287));
  nand23aa1n06x5               g192(.a(new_n285), .b(new_n286), .c(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  inv000aa1n02x5               g194(.a(new_n287), .o1(new_n290));
  aoi112aa1n02x5               g195(.a(new_n289), .b(new_n290), .c(new_n267), .d(new_n282), .o1(new_n291));
  aoi022aa1n02x5               g196(.a(new_n288), .b(new_n289), .c(new_n291), .d(new_n285), .o1(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  norp02aa1n02x5               g198(.a(\b[27] ), .b(\a[28] ), .o1(new_n294));
  nanp02aa1n02x5               g199(.a(\b[27] ), .b(\a[28] ), .o1(new_n295));
  nanb02aa1n02x5               g200(.a(new_n294), .b(new_n295), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n293), .c(new_n288), .d(new_n289), .o1(new_n297));
  oai022aa1n02x5               g202(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n298));
  aoi012aa1n09x5               g203(.a(new_n290), .b(new_n267), .c(new_n282), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n289), .o1(new_n300));
  aoai13aa1n02x5               g205(.a(new_n295), .b(new_n300), .c(new_n299), .d(new_n285), .o1(new_n301));
  oaih12aa1n02x5               g206(.a(new_n297), .b(new_n301), .c(new_n298), .o1(\s[28] ));
  norb02aa1n02x5               g207(.a(new_n289), .b(new_n296), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n288), .b(new_n303), .o1(new_n304));
  inv000aa1n03x5               g209(.a(new_n303), .o1(new_n305));
  and002aa1n02x5               g210(.a(\b[28] ), .b(\a[29] ), .o(new_n306));
  norp02aa1n02x5               g211(.a(\b[28] ), .b(\a[29] ), .o1(new_n307));
  aoi012aa1n02x5               g212(.a(new_n307), .b(new_n293), .c(new_n295), .o1(new_n308));
  norb03aa1n02x5               g213(.a(new_n308), .b(new_n294), .c(new_n306), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n299), .d(new_n285), .o1(new_n310));
  aoi012aa1n02x5               g215(.a(new_n294), .b(new_n293), .c(new_n295), .o1(new_n311));
  nor002aa1n02x5               g216(.a(new_n306), .b(new_n307), .o1(new_n312));
  aoai13aa1n03x5               g217(.a(new_n310), .b(new_n312), .c(new_n304), .d(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g219(.a(new_n296), .b(new_n289), .c(new_n312), .out0(new_n315));
  nanp02aa1n03x5               g220(.a(new_n288), .b(new_n315), .o1(new_n316));
  tech160nm_fioaoi03aa1n02p5x5 g221(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n317), .o1(new_n318));
  norp02aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .o1(new_n319));
  nanp02aa1n02x5               g224(.a(\b[29] ), .b(\a[30] ), .o1(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(new_n321));
  inv000aa1n02x5               g226(.a(new_n315), .o1(new_n322));
  nona22aa1n02x4               g227(.a(new_n320), .b(new_n319), .c(new_n307), .out0(new_n323));
  oab012aa1n02x4               g228(.a(new_n323), .b(new_n311), .c(new_n306), .out0(new_n324));
  aoai13aa1n02x5               g229(.a(new_n324), .b(new_n322), .c(new_n299), .d(new_n285), .o1(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n321), .c(new_n316), .d(new_n318), .o1(\s[30] ));
  nano22aa1n02x4               g231(.a(new_n305), .b(new_n312), .c(new_n321), .out0(new_n327));
  nanp02aa1n03x5               g232(.a(new_n288), .b(new_n327), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  inv000aa1n02x5               g234(.a(new_n327), .o1(new_n330));
  oai012aa1n02x5               g235(.a(new_n329), .b(\b[29] ), .c(\a[30] ), .o1(new_n331));
  aoi012aa1n02x5               g236(.a(new_n331), .b(new_n317), .c(new_n321), .o1(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n330), .c(new_n299), .d(new_n285), .o1(new_n333));
  aoi012aa1n02x5               g238(.a(new_n319), .b(new_n317), .c(new_n321), .o1(new_n334));
  aoai13aa1n03x5               g239(.a(new_n333), .b(new_n329), .c(new_n328), .d(new_n334), .o1(\s[31] ));
  nanp03aa1n02x5               g240(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n108), .b(new_n336), .c(new_n99), .out0(\s[3] ));
  aoi012aa1n02x5               g242(.a(new_n106), .b(new_n102), .c(new_n107), .o1(new_n338));
  xnrc02aa1n02x5               g243(.a(new_n338), .b(new_n105), .out0(\s[4] ));
  norb02aa1n02x5               g244(.a(new_n114), .b(new_n113), .out0(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n340), .b(new_n109), .c(new_n110), .out0(\s[5] ));
  nanp02aa1n02x5               g246(.a(new_n109), .b(new_n110), .o1(new_n342));
  aoi012aa1n02x5               g247(.a(new_n113), .b(new_n342), .c(new_n114), .o1(new_n343));
  xnrb03aa1n02x5               g248(.a(new_n343), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g249(.a(new_n119), .b(new_n118), .out0(new_n345));
  aobi12aa1n02x5               g250(.a(new_n115), .b(new_n109), .c(new_n110), .out0(new_n346));
  oa0012aa1n02x5               g251(.a(new_n345), .b(new_n346), .c(new_n123), .o(new_n347));
  aoi112aa1n02x5               g252(.a(new_n123), .b(new_n345), .c(new_n342), .d(new_n115), .o1(new_n348));
  norp02aa1n02x5               g253(.a(new_n347), .b(new_n348), .o1(\s[7] ));
  oaoi13aa1n02x5               g254(.a(new_n118), .b(new_n119), .c(new_n346), .d(new_n123), .o1(new_n350));
  xnrb03aa1n02x5               g255(.a(new_n350), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  inv000aa1d42x5               g256(.a(new_n146), .o1(new_n352));
  aoi112aa1n02x5               g257(.a(new_n352), .b(new_n124), .c(new_n120), .d(new_n123), .o1(new_n353));
  aoai13aa1n02x5               g258(.a(new_n353), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n354));
  aob012aa1n02x5               g259(.a(new_n354), .b(new_n126), .c(new_n352), .out0(\s[9] ));
endmodule


