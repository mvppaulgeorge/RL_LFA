// Benchmark "adder" written by ABC on Thu Jul 11 11:57:14 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n321, new_n322, new_n324, new_n325, new_n327, new_n328,
    new_n329, new_n330;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  norp02aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  160nm_ficinv00aa1n08x5       g005(.clk(new_n100), .clkout(new_n101));
  nanp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oai012aa1n02x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  norp02aa1n02x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n02x4               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  aoi012aa1n02x5               g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1n02x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  norp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .out0(new_n118));
  xnrc02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .out0(new_n119));
  norp03aa1n02x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  oai012aa1n02x5               g025(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n121));
  160nm_ficinv00aa1n08x5       g026(.clk(\b[5] ), .clkout(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  oaib12aa1n02x5               g028(.a(new_n123), .b(new_n122), .c(\a[6] ), .out0(new_n124));
  oai012aa1n02x5               g029(.a(new_n121), .b(new_n117), .c(new_n124), .o1(new_n125));
  nanp02aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n100), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n112), .d(new_n120), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n99), .b(new_n128), .c(new_n101), .out0(\s[10] ));
  aobi12aa1n02x5               g034(.a(new_n99), .b(new_n128), .c(new_n101), .out0(new_n130));
  norp02aa1n02x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  oaoi03aa1n02x5               g038(.a(\a[10] ), .b(\b[9] ), .c(new_n101), .o1(new_n134));
  oai012aa1n02x5               g039(.a(new_n133), .b(new_n130), .c(new_n134), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n131), .b(new_n132), .out0(new_n136));
  oai012aa1n02x5               g041(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n137));
  nano22aa1n02x4               g042(.a(new_n130), .b(new_n136), .c(new_n137), .out0(new_n138));
  norb02aa1n02x5               g043(.a(new_n135), .b(new_n138), .out0(\s[11] ));
  norp02aa1n02x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  nona22aa1n02x4               g047(.a(new_n135), .b(new_n142), .c(new_n131), .out0(new_n143));
  nanb02aa1n02x5               g048(.a(new_n140), .b(new_n141), .out0(new_n144));
  oaoi13aa1n02x5               g049(.a(new_n144), .b(new_n135), .c(\a[11] ), .d(\b[10] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n143), .b(new_n145), .out0(\s[12] ));
  nano23aa1n02x4               g051(.a(new_n97), .b(new_n100), .c(new_n126), .d(new_n98), .out0(new_n147));
  nona22aa1n02x4               g052(.a(new_n147), .b(new_n144), .c(new_n136), .out0(new_n148));
  160nm_ficinv00aa1n08x5       g053(.clk(new_n148), .clkout(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n125), .c(new_n112), .d(new_n120), .o1(new_n150));
  nona23aa1n02x4               g055(.a(new_n141), .b(new_n132), .c(new_n131), .d(new_n140), .out0(new_n151));
  aoi012aa1n02x5               g056(.a(new_n140), .b(new_n131), .c(new_n141), .o1(new_n152));
  oai012aa1n02x5               g057(.a(new_n152), .b(new_n151), .c(new_n137), .o1(new_n153));
  160nm_ficinv00aa1n08x5       g058(.clk(new_n153), .clkout(new_n154));
  norp02aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n150), .c(new_n154), .out0(\s[13] ));
  160nm_ficinv00aa1n08x5       g063(.clk(\a[13] ), .clkout(new_n159));
  160nm_ficinv00aa1n08x5       g064(.clk(\b[12] ), .clkout(new_n160));
  nanp02aa1n02x5               g065(.a(new_n150), .b(new_n154), .o1(new_n161));
  oaoi03aa1n02x5               g066(.a(new_n159), .b(new_n160), .c(new_n161), .o1(new_n162));
  norp02aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  xnrc02aa1n02x5               g070(.a(new_n162), .b(new_n165), .out0(\s[14] ));
  nona23aa1n02x4               g071(.a(new_n164), .b(new_n156), .c(new_n155), .d(new_n163), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n164), .b(new_n163), .c(new_n159), .d(new_n160), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n167), .c(new_n150), .d(new_n154), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  160nm_ficinv00aa1n08x5       g075(.clk(\a[15] ), .clkout(new_n171));
  160nm_ficinv00aa1n08x5       g076(.clk(\b[14] ), .clkout(new_n172));
  oaoi03aa1n02x5               g077(.a(new_n171), .b(new_n172), .c(new_n169), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  160nm_ficinv00aa1n08x5       g079(.clk(new_n174), .clkout(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n173), .b(new_n176), .c(new_n175), .out0(\s[16] ));
  norp02aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nano23aa1n02x4               g084(.a(new_n178), .b(new_n174), .c(new_n176), .d(new_n179), .out0(new_n180));
  nanp03aa1n02x5               g085(.a(new_n180), .b(new_n157), .c(new_n165), .o1(new_n181));
  norp02aa1n02x5               g086(.a(new_n181), .b(new_n148), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n125), .c(new_n112), .d(new_n120), .o1(new_n183));
  nanb02aa1n02x5               g088(.a(new_n168), .b(new_n180), .out0(new_n184));
  aoi112aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n185));
  160nm_ficinv00aa1n08x5       g090(.clk(new_n185), .clkout(new_n186));
  nanp03aa1n02x5               g091(.a(new_n134), .b(new_n133), .c(new_n142), .o1(new_n187));
  aoi012aa1n02x5               g092(.a(new_n181), .b(new_n187), .c(new_n152), .o1(new_n188));
  nano32aa1n02x4               g093(.a(new_n188), .b(new_n186), .c(new_n184), .d(new_n175), .out0(new_n189));
  nanp02aa1n02x5               g094(.a(new_n189), .b(new_n183), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g096(.clk(\a[18] ), .clkout(new_n192));
  160nm_ficinv00aa1n08x5       g097(.clk(\a[17] ), .clkout(new_n193));
  160nm_ficinv00aa1n08x5       g098(.clk(\b[16] ), .clkout(new_n194));
  oaoi03aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d04x5               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  nanp02aa1n02x5               g102(.a(new_n194), .b(new_n193), .o1(new_n198));
  oaoi03aa1n02x5               g103(.a(\a[18] ), .b(\b[17] ), .c(new_n198), .o1(new_n199));
  norp02aa1n02x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  aoai13aa1n02x5               g107(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n197), .o1(new_n203));
  aoi112aa1n02x5               g108(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n197), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  nona22aa1n02x4               g114(.a(new_n203), .b(new_n209), .c(new_n200), .out0(new_n210));
  160nm_ficinv00aa1n08x5       g115(.clk(new_n200), .clkout(new_n211));
  aobi12aa1n02x5               g116(.a(new_n209), .b(new_n203), .c(new_n211), .out0(new_n212));
  norb02aa1n02x5               g117(.a(new_n210), .b(new_n212), .out0(\s[20] ));
  nano23aa1n02x4               g118(.a(new_n200), .b(new_n207), .c(new_n208), .d(new_n201), .out0(new_n214));
  nanp02aa1n02x5               g119(.a(new_n197), .b(new_n214), .o1(new_n215));
  oai022aa1n02x5               g120(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n216));
  oaib12aa1n02x5               g121(.a(new_n216), .b(new_n192), .c(\b[17] ), .out0(new_n217));
  nona23aa1n02x4               g122(.a(new_n208), .b(new_n201), .c(new_n200), .d(new_n207), .out0(new_n218));
  aoi012aa1n02x5               g123(.a(new_n207), .b(new_n200), .c(new_n208), .o1(new_n219));
  oai012aa1n02x5               g124(.a(new_n219), .b(new_n218), .c(new_n217), .o1(new_n220));
  160nm_ficinv00aa1n08x5       g125(.clk(new_n220), .clkout(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n215), .c(new_n189), .d(new_n183), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xorc02aa1n02x5               g130(.a(\a[22] ), .b(\b[21] ), .out0(new_n226));
  aoi112aa1n02x5               g131(.a(new_n224), .b(new_n226), .c(new_n222), .d(new_n225), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n226), .b(new_n224), .c(new_n222), .d(new_n225), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(\s[22] ));
  160nm_ficinv00aa1n08x5       g134(.clk(\a[21] ), .clkout(new_n230));
  160nm_ficinv00aa1n08x5       g135(.clk(\a[22] ), .clkout(new_n231));
  xroi22aa1d04x5               g136(.a(new_n230), .b(\b[20] ), .c(new_n231), .d(\b[21] ), .out0(new_n232));
  nanp03aa1n02x5               g137(.a(new_n232), .b(new_n197), .c(new_n214), .o1(new_n233));
  160nm_ficinv00aa1n08x5       g138(.clk(\b[21] ), .clkout(new_n234));
  oaoi03aa1n02x5               g139(.a(new_n231), .b(new_n234), .c(new_n224), .o1(new_n235));
  160nm_ficinv00aa1n08x5       g140(.clk(new_n235), .clkout(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n220), .c(new_n232), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n233), .c(new_n189), .d(new_n183), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  xorc02aa1n02x5               g145(.a(\a[23] ), .b(\b[22] ), .out0(new_n241));
  xorc02aa1n02x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  aoi112aa1n02x5               g147(.a(new_n240), .b(new_n242), .c(new_n238), .d(new_n241), .o1(new_n243));
  aoai13aa1n02x5               g148(.a(new_n242), .b(new_n240), .c(new_n238), .d(new_n241), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n244), .b(new_n243), .out0(\s[24] ));
  and002aa1n02x5               g150(.a(new_n242), .b(new_n241), .o(new_n246));
  160nm_ficinv00aa1n08x5       g151(.clk(new_n246), .clkout(new_n247));
  nano32aa1n02x4               g152(.a(new_n247), .b(new_n232), .c(new_n197), .d(new_n214), .out0(new_n248));
  160nm_ficinv00aa1n08x5       g153(.clk(new_n219), .clkout(new_n249));
  aoai13aa1n02x5               g154(.a(new_n232), .b(new_n249), .c(new_n214), .d(new_n199), .o1(new_n250));
  norp02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  aoi012aa1n02x5               g157(.a(new_n251), .b(new_n240), .c(new_n252), .o1(new_n253));
  aoai13aa1n02x5               g158(.a(new_n253), .b(new_n247), .c(new_n250), .d(new_n235), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  aoai13aa1n02x5               g160(.a(new_n255), .b(new_n254), .c(new_n190), .d(new_n248), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n255), .b(new_n254), .c(new_n190), .d(new_n248), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n256), .b(new_n257), .out0(\s[25] ));
  norp02aa1n02x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  xorc02aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .out0(new_n260));
  nona22aa1n02x4               g165(.a(new_n256), .b(new_n260), .c(new_n259), .out0(new_n261));
  160nm_ficinv00aa1n08x5       g166(.clk(new_n259), .clkout(new_n262));
  aobi12aa1n02x5               g167(.a(new_n260), .b(new_n256), .c(new_n262), .out0(new_n263));
  norb02aa1n02x5               g168(.a(new_n261), .b(new_n263), .out0(\s[26] ));
  nanp02aa1n02x5               g169(.a(new_n112), .b(new_n120), .o1(new_n265));
  160nm_ficinv00aa1n08x5       g170(.clk(new_n125), .clkout(new_n266));
  nanp02aa1n02x5               g171(.a(new_n265), .b(new_n266), .o1(new_n267));
  nanb02aa1n02x5               g172(.a(new_n178), .b(new_n179), .out0(new_n268));
  nanb02aa1n02x5               g173(.a(new_n174), .b(new_n176), .out0(new_n269));
  norp03aa1n02x5               g174(.a(new_n168), .b(new_n269), .c(new_n268), .o1(new_n270));
  nona32aa1n02x4               g175(.a(new_n153), .b(new_n269), .c(new_n167), .d(new_n268), .out0(new_n271));
  nona32aa1n02x4               g176(.a(new_n271), .b(new_n185), .c(new_n270), .d(new_n174), .out0(new_n272));
  and002aa1n02x5               g177(.a(new_n260), .b(new_n255), .o(new_n273));
  nano22aa1n02x4               g178(.a(new_n233), .b(new_n246), .c(new_n273), .out0(new_n274));
  aoai13aa1n02x5               g179(.a(new_n274), .b(new_n272), .c(new_n267), .d(new_n182), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .c(new_n262), .carry(new_n276));
  aobi12aa1n02x5               g181(.a(new_n276), .b(new_n254), .c(new_n273), .out0(new_n277));
  xorc02aa1n02x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n277), .c(new_n275), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  160nm_ficinv00aa1n08x5       g185(.clk(new_n280), .clkout(new_n281));
  aobi12aa1n02x5               g186(.a(new_n278), .b(new_n277), .c(new_n275), .out0(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  nano22aa1n02x4               g188(.a(new_n282), .b(new_n281), .c(new_n283), .out0(new_n284));
  aobi12aa1n02x5               g189(.a(new_n274), .b(new_n189), .c(new_n183), .out0(new_n285));
  aoai13aa1n02x5               g190(.a(new_n246), .b(new_n236), .c(new_n220), .d(new_n232), .o1(new_n286));
  160nm_ficinv00aa1n08x5       g191(.clk(new_n273), .clkout(new_n287));
  aoai13aa1n02x5               g192(.a(new_n276), .b(new_n287), .c(new_n286), .d(new_n253), .o1(new_n288));
  oai012aa1n02x5               g193(.a(new_n278), .b(new_n288), .c(new_n285), .o1(new_n289));
  aoi012aa1n02x5               g194(.a(new_n283), .b(new_n289), .c(new_n281), .o1(new_n290));
  norp02aa1n02x5               g195(.a(new_n290), .b(new_n284), .o1(\s[28] ));
  norb02aa1n02x5               g196(.a(new_n278), .b(new_n283), .out0(new_n292));
  oai012aa1n02x5               g197(.a(new_n292), .b(new_n288), .c(new_n285), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n281), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  aoi012aa1n02x5               g200(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n296));
  aobi12aa1n02x5               g201(.a(new_n292), .b(new_n277), .c(new_n275), .out0(new_n297));
  nano22aa1n02x4               g202(.a(new_n297), .b(new_n294), .c(new_n295), .out0(new_n298));
  norp02aa1n02x5               g203(.a(new_n296), .b(new_n298), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g205(.a(new_n278), .b(new_n295), .c(new_n283), .out0(new_n301));
  oai012aa1n02x5               g206(.a(new_n301), .b(new_n288), .c(new_n285), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[29] ), .b(\a[30] ), .out0(new_n304));
  aoi012aa1n02x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  aobi12aa1n02x5               g210(.a(new_n301), .b(new_n277), .c(new_n275), .out0(new_n306));
  nano22aa1n02x4               g211(.a(new_n306), .b(new_n303), .c(new_n304), .out0(new_n307));
  norp02aa1n02x5               g212(.a(new_n305), .b(new_n307), .o1(\s[30] ));
  xnrc02aa1n02x5               g213(.a(\b[30] ), .b(\a[31] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n301), .b(new_n304), .out0(new_n310));
  aobi12aa1n02x5               g215(.a(new_n310), .b(new_n277), .c(new_n275), .out0(new_n311));
  oao003aa1n02x5               g216(.a(\a[30] ), .b(\b[29] ), .c(new_n303), .carry(new_n312));
  nano22aa1n02x4               g217(.a(new_n311), .b(new_n309), .c(new_n312), .out0(new_n313));
  oai012aa1n02x5               g218(.a(new_n310), .b(new_n288), .c(new_n285), .o1(new_n314));
  aoi012aa1n02x5               g219(.a(new_n309), .b(new_n314), .c(new_n312), .o1(new_n315));
  norp02aa1n02x5               g220(.a(new_n315), .b(new_n313), .o1(\s[31] ));
  xnrb03aa1n02x5               g221(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g222(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g224(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g225(.a(new_n119), .b(new_n112), .out0(new_n321));
  oai012aa1n02x5               g226(.a(new_n321), .b(\b[4] ), .c(\a[5] ), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g228(.a(new_n118), .b(new_n322), .out0(new_n324));
  oaib12aa1n02x5               g229(.a(new_n324), .b(\a[6] ), .c(new_n122), .out0(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g231(.a(new_n113), .b(new_n114), .out0(new_n327));
  160nm_ficinv00aa1n08x5       g232(.clk(new_n327), .clkout(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n115), .c(new_n325), .d(new_n116), .o1(new_n329));
  aoi112aa1n02x5               g234(.a(new_n328), .b(new_n115), .c(new_n325), .d(new_n116), .o1(new_n330));
  norb02aa1n02x5               g235(.a(new_n329), .b(new_n330), .out0(\s[8] ));
  xnbna2aa1n03x5               g236(.a(new_n127), .b(new_n265), .c(new_n266), .out0(\s[9] ));
endmodule


