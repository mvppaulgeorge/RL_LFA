// Benchmark "adder" written by ABC on Thu Jul 18 12:28:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n350, new_n351,
    new_n352, new_n354, new_n355, new_n357, new_n359, new_n360, new_n361,
    new_n362, new_n364, new_n365, new_n367, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nand02aa1d28x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n02x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor022aa1n06x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1n03x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1d32x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n03x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  tech160nm_fioai012aa1n05x5   g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oai012aa1n04x7               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand02aa1n08x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  norp02aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nona23aa1n02x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .d(new_n110), .out0(new_n114));
  xnrc02aa1n12x5               g019(.a(\b[4] ), .b(\a[5] ), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  nor043aa1n03x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  inv000aa1d42x5               g022(.a(new_n110), .o1(new_n118));
  inv000aa1d42x5               g023(.a(new_n112), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[8] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[7] ), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  norp02aa1n06x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  nor002aa1n02x5               g028(.a(\b[5] ), .b(\a[6] ), .o1(new_n124));
  aoi022aa1n09x5               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  oai012aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n123), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n122), .b(new_n119), .c(new_n126), .d(new_n118), .o1(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n127), .c(new_n109), .d(new_n117), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  oai022aa1d24x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n131), .b(new_n129), .out0(new_n132));
  nand02aa1d08x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1n10x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  tech160nm_fioai012aa1n04x5   g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .o1(new_n135));
  nanb03aa1n06x5               g040(.a(new_n135), .b(new_n132), .c(new_n133), .out0(new_n136));
  orn002aa1n02x5               g041(.a(\a[11] ), .b(\b[10] ), .o(new_n137));
  aoi022aa1n02x5               g042(.a(new_n132), .b(new_n134), .c(new_n137), .d(new_n133), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n136), .b(new_n138), .out0(\s[11] ));
  tech160nm_fixorc02aa1n03p5x5 g044(.a(\a[12] ), .b(\b[11] ), .out0(new_n140));
  oai022aa1n03x5               g045(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n141));
  aoi012aa1n06x5               g046(.a(new_n141), .b(\a[12] ), .c(\b[11] ), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(new_n136), .b(new_n142), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n140), .c(new_n136), .d(new_n137), .o1(\s[12] ));
  inv000aa1n03x5               g049(.a(new_n101), .o1(new_n145));
  oaoi03aa1n02x5               g050(.a(\a[2] ), .b(\b[1] ), .c(new_n145), .o1(new_n146));
  norb02aa1n06x5               g051(.a(new_n104), .b(new_n103), .out0(new_n147));
  norb02aa1n09x5               g052(.a(new_n106), .b(new_n105), .out0(new_n148));
  nand23aa1n04x5               g053(.a(new_n146), .b(new_n147), .c(new_n148), .o1(new_n149));
  nano23aa1n02x4               g054(.a(new_n113), .b(new_n110), .c(new_n111), .d(new_n112), .out0(new_n150));
  nona22aa1n02x4               g055(.a(new_n150), .b(new_n115), .c(new_n116), .out0(new_n151));
  nand02aa1n04x5               g056(.a(new_n126), .b(new_n118), .o1(new_n152));
  oaoi03aa1n09x5               g057(.a(new_n120), .b(new_n121), .c(new_n152), .o1(new_n153));
  aoai13aa1n09x5               g058(.a(new_n153), .b(new_n151), .c(new_n149), .d(new_n108), .o1(new_n154));
  nand23aa1n04x5               g059(.a(new_n131), .b(new_n134), .c(new_n133), .o1(new_n155));
  aob012aa1n06x5               g060(.a(new_n133), .b(\b[8] ), .c(\a[9] ), .out0(new_n156));
  nona23aa1n09x5               g061(.a(new_n155), .b(new_n140), .c(new_n156), .d(new_n135), .out0(new_n157));
  nanb02aa1n02x5               g062(.a(new_n157), .b(new_n154), .out0(new_n158));
  inv000aa1d42x5               g063(.a(\b[11] ), .o1(new_n159));
  nand42aa1n02x5               g064(.a(new_n155), .b(new_n142), .o1(new_n160));
  oaib12aa1n02x5               g065(.a(new_n160), .b(new_n159), .c(\a[12] ), .out0(new_n161));
  nor022aa1n12x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand02aa1n06x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n158), .c(new_n161), .out0(\s[13] ));
  inv000aa1d42x5               g070(.a(new_n162), .o1(new_n166));
  nanp02aa1n03x5               g071(.a(new_n109), .b(new_n117), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n161), .b(new_n157), .c(new_n167), .d(new_n153), .o1(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n164), .o1(new_n169));
  nor002aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand02aa1n10x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  oaih22aa1d12x5               g077(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n173));
  nanb03aa1n02x5               g078(.a(new_n173), .b(new_n169), .c(new_n171), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n172), .c(new_n166), .d(new_n169), .o1(\s[14] ));
  nano23aa1n06x5               g080(.a(new_n162), .b(new_n170), .c(new_n171), .d(new_n163), .out0(new_n176));
  oaoi03aa1n02x5               g081(.a(\a[14] ), .b(\b[13] ), .c(new_n166), .o1(new_n177));
  tech160nm_fixorc02aa1n03p5x5 g082(.a(\a[15] ), .b(\b[14] ), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n177), .c(new_n168), .d(new_n176), .o1(new_n179));
  aoi112aa1n02x5               g084(.a(new_n178), .b(new_n177), .c(new_n168), .d(new_n176), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(\a[15] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[14] ), .o1(new_n183));
  nand22aa1n02x5               g088(.a(new_n183), .b(new_n182), .o1(new_n184));
  norp02aa1n04x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  and002aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o(new_n186));
  nor002aa1n02x5               g091(.a(new_n186), .b(new_n185), .o1(new_n187));
  oai022aa1n02x5               g092(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n188));
  nona22aa1n03x5               g093(.a(new_n179), .b(new_n186), .c(new_n188), .out0(new_n189));
  aoai13aa1n02x5               g094(.a(new_n189), .b(new_n187), .c(new_n184), .d(new_n179), .o1(\s[16] ));
  nano32aa1n03x7               g095(.a(new_n157), .b(new_n187), .c(new_n176), .d(new_n178), .out0(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n127), .c(new_n109), .d(new_n117), .o1(new_n192));
  aoi112aa1n03x5               g097(.a(new_n186), .b(new_n185), .c(\a[15] ), .d(\b[14] ), .o1(new_n193));
  obai22aa1n02x7               g098(.a(\a[12] ), .b(new_n159), .c(\b[12] ), .d(\a[13] ), .out0(new_n194));
  oai012aa1n02x5               g099(.a(new_n163), .b(\b[13] ), .c(\a[14] ), .o1(new_n195));
  nano23aa1n06x5               g100(.a(new_n194), .b(new_n195), .c(new_n184), .d(new_n171), .out0(new_n196));
  oai112aa1n02x5               g101(.a(new_n173), .b(new_n171), .c(new_n183), .d(new_n182), .o1(new_n197));
  aoi022aa1n03x5               g102(.a(new_n197), .b(new_n184), .c(\a[16] ), .d(\b[15] ), .o1(new_n198));
  aoi113aa1n09x5               g103(.a(new_n198), .b(new_n185), .c(new_n160), .d(new_n196), .e(new_n193), .o1(new_n199));
  nanp02aa1n09x5               g104(.a(new_n192), .b(new_n199), .o1(new_n200));
  nor042aa1n09x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  nand42aa1n03x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  obai22aa1n02x7               g108(.a(new_n202), .b(new_n201), .c(\a[16] ), .d(\b[15] ), .out0(new_n204));
  aoi113aa1n02x5               g109(.a(new_n198), .b(new_n204), .c(new_n160), .d(new_n196), .e(new_n193), .o1(new_n205));
  aoi022aa1n02x5               g110(.a(new_n200), .b(new_n203), .c(new_n192), .d(new_n205), .o1(\s[17] ));
  inv000aa1d42x5               g111(.a(new_n201), .o1(new_n207));
  nanp03aa1n02x5               g112(.a(new_n160), .b(new_n196), .c(new_n193), .o1(new_n208));
  nona22aa1n02x4               g113(.a(new_n208), .b(new_n198), .c(new_n185), .out0(new_n209));
  aoai13aa1n02x5               g114(.a(new_n203), .b(new_n209), .c(new_n154), .d(new_n191), .o1(new_n210));
  nor042aa1n02x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nand42aa1n04x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  oaih22aa1n04x5               g118(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n214));
  nanb03aa1n02x5               g119(.a(new_n214), .b(new_n210), .c(new_n212), .out0(new_n215));
  aoai13aa1n02x5               g120(.a(new_n215), .b(new_n213), .c(new_n207), .d(new_n210), .o1(\s[18] ));
  nano23aa1n06x5               g121(.a(new_n201), .b(new_n211), .c(new_n212), .d(new_n202), .out0(new_n217));
  oaoi03aa1n02x5               g122(.a(\a[18] ), .b(\b[17] ), .c(new_n207), .o1(new_n218));
  nor002aa1d32x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  nand42aa1n02x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  norb02aa1n03x5               g125(.a(new_n220), .b(new_n219), .out0(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n218), .c(new_n200), .d(new_n217), .o1(new_n222));
  aoi112aa1n02x5               g127(.a(new_n221), .b(new_n218), .c(new_n200), .d(new_n217), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n222), .b(new_n223), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g130(.a(new_n219), .o1(new_n226));
  nor002aa1n06x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  tech160nm_finand02aa1n03p5x5 g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  norb02aa1n03x5               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  norb03aa1n02x5               g134(.a(new_n228), .b(new_n219), .c(new_n227), .out0(new_n230));
  nanp02aa1n03x5               g135(.a(new_n222), .b(new_n230), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n229), .c(new_n226), .d(new_n222), .o1(\s[20] ));
  nand03aa1n06x5               g137(.a(new_n217), .b(new_n221), .c(new_n229), .o1(new_n233));
  inv040aa1n03x5               g138(.a(new_n233), .o1(new_n234));
  tech160nm_fioai012aa1n03p5x5 g139(.a(new_n228), .b(new_n227), .c(new_n219), .o1(new_n235));
  nanb03aa1n02x5               g140(.a(new_n227), .b(new_n228), .c(new_n220), .out0(new_n236));
  oai112aa1n02x5               g141(.a(new_n214), .b(new_n212), .c(\b[18] ), .d(\a[19] ), .o1(new_n237));
  oai012aa1n04x7               g142(.a(new_n235), .b(new_n237), .c(new_n236), .o1(new_n238));
  nor042aa1n06x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  nand02aa1n03x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n238), .c(new_n200), .d(new_n234), .o1(new_n242));
  inv000aa1n06x5               g147(.a(new_n235), .o1(new_n243));
  nano22aa1n03x5               g148(.a(new_n227), .b(new_n220), .c(new_n228), .out0(new_n244));
  oai012aa1n02x7               g149(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .o1(new_n245));
  oab012aa1n06x5               g150(.a(new_n245), .b(new_n201), .c(new_n211), .out0(new_n246));
  aoi112aa1n02x5               g151(.a(new_n241), .b(new_n243), .c(new_n246), .d(new_n244), .o1(new_n247));
  aobi12aa1n02x5               g152(.a(new_n247), .b(new_n200), .c(new_n234), .out0(new_n248));
  norb02aa1n03x4               g153(.a(new_n242), .b(new_n248), .out0(\s[21] ));
  inv020aa1n02x5               g154(.a(new_n239), .o1(new_n250));
  nor042aa1n02x5               g155(.a(\b[21] ), .b(\a[22] ), .o1(new_n251));
  nand02aa1n03x5               g156(.a(\b[21] ), .b(\a[22] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  norb03aa1n02x5               g158(.a(new_n252), .b(new_n239), .c(new_n251), .out0(new_n254));
  nanp02aa1n03x5               g159(.a(new_n242), .b(new_n254), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n253), .c(new_n250), .d(new_n242), .o1(\s[22] ));
  nano23aa1d15x5               g161(.a(new_n239), .b(new_n251), .c(new_n252), .d(new_n240), .out0(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  nano32aa1n02x4               g163(.a(new_n258), .b(new_n217), .c(new_n221), .d(new_n229), .out0(new_n259));
  aoai13aa1n06x5               g164(.a(new_n257), .b(new_n243), .c(new_n246), .d(new_n244), .o1(new_n260));
  oaoi03aa1n12x5               g165(.a(\a[22] ), .b(\b[21] ), .c(new_n250), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(new_n260), .b(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n263), .c(new_n200), .d(new_n259), .o1(new_n265));
  nona22aa1n02x4               g170(.a(new_n260), .b(new_n261), .c(new_n264), .out0(new_n266));
  aoi012aa1n02x5               g171(.a(new_n266), .b(new_n200), .c(new_n259), .o1(new_n267));
  norb02aa1n02x5               g172(.a(new_n265), .b(new_n267), .out0(\s[23] ));
  norp02aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[24] ), .b(\b[23] ), .out0(new_n271));
  oai022aa1n02x5               g176(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n272));
  aoi012aa1n02x5               g177(.a(new_n272), .b(\a[24] ), .c(\b[23] ), .o1(new_n273));
  nanp02aa1n03x5               g178(.a(new_n265), .b(new_n273), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n271), .c(new_n270), .d(new_n265), .o1(\s[24] ));
  nano32aa1n02x5               g180(.a(new_n233), .b(new_n271), .c(new_n257), .d(new_n264), .out0(new_n276));
  nanp02aa1n02x5               g181(.a(new_n271), .b(new_n264), .o1(new_n277));
  aob012aa1n02x5               g182(.a(new_n272), .b(\b[23] ), .c(\a[24] ), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n260), .d(new_n262), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[25] ), .b(\b[24] ), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n279), .c(new_n200), .d(new_n276), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n277), .o1(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n261), .c(new_n238), .d(new_n257), .o1(new_n283));
  nanb03aa1n02x5               g188(.a(new_n280), .b(new_n283), .c(new_n278), .out0(new_n284));
  aoi012aa1n02x5               g189(.a(new_n284), .b(new_n200), .c(new_n276), .o1(new_n285));
  norb02aa1n02x5               g190(.a(new_n281), .b(new_n285), .out0(\s[25] ));
  norp02aa1n02x5               g191(.a(\b[24] ), .b(\a[25] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  tech160nm_fixorc02aa1n02p5x5 g193(.a(\a[26] ), .b(\b[25] ), .out0(new_n289));
  nanp02aa1n02x5               g194(.a(\b[25] ), .b(\a[26] ), .o1(new_n290));
  oai022aa1n02x5               g195(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n291));
  norb02aa1n02x5               g196(.a(new_n290), .b(new_n291), .out0(new_n292));
  nanp02aa1n03x5               g197(.a(new_n281), .b(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n288), .d(new_n281), .o1(\s[26] ));
  nand02aa1d04x5               g199(.a(new_n289), .b(new_n280), .o1(new_n295));
  nano23aa1n06x5               g200(.a(new_n233), .b(new_n295), .c(new_n282), .d(new_n257), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n209), .c(new_n154), .d(new_n191), .o1(new_n297));
  nona32aa1n03x5               g202(.a(new_n234), .b(new_n295), .c(new_n277), .d(new_n258), .out0(new_n298));
  tech160nm_fiaoi012aa1n05x5   g203(.a(new_n298), .b(new_n192), .c(new_n199), .o1(new_n299));
  nanp02aa1n02x5               g204(.a(new_n291), .b(new_n290), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n295), .c(new_n283), .d(new_n278), .o1(new_n301));
  xorc02aa1n12x5               g206(.a(\a[27] ), .b(\b[26] ), .out0(new_n302));
  tech160nm_fioai012aa1n03p5x5 g207(.a(new_n302), .b(new_n301), .c(new_n299), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n295), .o1(new_n304));
  aoi122aa1n02x5               g209(.a(new_n302), .b(new_n290), .c(new_n291), .d(new_n279), .e(new_n304), .o1(new_n305));
  aobi12aa1n02x7               g210(.a(new_n303), .b(new_n305), .c(new_n297), .out0(\s[27] ));
  norp02aa1n02x5               g211(.a(\b[26] ), .b(\a[27] ), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[28] ), .b(\b[27] ), .out0(new_n309));
  aoi022aa1n06x5               g214(.a(new_n279), .b(new_n304), .c(new_n290), .d(new_n291), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n302), .o1(new_n311));
  nanp02aa1n02x5               g216(.a(\b[27] ), .b(\a[28] ), .o1(new_n312));
  oai022aa1d18x5               g217(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n313));
  norb02aa1n02x5               g218(.a(new_n312), .b(new_n313), .out0(new_n314));
  aoai13aa1n04x5               g219(.a(new_n314), .b(new_n311), .c(new_n310), .d(new_n297), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n309), .c(new_n303), .d(new_n308), .o1(\s[28] ));
  and002aa1n02x5               g221(.a(new_n309), .b(new_n302), .o(new_n317));
  oaih12aa1n02x5               g222(.a(new_n317), .b(new_n301), .c(new_n299), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  nanp02aa1n02x5               g224(.a(new_n313), .b(new_n312), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n319), .c(new_n310), .d(new_n297), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .out0(new_n322));
  aoi012aa1n02x5               g227(.a(new_n322), .b(new_n312), .c(new_n313), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g230(.a(new_n311), .b(new_n309), .c(new_n322), .out0(new_n326));
  oai012aa1n02x5               g231(.a(new_n326), .b(new_n301), .c(new_n299), .o1(new_n327));
  inv000aa1n02x5               g232(.a(new_n326), .o1(new_n328));
  inv000aa1d42x5               g233(.a(\a[29] ), .o1(new_n329));
  inv000aa1d42x5               g234(.a(\b[28] ), .o1(new_n330));
  nanp02aa1n02x5               g235(.a(new_n330), .b(new_n329), .o1(new_n331));
  oai112aa1n02x5               g236(.a(new_n313), .b(new_n312), .c(new_n330), .d(new_n329), .o1(new_n332));
  nanp02aa1n02x5               g237(.a(new_n332), .b(new_n331), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n333), .o1(new_n334));
  aoai13aa1n02x7               g239(.a(new_n334), .b(new_n328), .c(new_n310), .d(new_n297), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[30] ), .b(\b[29] ), .out0(new_n336));
  nano22aa1n02x4               g241(.a(new_n336), .b(new_n332), .c(new_n331), .out0(new_n337));
  aoi022aa1n03x5               g242(.a(new_n335), .b(new_n336), .c(new_n327), .d(new_n337), .o1(\s[30] ));
  nano32aa1n03x7               g243(.a(new_n311), .b(new_n336), .c(new_n309), .d(new_n322), .out0(new_n339));
  tech160nm_fioai012aa1n04x5   g244(.a(new_n339), .b(new_n301), .c(new_n299), .o1(new_n340));
  inv000aa1d42x5               g245(.a(new_n339), .o1(new_n341));
  inv000aa1d42x5               g246(.a(\a[30] ), .o1(new_n342));
  inv000aa1d42x5               g247(.a(\b[29] ), .o1(new_n343));
  oaoi03aa1n02x5               g248(.a(new_n342), .b(new_n343), .c(new_n333), .o1(new_n344));
  aoai13aa1n03x5               g249(.a(new_n344), .b(new_n341), .c(new_n310), .d(new_n297), .o1(new_n345));
  xorc02aa1n02x5               g250(.a(\a[31] ), .b(\b[30] ), .out0(new_n346));
  aoi022aa1n02x5               g251(.a(new_n332), .b(new_n331), .c(\a[30] ), .d(\b[29] ), .o1(new_n347));
  aoi112aa1n02x5               g252(.a(new_n347), .b(new_n346), .c(new_n342), .d(new_n343), .o1(new_n348));
  aoi022aa1n03x5               g253(.a(new_n345), .b(new_n346), .c(new_n340), .d(new_n348), .o1(\s[31] ));
  aoi022aa1n02x5               g254(.a(new_n100), .b(new_n99), .c(\a[1] ), .d(\b[0] ), .o1(new_n350));
  oaib12aa1n02x5               g255(.a(new_n350), .b(new_n100), .c(\a[2] ), .out0(new_n351));
  aboi22aa1n03x5               g256(.a(new_n105), .b(new_n106), .c(new_n99), .d(new_n100), .out0(new_n352));
  aoi022aa1n02x5               g257(.a(new_n351), .b(new_n352), .c(new_n146), .d(new_n148), .o1(\s[3] ));
  inv000aa1d42x5               g258(.a(new_n105), .o1(new_n354));
  nanp02aa1n02x5               g259(.a(new_n146), .b(new_n148), .o1(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n147), .b(new_n355), .c(new_n354), .out0(\s[4] ));
  inv000aa1d42x5               g261(.a(new_n115), .o1(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n357), .b(new_n149), .c(new_n108), .out0(\s[5] ));
  aoai13aa1n02x5               g263(.a(new_n116), .b(new_n123), .c(new_n109), .d(new_n357), .o1(new_n359));
  and002aa1n02x5               g264(.a(\b[5] ), .b(\a[6] ), .o(new_n360));
  norp03aa1n02x5               g265(.a(new_n360), .b(new_n124), .c(new_n123), .o1(new_n361));
  aoai13aa1n06x5               g266(.a(new_n361), .b(new_n115), .c(new_n149), .d(new_n108), .o1(new_n362));
  nanp02aa1n02x5               g267(.a(new_n359), .b(new_n362), .o1(\s[6] ));
  aboi22aa1n03x5               g268(.a(new_n360), .b(new_n362), .c(new_n118), .d(new_n111), .out0(new_n364));
  nanp03aa1n02x5               g269(.a(new_n362), .b(new_n118), .c(new_n125), .o1(new_n365));
  norb02aa1n02x5               g270(.a(new_n365), .b(new_n364), .out0(\s[7] ));
  norb02aa1n02x5               g271(.a(new_n112), .b(new_n113), .out0(new_n367));
  xnbna2aa1n03x5               g272(.a(new_n367), .b(new_n365), .c(new_n118), .out0(\s[8] ));
  aoi112aa1n02x5               g273(.a(new_n128), .b(new_n113), .c(new_n152), .d(new_n112), .o1(new_n369));
  aoi022aa1n02x5               g274(.a(new_n154), .b(new_n128), .c(new_n167), .d(new_n369), .o1(\s[9] ));
endmodule


