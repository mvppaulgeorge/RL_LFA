// Benchmark "adder" written by ABC on Thu Jul 18 05:28:58 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n332, new_n333, new_n336, new_n338, new_n339, new_n340,
    new_n342, new_n343, new_n344, new_n346, new_n348, new_n349, new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nand42aa1n03x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  orn002aa1n03x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nand42aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aob012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  nor002aa1n03x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n09x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor002aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n06x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nanp03aa1d12x5               g013(.a(new_n102), .b(new_n105), .c(new_n108), .o1(new_n109));
  tech160nm_fiaoi012aa1n05x5   g014(.a(new_n103), .b(new_n106), .c(new_n104), .o1(new_n110));
  nor042aa1n03x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanp02aa1n24x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n10x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nano23aa1n09x5               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  nor022aa1n04x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand02aa1n06x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor002aa1d32x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nand02aa1n04x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nand02aa1n04x5               g025(.a(new_n120), .b(new_n115), .o1(new_n121));
  inv040aa1n09x5               g026(.a(new_n118), .o1(new_n122));
  oaoi03aa1n06x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n113), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  aoi012aa1n06x5               g030(.a(new_n125), .b(new_n115), .c(new_n123), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n126), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n127));
  xorc02aa1n02x5               g032(.a(\a[10] ), .b(\b[9] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n97), .c(new_n127), .d(new_n98), .o1(new_n129));
  aoi112aa1n02x5               g034(.a(new_n128), .b(new_n97), .c(new_n127), .d(new_n98), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(\s[10] ));
  inv000aa1n03x5               g036(.a(new_n97), .o1(new_n132));
  tech160nm_fioaoi03aa1n03p5x5 g037(.a(\a[10] ), .b(\b[9] ), .c(new_n132), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  xorc02aa1n12x5               g039(.a(\a[11] ), .b(\b[10] ), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n129), .c(new_n134), .out0(\s[11] ));
  nor042aa1n06x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  aob012aa1n02x5               g043(.a(new_n135), .b(new_n129), .c(new_n134), .out0(new_n139));
  nor022aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  and002aa1n12x5               g045(.a(\b[11] ), .b(\a[12] ), .o(new_n141));
  nor002aa1n02x5               g046(.a(new_n141), .b(new_n140), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n135), .o1(new_n143));
  norp03aa1n02x5               g048(.a(new_n141), .b(new_n140), .c(new_n137), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n143), .c(new_n129), .d(new_n134), .o1(new_n145));
  aoai13aa1n03x5               g050(.a(new_n145), .b(new_n142), .c(new_n139), .d(new_n138), .o1(\s[12] ));
  nand42aa1n04x5               g051(.a(\b[9] ), .b(\a[10] ), .o1(new_n147));
  oai022aa1n04x5               g052(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n148));
  nano22aa1n02x4               g053(.a(new_n148), .b(new_n98), .c(new_n147), .out0(new_n149));
  nano22aa1n02x4               g054(.a(new_n143), .b(new_n149), .c(new_n142), .out0(new_n150));
  aoi012aa1n02x5               g055(.a(new_n140), .b(\a[11] ), .c(\b[10] ), .o1(new_n151));
  oai012aa1n02x5               g056(.a(new_n147), .b(\b[10] ), .c(\a[11] ), .o1(new_n152));
  nona23aa1n03x5               g057(.a(new_n151), .b(new_n148), .c(new_n152), .d(new_n141), .out0(new_n153));
  oabi12aa1n02x5               g058(.a(new_n141), .b(new_n137), .c(new_n140), .out0(new_n154));
  nanp02aa1n02x5               g059(.a(new_n153), .b(new_n154), .o1(new_n155));
  nor042aa1n04x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n157), .b(new_n156), .out0(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n155), .c(new_n127), .d(new_n150), .o1(new_n159));
  nano22aa1n02x4               g064(.a(new_n158), .b(new_n153), .c(new_n154), .out0(new_n160));
  aobi12aa1n02x5               g065(.a(new_n160), .b(new_n127), .c(new_n150), .out0(new_n161));
  norb02aa1n02x5               g066(.a(new_n159), .b(new_n161), .out0(\s[13] ));
  nor002aa1n04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand22aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  aoib12aa1n02x5               g069(.a(new_n156), .b(new_n164), .c(new_n163), .out0(new_n165));
  nano23aa1n06x5               g070(.a(new_n156), .b(new_n163), .c(new_n164), .d(new_n157), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n155), .c(new_n127), .d(new_n150), .o1(new_n167));
  aoi012aa1n12x5               g072(.a(new_n163), .b(new_n156), .c(new_n164), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n163), .b(new_n167), .c(new_n168), .o1(new_n169));
  aoi012aa1n02x5               g074(.a(new_n169), .b(new_n159), .c(new_n165), .o1(\s[14] ));
  nor042aa1n09x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n167), .c(new_n168), .out0(\s[15] ));
  inv000aa1d42x5               g079(.a(new_n171), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n173), .o1(new_n176));
  aoai13aa1n02x7               g081(.a(new_n175), .b(new_n176), .c(new_n167), .d(new_n168), .o1(new_n177));
  nor042aa1n02x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanp02aa1n04x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  norb03aa1n02x5               g085(.a(new_n179), .b(new_n171), .c(new_n178), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n176), .c(new_n167), .d(new_n168), .o1(new_n182));
  aob012aa1n03x5               g087(.a(new_n182), .b(new_n177), .c(new_n180), .out0(\s[16] ));
  nano23aa1n06x5               g088(.a(new_n171), .b(new_n178), .c(new_n179), .d(new_n172), .out0(new_n184));
  nand02aa1d04x5               g089(.a(new_n184), .b(new_n166), .o1(new_n185));
  nano32aa1n03x7               g090(.a(new_n185), .b(new_n149), .c(new_n142), .d(new_n135), .out0(new_n186));
  nanp02aa1n09x5               g091(.a(new_n127), .b(new_n186), .o1(new_n187));
  inv040aa1n03x5               g092(.a(new_n168), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n179), .b(new_n178), .c(new_n171), .o1(new_n189));
  aobi12aa1n06x5               g094(.a(new_n189), .b(new_n184), .c(new_n188), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n185), .c(new_n153), .d(new_n154), .o1(new_n191));
  inv000aa1n09x5               g096(.a(new_n191), .o1(new_n192));
  nanp02aa1n09x5               g097(.a(new_n187), .b(new_n192), .o1(new_n193));
  nor042aa1n03x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  nand42aa1n03x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aob012aa1n02x5               g101(.a(new_n184), .b(new_n167), .c(new_n168), .out0(new_n197));
  oaoi13aa1n02x5               g102(.a(new_n196), .b(new_n179), .c(new_n171), .d(new_n178), .o1(new_n198));
  aoi022aa1n02x5               g103(.a(new_n197), .b(new_n198), .c(new_n196), .d(new_n193), .o1(\s[17] ));
  nor042aa1n04x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nand42aa1n06x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  obai22aa1n02x7               g106(.a(new_n201), .b(new_n200), .c(\a[17] ), .d(\b[16] ), .out0(new_n202));
  aoi012aa1n02x5               g107(.a(new_n202), .b(new_n193), .c(new_n196), .o1(new_n203));
  nano23aa1n09x5               g108(.a(new_n194), .b(new_n200), .c(new_n201), .d(new_n195), .out0(new_n204));
  aoai13aa1n02x5               g109(.a(new_n204), .b(new_n191), .c(new_n127), .d(new_n186), .o1(new_n205));
  aoi012aa1n06x5               g110(.a(new_n200), .b(new_n194), .c(new_n201), .o1(new_n206));
  aoi012aa1n02x5               g111(.a(new_n200), .b(new_n205), .c(new_n206), .o1(new_n207));
  norp02aa1n02x5               g112(.a(new_n207), .b(new_n203), .o1(\s[18] ));
  nor002aa1d32x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand02aa1n03x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  norb02aa1n06x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n205), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g118(.a(new_n209), .o1(new_n214));
  inv040aa1n03x5               g119(.a(new_n206), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n211), .b(new_n215), .c(new_n193), .d(new_n204), .o1(new_n216));
  nor042aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand42aa1n02x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n06x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  norb03aa1n02x5               g124(.a(new_n218), .b(new_n209), .c(new_n217), .out0(new_n220));
  nanp02aa1n02x5               g125(.a(new_n216), .b(new_n220), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n219), .c(new_n214), .d(new_n216), .o1(\s[20] ));
  nano23aa1n06x5               g127(.a(new_n209), .b(new_n217), .c(new_n218), .d(new_n210), .out0(new_n223));
  and002aa1n02x5               g128(.a(new_n223), .b(new_n204), .o(new_n224));
  aoi112aa1n03x5               g129(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n225));
  oai112aa1n06x5               g130(.a(new_n211), .b(new_n219), .c(new_n225), .d(new_n200), .o1(new_n226));
  tech160nm_fioaoi03aa1n03p5x5 g131(.a(\a[20] ), .b(\b[19] ), .c(new_n214), .o1(new_n227));
  inv040aa1n02x5               g132(.a(new_n227), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(new_n226), .b(new_n228), .o1(new_n229));
  xorc02aa1n02x5               g134(.a(\a[21] ), .b(\b[20] ), .out0(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n229), .c(new_n193), .d(new_n224), .o1(new_n231));
  nona22aa1n02x4               g136(.a(new_n226), .b(new_n227), .c(new_n230), .out0(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n193), .c(new_n224), .o1(new_n233));
  norb02aa1n03x4               g138(.a(new_n231), .b(new_n233), .out0(\s[21] ));
  norp02aa1n02x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  xorc02aa1n02x5               g141(.a(\a[22] ), .b(\b[21] ), .out0(new_n237));
  oai022aa1n02x7               g142(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(\a[22] ), .c(\b[21] ), .o1(new_n239));
  nanp02aa1n03x5               g144(.a(new_n231), .b(new_n239), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n237), .c(new_n236), .d(new_n231), .o1(\s[22] ));
  nand22aa1n03x5               g146(.a(new_n237), .b(new_n230), .o1(new_n242));
  nano22aa1n02x4               g147(.a(new_n242), .b(new_n204), .c(new_n223), .out0(new_n243));
  inv000aa1d42x5               g148(.a(\a[22] ), .o1(new_n244));
  oaib12aa1n18x5               g149(.a(new_n238), .b(new_n244), .c(\b[21] ), .out0(new_n245));
  aoai13aa1n12x5               g150(.a(new_n245), .b(new_n242), .c(new_n226), .d(new_n228), .o1(new_n246));
  xorc02aa1n02x5               g151(.a(\a[23] ), .b(\b[22] ), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n246), .c(new_n193), .d(new_n243), .o1(new_n248));
  inv000aa1d42x5               g153(.a(\a[21] ), .o1(new_n249));
  xroi22aa1d04x5               g154(.a(new_n249), .b(\b[20] ), .c(new_n244), .d(\b[21] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n227), .c(new_n223), .d(new_n215), .o1(new_n251));
  nano22aa1n02x4               g156(.a(new_n247), .b(new_n251), .c(new_n245), .out0(new_n252));
  aobi12aa1n02x5               g157(.a(new_n252), .b(new_n193), .c(new_n243), .out0(new_n253));
  norb02aa1n02x5               g158(.a(new_n248), .b(new_n253), .out0(\s[23] ));
  nor042aa1d18x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  inv000aa1n09x5               g160(.a(new_n255), .o1(new_n256));
  xorc02aa1n02x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  oai022aa1n02x5               g162(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(\a[24] ), .c(\b[23] ), .o1(new_n259));
  nanp02aa1n03x5               g164(.a(new_n248), .b(new_n259), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n257), .c(new_n256), .d(new_n248), .o1(\s[24] ));
  nanp02aa1n02x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[23] ), .b(\a[24] ), .out0(new_n263));
  nano22aa1n12x5               g168(.a(new_n263), .b(new_n256), .c(new_n262), .out0(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  nano23aa1n02x4               g170(.a(new_n265), .b(new_n242), .c(new_n223), .d(new_n204), .out0(new_n266));
  tech160nm_fioaoi03aa1n03p5x5 g171(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n265), .c(new_n251), .d(new_n245), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n193), .d(new_n266), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(new_n270), .b(new_n267), .c(new_n246), .d(new_n264), .o1(new_n272));
  aobi12aa1n02x5               g177(.a(new_n272), .b(new_n193), .c(new_n266), .out0(new_n273));
  norb02aa1n03x4               g178(.a(new_n271), .b(new_n273), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  tech160nm_fixorc02aa1n03p5x5 g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  oai022aa1n02x5               g182(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n278));
  aoi012aa1n02x5               g183(.a(new_n278), .b(\a[26] ), .c(\b[25] ), .o1(new_n279));
  nand02aa1d04x5               g184(.a(new_n271), .b(new_n279), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n277), .c(new_n276), .d(new_n271), .o1(\s[26] ));
  nanp02aa1n02x5               g186(.a(new_n250), .b(new_n264), .o1(new_n282));
  and002aa1n02x5               g187(.a(new_n277), .b(new_n270), .o(new_n283));
  nano32aa1n03x7               g188(.a(new_n282), .b(new_n283), .c(new_n204), .d(new_n223), .out0(new_n284));
  aoai13aa1n09x5               g189(.a(new_n284), .b(new_n191), .c(new_n127), .d(new_n186), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n283), .b(new_n267), .c(new_n246), .d(new_n264), .o1(new_n286));
  aob012aa1n02x5               g191(.a(new_n278), .b(\b[25] ), .c(\a[26] ), .out0(new_n287));
  nand23aa1n06x5               g192(.a(new_n285), .b(new_n286), .c(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  and003aa1n02x5               g195(.a(new_n286), .b(new_n290), .c(new_n287), .o(new_n291));
  aoi022aa1n02x5               g196(.a(new_n291), .b(new_n285), .c(new_n288), .d(new_n289), .o1(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  nanp02aa1n03x5               g199(.a(new_n288), .b(new_n289), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .out0(new_n296));
  aobi12aa1n03x5               g201(.a(new_n287), .b(new_n269), .c(new_n283), .out0(new_n297));
  oai022aa1n02x5               g202(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n298));
  aoi012aa1n02x5               g203(.a(new_n298), .b(\a[28] ), .c(\b[27] ), .o1(new_n299));
  aoai13aa1n02x5               g204(.a(new_n299), .b(new_n290), .c(new_n297), .d(new_n285), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n294), .o1(\s[28] ));
  and002aa1n02x5               g206(.a(new_n296), .b(new_n289), .o(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  oaoi03aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n294), .o1(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[28] ), .b(\a[29] ), .out0(new_n305));
  norp02aa1n02x5               g210(.a(new_n304), .b(new_n305), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n306), .b(new_n303), .c(new_n297), .d(new_n285), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n305), .b(new_n304), .c(new_n288), .d(new_n302), .o1(new_n308));
  nanp02aa1n03x5               g213(.a(new_n308), .b(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g215(.a(new_n305), .b(new_n289), .c(new_n296), .out0(new_n311));
  nanp02aa1n03x5               g216(.a(new_n288), .b(new_n311), .o1(new_n312));
  norp02aa1n02x5               g217(.a(\b[28] ), .b(\a[29] ), .o1(new_n313));
  aoi022aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n314));
  aoi012aa1n02x5               g219(.a(new_n313), .b(new_n298), .c(new_n314), .o1(new_n315));
  norp02aa1n02x5               g220(.a(\b[29] ), .b(\a[30] ), .o1(new_n316));
  nanp02aa1n02x5               g221(.a(\b[29] ), .b(\a[30] ), .o1(new_n317));
  norb02aa1n02x5               g222(.a(new_n317), .b(new_n316), .out0(new_n318));
  inv000aa1n02x5               g223(.a(new_n311), .o1(new_n319));
  nona22aa1n02x4               g224(.a(new_n317), .b(new_n316), .c(new_n313), .out0(new_n320));
  aoi012aa1n02x5               g225(.a(new_n320), .b(new_n298), .c(new_n314), .o1(new_n321));
  aoai13aa1n02x5               g226(.a(new_n321), .b(new_n319), .c(new_n297), .d(new_n285), .o1(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n318), .c(new_n312), .d(new_n315), .o1(\s[30] ));
  nano32aa1n09x5               g228(.a(new_n305), .b(new_n296), .c(new_n289), .d(new_n318), .out0(new_n324));
  inv000aa1d42x5               g229(.a(new_n324), .o1(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[30] ), .b(\a[31] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n317), .b(new_n321), .out0(new_n327));
  norp02aa1n02x5               g232(.a(new_n327), .b(new_n326), .o1(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n325), .c(new_n297), .d(new_n285), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n326), .b(new_n327), .c(new_n288), .d(new_n324), .o1(new_n330));
  nanp02aa1n03x5               g235(.a(new_n330), .b(new_n329), .o1(\s[31] ));
  and003aa1n02x5               g236(.a(new_n99), .b(new_n101), .c(new_n100), .o(new_n332));
  nona23aa1n02x4               g237(.a(new_n107), .b(new_n99), .c(new_n332), .d(new_n106), .out0(new_n333));
  oaib12aa1n02x5               g238(.a(new_n333), .b(new_n108), .c(new_n102), .out0(\s[3] ));
  xobna2aa1n03x5               g239(.a(new_n105), .b(new_n333), .c(new_n107), .out0(\s[4] ));
  norb02aa1n02x5               g240(.a(new_n119), .b(new_n118), .out0(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n336), .b(new_n109), .c(new_n110), .out0(\s[5] ));
  norb02aa1n02x5               g242(.a(new_n117), .b(new_n116), .out0(new_n338));
  nanp02aa1n02x5               g243(.a(new_n109), .b(new_n110), .o1(new_n339));
  nanp02aa1n02x5               g244(.a(new_n339), .b(new_n336), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n338), .b(new_n340), .c(new_n122), .out0(\s[6] ));
  norb02aa1n02x5               g246(.a(new_n114), .b(new_n113), .out0(new_n342));
  aoai13aa1n02x5               g247(.a(new_n342), .b(new_n123), .c(new_n339), .d(new_n120), .o1(new_n343));
  aoi112aa1n02x5               g248(.a(new_n342), .b(new_n123), .c(new_n339), .d(new_n120), .o1(new_n344));
  norb02aa1n02x5               g249(.a(new_n343), .b(new_n344), .out0(\s[7] ));
  norb02aa1n02x5               g250(.a(new_n112), .b(new_n111), .out0(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n343), .c(new_n124), .out0(\s[8] ));
  nanb02aa1n02x5               g252(.a(new_n97), .b(new_n98), .out0(new_n348));
  aoi112aa1n02x5               g253(.a(new_n348), .b(new_n125), .c(new_n115), .d(new_n123), .o1(new_n349));
  aoai13aa1n02x5               g254(.a(new_n349), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n350));
  aob012aa1n02x5               g255(.a(new_n350), .b(new_n127), .c(new_n348), .out0(\s[9] ));
endmodule


