// Benchmark "adder" written by ABC on Thu Jul 18 05:38:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n349, new_n351, new_n353, new_n355,
    new_n357, new_n358;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n12x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nand02aa1d28x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  nanb02aa1n02x5               g004(.a(new_n98), .b(new_n99), .out0(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[1] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand22aa1n12x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  aob012aa1n06x5               g010(.a(new_n103), .b(new_n104), .c(new_n105), .out0(new_n106));
  nor002aa1d24x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nand22aa1n12x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nor022aa1n16x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nand42aa1n04x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  norb02aa1n02x5               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  nand23aa1n04x5               g017(.a(new_n106), .b(new_n109), .c(new_n112), .o1(new_n113));
  aoi012aa1n06x5               g018(.a(new_n107), .b(new_n110), .c(new_n108), .o1(new_n114));
  nor022aa1n16x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand42aa1n16x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor002aa1d32x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nanp02aa1n04x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nano23aa1n02x5               g023(.a(new_n115), .b(new_n117), .c(new_n118), .d(new_n116), .out0(new_n119));
  nor042aa1d18x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nand22aa1n09x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nanb02aa1n03x5               g026(.a(new_n120), .b(new_n121), .out0(new_n122));
  nor042aa1d18x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nand02aa1d28x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nanb02aa1n12x5               g029(.a(new_n123), .b(new_n124), .out0(new_n125));
  nona22aa1n03x5               g030(.a(new_n119), .b(new_n122), .c(new_n125), .out0(new_n126));
  norb02aa1n15x5               g031(.a(new_n121), .b(new_n120), .out0(new_n127));
  nano22aa1n12x5               g032(.a(new_n123), .b(new_n116), .c(new_n124), .out0(new_n128));
  oai022aa1d18x5               g033(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n129));
  oa0012aa1n03x5               g034(.a(new_n121), .b(new_n123), .c(new_n120), .o(new_n130));
  aoi013aa1n06x4               g035(.a(new_n130), .b(new_n128), .c(new_n129), .d(new_n127), .o1(new_n131));
  aoai13aa1n12x5               g036(.a(new_n131), .b(new_n126), .c(new_n113), .d(new_n114), .o1(new_n132));
  oabi12aa1n02x5               g037(.a(new_n132), .b(\a[9] ), .c(\b[8] ), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n100), .b(new_n133), .c(new_n97), .out0(\s[10] ));
  nano22aa1n02x4               g039(.a(new_n98), .b(new_n97), .c(new_n99), .out0(new_n135));
  nor042aa1d18x5               g040(.a(\b[8] ), .b(\a[9] ), .o1(new_n136));
  tech160nm_fioai012aa1n05x5   g041(.a(new_n135), .b(new_n132), .c(new_n136), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n98), .b(new_n136), .c(new_n99), .o1(new_n138));
  nor042aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1d28x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n137), .c(new_n138), .out0(\s[11] ));
  aob012aa1n03x5               g047(.a(new_n141), .b(new_n137), .c(new_n138), .out0(new_n143));
  inv000aa1d42x5               g048(.a(\a[11] ), .o1(new_n144));
  oaib12aa1n03x5               g049(.a(new_n143), .b(\b[10] ), .c(new_n144), .out0(new_n145));
  nor042aa1n09x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1d28x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  aoib12aa1n02x5               g053(.a(new_n139), .b(new_n147), .c(new_n146), .out0(new_n149));
  aoi022aa1n02x5               g054(.a(new_n145), .b(new_n148), .c(new_n143), .d(new_n149), .o1(\s[12] ));
  nano23aa1n09x5               g055(.a(new_n139), .b(new_n146), .c(new_n147), .d(new_n140), .out0(new_n151));
  nano23aa1n09x5               g056(.a(new_n136), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n152));
  nand22aa1n09x5               g057(.a(new_n152), .b(new_n151), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n03x5               g059(.a(new_n140), .b(new_n98), .c(new_n136), .d(new_n99), .o1(new_n155));
  nona22aa1n03x5               g060(.a(new_n155), .b(new_n146), .c(new_n139), .out0(new_n156));
  and002aa1n02x5               g061(.a(new_n156), .b(new_n147), .o(new_n157));
  nor042aa1n09x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand02aa1n16x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n159), .b(new_n158), .out0(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n157), .c(new_n132), .d(new_n154), .o1(new_n161));
  aoi112aa1n02x5               g066(.a(new_n160), .b(new_n157), .c(new_n132), .d(new_n154), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n161), .b(new_n162), .out0(\s[13] ));
  nor002aa1d32x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  inv000aa1d42x5               g069(.a(\a[13] ), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[12] ), .o1(new_n166));
  nand42aa1d28x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  aboi22aa1n03x5               g072(.a(new_n164), .b(new_n167), .c(new_n165), .d(new_n166), .out0(new_n168));
  nano23aa1d15x5               g073(.a(new_n158), .b(new_n164), .c(new_n167), .d(new_n159), .out0(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n157), .c(new_n132), .d(new_n154), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n167), .b(new_n164), .c(new_n165), .d(new_n166), .o1(new_n171));
  nand22aa1n03x5               g076(.a(new_n170), .b(new_n171), .o1(new_n172));
  aboi22aa1n03x5               g077(.a(new_n164), .b(new_n172), .c(new_n161), .d(new_n168), .out0(\s[14] ));
  nor022aa1n08x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nand02aa1d20x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n170), .c(new_n171), .out0(\s[15] ));
  aoi012aa1n03x5               g082(.a(new_n174), .b(new_n172), .c(new_n175), .o1(new_n178));
  nor042aa1n09x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand02aa1d28x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n176), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n180), .o1(new_n183));
  oai022aa1d24x5               g088(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n184));
  norp02aa1n02x5               g089(.a(new_n184), .b(new_n183), .o1(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n182), .c(new_n170), .d(new_n171), .o1(new_n186));
  tech160nm_fioai012aa1n02p5x5 g091(.a(new_n186), .b(new_n178), .c(new_n181), .o1(\s[16] ));
  tech160nm_fioaoi03aa1n02p5x5 g092(.a(new_n101), .b(new_n102), .c(new_n105), .o1(new_n188));
  nona23aa1n03x5               g093(.a(new_n111), .b(new_n108), .c(new_n107), .d(new_n110), .out0(new_n189));
  oaih12aa1n06x5               g094(.a(new_n114), .b(new_n189), .c(new_n188), .o1(new_n190));
  nona23aa1n02x4               g095(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n191));
  nor043aa1n03x5               g096(.a(new_n191), .b(new_n122), .c(new_n125), .o1(new_n192));
  nand43aa1n02x5               g097(.a(new_n128), .b(new_n127), .c(new_n129), .o1(new_n193));
  norb03aa1n03x5               g098(.a(new_n121), .b(new_n120), .c(new_n123), .out0(new_n194));
  oaib12aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n121), .out0(new_n195));
  nano23aa1n06x5               g100(.a(new_n174), .b(new_n179), .c(new_n180), .d(new_n175), .out0(new_n196));
  nano22aa1d15x5               g101(.a(new_n153), .b(new_n169), .c(new_n196), .out0(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n195), .c(new_n190), .d(new_n192), .o1(new_n198));
  nano22aa1n12x5               g103(.a(new_n179), .b(new_n175), .c(new_n180), .out0(new_n199));
  oai012aa1n02x5               g104(.a(new_n147), .b(\b[12] ), .c(\a[13] ), .o1(new_n200));
  oai012aa1n02x5               g105(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .o1(new_n201));
  oai012aa1n06x5               g106(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .o1(new_n202));
  norp03aa1n06x5               g107(.a(new_n202), .b(new_n201), .c(new_n200), .o1(new_n203));
  oab012aa1n06x5               g108(.a(new_n202), .b(new_n158), .c(new_n164), .out0(new_n204));
  aoi022aa1n09x5               g109(.a(new_n204), .b(new_n199), .c(new_n180), .d(new_n184), .o1(new_n205));
  inv020aa1n03x5               g110(.a(new_n205), .o1(new_n206));
  aoi013aa1n09x5               g111(.a(new_n206), .b(new_n156), .c(new_n199), .d(new_n203), .o1(new_n207));
  nanp02aa1n09x5               g112(.a(new_n198), .b(new_n207), .o1(new_n208));
  nor002aa1d32x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(\b[16] ), .b(\a[17] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  nanp02aa1n03x5               g116(.a(new_n172), .b(new_n196), .o1(new_n212));
  aboi22aa1n03x5               g117(.a(new_n209), .b(new_n210), .c(new_n184), .d(new_n180), .out0(new_n213));
  aoi022aa1n02x7               g118(.a(new_n212), .b(new_n213), .c(new_n211), .d(new_n208), .o1(\s[17] ));
  nor042aa1d18x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  nanp02aa1n24x5               g120(.a(\b[17] ), .b(\a[18] ), .o1(new_n216));
  obai22aa1n02x7               g121(.a(new_n216), .b(new_n215), .c(\a[17] ), .d(\b[16] ), .out0(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(new_n208), .c(new_n211), .o1(new_n218));
  nand43aa1n02x5               g123(.a(new_n156), .b(new_n199), .c(new_n203), .o1(new_n219));
  nand02aa1n03x5               g124(.a(new_n219), .b(new_n205), .o1(new_n220));
  nano23aa1n09x5               g125(.a(new_n209), .b(new_n215), .c(new_n216), .d(new_n210), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n220), .c(new_n132), .d(new_n197), .o1(new_n222));
  nor002aa1n03x5               g127(.a(new_n215), .b(new_n209), .o1(new_n223));
  norb02aa1n06x4               g128(.a(new_n216), .b(new_n223), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  nanp02aa1n02x5               g130(.a(new_n222), .b(new_n225), .o1(new_n226));
  aoib12aa1n02x5               g131(.a(new_n218), .b(new_n226), .c(new_n215), .out0(\s[18] ));
  xorc02aa1n02x5               g132(.a(\a[19] ), .b(\b[18] ), .out0(new_n228));
  xnbna2aa1n03x5               g133(.a(new_n228), .b(new_n222), .c(new_n225), .out0(\s[19] ));
  xnrc02aa1n02x5               g134(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g135(.a(\b[18] ), .b(\a[19] ), .o1(new_n231));
  inv030aa1n02x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n228), .b(new_n224), .c(new_n208), .d(new_n221), .o1(new_n233));
  nor002aa1n20x5               g138(.a(\b[19] ), .b(\a[20] ), .o1(new_n234));
  nanp02aa1n12x5               g139(.a(\b[19] ), .b(\a[20] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n235), .b(new_n234), .out0(new_n236));
  and002aa1n02x5               g141(.a(\b[19] ), .b(\a[20] ), .o(new_n237));
  oai022aa1n02x5               g142(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n238));
  nona22aa1n02x5               g143(.a(new_n233), .b(new_n237), .c(new_n238), .out0(new_n239));
  aoai13aa1n03x5               g144(.a(new_n239), .b(new_n236), .c(new_n233), .d(new_n232), .o1(\s[20] ));
  nand42aa1n04x5               g145(.a(\b[18] ), .b(\a[19] ), .o1(new_n241));
  nano23aa1n09x5               g146(.a(new_n231), .b(new_n234), .c(new_n235), .d(new_n241), .out0(new_n242));
  tech160nm_finand02aa1n05x5   g147(.a(new_n242), .b(new_n221), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  nanb03aa1n03x5               g149(.a(new_n234), .b(new_n235), .c(new_n241), .out0(new_n245));
  oai112aa1n03x5               g150(.a(new_n232), .b(new_n216), .c(new_n215), .d(new_n209), .o1(new_n246));
  oaih12aa1n06x5               g151(.a(new_n235), .b(new_n234), .c(new_n231), .o1(new_n247));
  tech160nm_fioai012aa1n05x5   g152(.a(new_n247), .b(new_n246), .c(new_n245), .o1(new_n248));
  xorc02aa1n12x5               g153(.a(\a[21] ), .b(\b[20] ), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n248), .c(new_n208), .d(new_n244), .o1(new_n250));
  aoi112aa1n02x5               g155(.a(new_n249), .b(new_n248), .c(new_n208), .d(new_n244), .o1(new_n251));
  norb02aa1n03x4               g156(.a(new_n250), .b(new_n251), .out0(\s[21] ));
  inv000aa1d42x5               g157(.a(\a[21] ), .o1(new_n253));
  nanb02aa1n12x5               g158(.a(\b[20] ), .b(new_n253), .out0(new_n254));
  xorc02aa1n02x5               g159(.a(\a[22] ), .b(\b[21] ), .out0(new_n255));
  nanp02aa1n02x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  oai022aa1n02x5               g161(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n256), .b(new_n257), .out0(new_n258));
  tech160nm_finand02aa1n03p5x5 g163(.a(new_n250), .b(new_n258), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n255), .c(new_n250), .d(new_n254), .o1(\s[22] ));
  nanp02aa1n02x5               g165(.a(new_n255), .b(new_n249), .o1(new_n261));
  nano22aa1n02x4               g166(.a(new_n261), .b(new_n242), .c(new_n221), .out0(new_n262));
  nano22aa1n02x5               g167(.a(new_n234), .b(new_n241), .c(new_n235), .out0(new_n263));
  oai012aa1n02x5               g168(.a(new_n216), .b(\b[18] ), .c(\a[19] ), .o1(new_n264));
  nona22aa1n03x5               g169(.a(new_n263), .b(new_n223), .c(new_n264), .out0(new_n265));
  oaoi03aa1n12x5               g170(.a(\a[22] ), .b(\b[21] ), .c(new_n254), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n261), .c(new_n265), .d(new_n247), .o1(new_n268));
  nor042aa1n06x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(\b[22] ), .b(\a[23] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n270), .b(new_n269), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n268), .c(new_n208), .d(new_n262), .o1(new_n272));
  aoi112aa1n02x5               g177(.a(new_n271), .b(new_n268), .c(new_n208), .d(new_n262), .o1(new_n273));
  norb02aa1n03x4               g178(.a(new_n272), .b(new_n273), .out0(\s[23] ));
  inv040aa1n06x5               g179(.a(new_n269), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[24] ), .b(\b[23] ), .out0(new_n276));
  and002aa1n02x5               g181(.a(\b[23] ), .b(\a[24] ), .o(new_n277));
  oai022aa1n02x5               g182(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n278));
  nona22aa1n02x5               g183(.a(new_n272), .b(new_n277), .c(new_n278), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n272), .d(new_n275), .o1(\s[24] ));
  inv000aa1d42x5               g185(.a(\a[22] ), .o1(new_n281));
  xroi22aa1d04x5               g186(.a(new_n253), .b(\b[20] ), .c(new_n281), .d(\b[21] ), .out0(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[23] ), .b(\a[24] ), .out0(new_n283));
  nano22aa1n06x5               g188(.a(new_n283), .b(new_n275), .c(new_n270), .out0(new_n284));
  nano22aa1n03x7               g189(.a(new_n243), .b(new_n282), .c(new_n284), .out0(new_n285));
  aobi12aa1n06x5               g190(.a(new_n285), .b(new_n198), .c(new_n207), .out0(new_n286));
  inv000aa1n03x5               g191(.a(new_n286), .o1(new_n287));
  tech160nm_fioaoi03aa1n03p5x5 g192(.a(\a[24] ), .b(\b[23] ), .c(new_n275), .o1(new_n288));
  tech160nm_fiaoi012aa1n02p5x5 g193(.a(new_n288), .b(new_n268), .c(new_n284), .o1(new_n289));
  xnrc02aa1n12x5               g194(.a(\b[24] ), .b(\a[25] ), .out0(new_n290));
  xobna2aa1n03x5               g195(.a(new_n290), .b(new_n287), .c(new_n289), .out0(\s[25] ));
  norp02aa1n02x5               g196(.a(\b[24] ), .b(\a[25] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  inv020aa1n02x5               g198(.a(new_n289), .o1(new_n294));
  oabi12aa1n03x5               g199(.a(new_n290), .b(new_n286), .c(new_n294), .out0(new_n295));
  xorc02aa1n06x5               g200(.a(\a[26] ), .b(\b[25] ), .out0(new_n296));
  nanp02aa1n02x5               g201(.a(\b[25] ), .b(\a[26] ), .o1(new_n297));
  oai022aa1n02x5               g202(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n298));
  norb02aa1n02x5               g203(.a(new_n297), .b(new_n298), .out0(new_n299));
  nand42aa1n02x5               g204(.a(new_n295), .b(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n293), .o1(\s[26] ));
  norb02aa1n02x5               g206(.a(new_n296), .b(new_n290), .out0(new_n302));
  nano32aa1n03x7               g207(.a(new_n243), .b(new_n302), .c(new_n282), .d(new_n284), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n220), .c(new_n132), .d(new_n197), .o1(new_n304));
  aoai13aa1n02x5               g209(.a(new_n302), .b(new_n288), .c(new_n268), .d(new_n284), .o1(new_n305));
  nanp02aa1n02x5               g210(.a(new_n298), .b(new_n297), .o1(new_n306));
  nanp03aa1n03x5               g211(.a(new_n304), .b(new_n305), .c(new_n306), .o1(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g213(.a(\b[26] ), .b(\a[27] ), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  aobi12aa1n09x5               g215(.a(new_n303), .b(new_n198), .c(new_n207), .out0(new_n311));
  aoai13aa1n02x7               g216(.a(new_n284), .b(new_n266), .c(new_n248), .d(new_n282), .o1(new_n312));
  inv000aa1n02x5               g217(.a(new_n288), .o1(new_n313));
  inv000aa1n02x5               g218(.a(new_n302), .o1(new_n314));
  aoai13aa1n09x5               g219(.a(new_n306), .b(new_n314), .c(new_n312), .d(new_n313), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[27] ), .b(\b[26] ), .out0(new_n316));
  oaih12aa1n02x5               g221(.a(new_n316), .b(new_n315), .c(new_n311), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[28] ), .b(\b[27] ), .out0(new_n318));
  oai022aa1d24x5               g223(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n319), .b(\a[28] ), .c(\b[27] ), .o1(new_n320));
  tech160nm_finand02aa1n03p5x5 g225(.a(new_n317), .b(new_n320), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n318), .c(new_n317), .d(new_n310), .o1(\s[28] ));
  xorc02aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(new_n318), .b(new_n316), .o(new_n324));
  oaih12aa1n02x5               g229(.a(new_n324), .b(new_n315), .c(new_n311), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[27] ), .o1(new_n326));
  oaib12aa1n09x5               g231(.a(new_n319), .b(new_n326), .c(\a[28] ), .out0(new_n327));
  nanp03aa1n03x5               g232(.a(new_n325), .b(new_n327), .c(new_n323), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n327), .o1(new_n329));
  oaoi13aa1n03x5               g234(.a(new_n329), .b(new_n324), .c(new_n315), .d(new_n311), .o1(new_n330));
  oaih12aa1n02x5               g235(.a(new_n328), .b(new_n330), .c(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g236(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g237(.a(new_n316), .b(new_n323), .c(new_n318), .o(new_n333));
  tech160nm_fioaoi03aa1n03p5x5 g238(.a(\a[29] ), .b(\b[28] ), .c(new_n327), .o1(new_n334));
  oaoi13aa1n03x5               g239(.a(new_n334), .b(new_n333), .c(new_n315), .d(new_n311), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[30] ), .b(\b[29] ), .out0(new_n336));
  oaih12aa1n02x5               g241(.a(new_n333), .b(new_n315), .c(new_n311), .o1(new_n337));
  norb02aa1n03x5               g242(.a(new_n336), .b(new_n334), .out0(new_n338));
  nand42aa1n04x5               g243(.a(new_n337), .b(new_n338), .o1(new_n339));
  oaih12aa1n02x5               g244(.a(new_n339), .b(new_n335), .c(new_n336), .o1(\s[30] ));
  xnrc02aa1n02x5               g245(.a(\b[30] ), .b(\a[31] ), .out0(new_n341));
  and003aa1n02x5               g246(.a(new_n324), .b(new_n336), .c(new_n323), .o(new_n342));
  tech160nm_fiaoi012aa1n03p5x5 g247(.a(new_n338), .b(\a[30] ), .c(\b[29] ), .o1(new_n343));
  aoai13aa1n03x5               g248(.a(new_n341), .b(new_n343), .c(new_n307), .d(new_n342), .o1(new_n344));
  oaih12aa1n02x5               g249(.a(new_n342), .b(new_n315), .c(new_n311), .o1(new_n345));
  nona22aa1n03x5               g250(.a(new_n345), .b(new_n343), .c(new_n341), .out0(new_n346));
  nanp02aa1n03x5               g251(.a(new_n344), .b(new_n346), .o1(\s[31] ));
  xorb03aa1n02x5               g252(.a(new_n106), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi13aa1n02x5               g253(.a(new_n109), .b(new_n111), .c(new_n106), .d(new_n110), .o1(new_n349));
  aoib12aa1n02x5               g254(.a(new_n349), .b(new_n190), .c(new_n107), .out0(\s[4] ));
  norb02aa1n02x5               g255(.a(new_n118), .b(new_n117), .out0(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n351), .b(new_n113), .c(new_n114), .out0(\s[5] ));
  aoi012aa1n02x5               g257(.a(new_n117), .b(new_n190), .c(new_n118), .o1(new_n353));
  xnrb03aa1n02x5               g258(.a(new_n353), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g259(.a(\a[6] ), .b(\b[5] ), .c(new_n353), .o1(new_n355));
  xorb03aa1n02x5               g260(.a(new_n355), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g261(.a(new_n125), .b(new_n355), .out0(new_n357));
  aoai13aa1n02x5               g262(.a(new_n122), .b(new_n123), .c(new_n355), .d(new_n124), .o1(new_n358));
  aob012aa1n02x5               g263(.a(new_n358), .b(new_n357), .c(new_n194), .out0(\s[8] ));
  xorb03aa1n02x5               g264(.a(new_n132), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


