// Benchmark "adder" written by ABC on Thu Jul 11 11:56:47 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n304, new_n307, new_n309, new_n311;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  160nm_ficinv00aa1n08x5       g001(.clk(\a[9] ), .clkout(new_n97));
  160nm_ficinv00aa1n08x5       g002(.clk(\b[8] ), .clkout(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  and002aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  norp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oai012aa1n02x5               g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norp02aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nona23aa1n02x4               g013(.a(new_n108), .b(new_n106), .c(new_n105), .d(new_n107), .out0(new_n109));
  aoi012aa1n02x5               g014(.a(new_n105), .b(new_n107), .c(new_n106), .o1(new_n110));
  oai012aa1n02x5               g015(.a(new_n110), .b(new_n109), .c(new_n104), .o1(new_n111));
  xnrc02aa1n02x5               g016(.a(\b[5] ), .b(\a[6] ), .out0(new_n112));
  norp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  norp03aa1n02x5               g023(.a(new_n117), .b(new_n118), .c(new_n112), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n111), .b(new_n119), .o1(new_n120));
  oai022aa1n02x5               g025(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n121));
  160nm_ficinv00aa1n08x5       g026(.clk(\a[5] ), .clkout(new_n122));
  160nm_ficinv00aa1n08x5       g027(.clk(\b[4] ), .clkout(new_n123));
  nanp02aa1n02x5               g028(.a(new_n123), .b(new_n122), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[6] ), .b(\b[5] ), .c(new_n124), .o1(new_n125));
  aboi22aa1n03x5               g030(.a(new_n117), .b(new_n125), .c(new_n114), .d(new_n121), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n99), .b(new_n100), .c(new_n120), .d(new_n126), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  norp02aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  160nm_ficinv00aa1n08x5       g036(.clk(new_n131), .clkout(new_n132));
  norp02aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n136));
  160nm_ficinv00aa1n08x5       g041(.clk(new_n136), .clkout(new_n137));
  aoai13aa1n02x5               g042(.a(new_n135), .b(new_n137), .c(new_n127), .d(new_n132), .o1(new_n138));
  aoi112aa1n02x5               g043(.a(new_n135), .b(new_n137), .c(new_n127), .d(new_n132), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n138), .b(new_n139), .out0(\s[11] ));
  160nm_ficinv00aa1n08x5       g045(.clk(new_n133), .clkout(new_n141));
  norp02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n138), .c(new_n141), .out0(\s[12] ));
  xnrc02aa1n02x5               g050(.a(\b[8] ), .b(\a[9] ), .out0(new_n146));
  nano23aa1n02x4               g051(.a(new_n133), .b(new_n142), .c(new_n143), .d(new_n134), .out0(new_n147));
  nona22aa1n02x4               g052(.a(new_n147), .b(new_n146), .c(new_n131), .out0(new_n148));
  160nm_ficinv00aa1n08x5       g053(.clk(new_n142), .clkout(new_n149));
  nona23aa1n02x4               g054(.a(new_n143), .b(new_n134), .c(new_n133), .d(new_n142), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n133), .b(new_n143), .o1(new_n151));
  oai112aa1n02x5               g056(.a(new_n151), .b(new_n149), .c(new_n150), .d(new_n136), .o1(new_n152));
  160nm_ficinv00aa1n08x5       g057(.clk(new_n152), .clkout(new_n153));
  aoai13aa1n02x5               g058(.a(new_n153), .b(new_n148), .c(new_n120), .d(new_n126), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n156), .b(new_n154), .c(new_n157), .o1(new_n158));
  xnrb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n02x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  norp02aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1n02x4               g069(.a(new_n156), .b(new_n163), .c(new_n164), .d(new_n157), .out0(new_n165));
  oai012aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n156), .o1(new_n166));
  160nm_ficinv00aa1n08x5       g071(.clk(new_n166), .clkout(new_n167));
  aoai13aa1n02x5               g072(.a(new_n162), .b(new_n167), .c(new_n154), .d(new_n165), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n162), .b(new_n167), .c(new_n154), .d(new_n165), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(\s[15] ));
  160nm_ficinv00aa1n08x5       g075(.clk(new_n160), .clkout(new_n171));
  norp02aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n168), .c(new_n171), .out0(\s[16] ));
  oai012aa1n02x5               g080(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n176));
  oaib12aa1n02x5               g081(.a(new_n176), .b(new_n117), .c(new_n125), .out0(new_n177));
  nano32aa1n02x4               g082(.a(new_n148), .b(new_n174), .c(new_n162), .d(new_n165), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n177), .c(new_n111), .d(new_n119), .o1(new_n179));
  nona23aa1n02x4               g084(.a(new_n173), .b(new_n161), .c(new_n160), .d(new_n172), .out0(new_n180));
  norb02aa1n02x5               g085(.a(new_n165), .b(new_n180), .out0(new_n181));
  aoi112aa1n02x5               g086(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n182));
  oai022aa1n02x5               g087(.a(new_n180), .b(new_n166), .c(\b[15] ), .d(\a[16] ), .o1(new_n183));
  aoi112aa1n02x5               g088(.a(new_n183), .b(new_n182), .c(new_n152), .d(new_n181), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n184), .b(new_n179), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g091(.clk(\a[18] ), .clkout(new_n187));
  160nm_ficinv00aa1n08x5       g092(.clk(\a[17] ), .clkout(new_n188));
  160nm_ficinv00aa1n08x5       g093(.clk(\b[16] ), .clkout(new_n189));
  oaoi03aa1n02x5               g094(.a(new_n188), .b(new_n189), .c(new_n185), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(new_n187), .out0(\s[18] ));
  xroi22aa1d04x5               g096(.a(new_n188), .b(\b[16] ), .c(new_n187), .d(\b[17] ), .out0(new_n192));
  nanp02aa1n02x5               g097(.a(new_n189), .b(new_n188), .o1(new_n193));
  oaoi03aa1n02x5               g098(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n194));
  norp02aa1n02x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nanp02aa1n02x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  norb02aa1n02x5               g101(.a(new_n196), .b(new_n195), .out0(new_n197));
  aoai13aa1n02x5               g102(.a(new_n197), .b(new_n194), .c(new_n185), .d(new_n192), .o1(new_n198));
  aoi112aa1n02x5               g103(.a(new_n197), .b(new_n194), .c(new_n185), .d(new_n192), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  nona22aa1n02x4               g109(.a(new_n198), .b(new_n204), .c(new_n195), .out0(new_n205));
  orn002aa1n02x5               g110(.a(\a[19] ), .b(\b[18] ), .o(new_n206));
  aobi12aa1n02x5               g111(.a(new_n204), .b(new_n198), .c(new_n206), .out0(new_n207));
  norb02aa1n02x5               g112(.a(new_n205), .b(new_n207), .out0(\s[20] ));
  nano23aa1n02x4               g113(.a(new_n195), .b(new_n202), .c(new_n203), .d(new_n196), .out0(new_n209));
  nanp02aa1n02x5               g114(.a(new_n192), .b(new_n209), .o1(new_n210));
  oai022aa1n02x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  oaib12aa1n02x5               g116(.a(new_n211), .b(new_n187), .c(\b[17] ), .out0(new_n212));
  nona23aa1n02x4               g117(.a(new_n203), .b(new_n196), .c(new_n195), .d(new_n202), .out0(new_n213));
  oaoi03aa1n02x5               g118(.a(\a[20] ), .b(\b[19] ), .c(new_n206), .o1(new_n214));
  oabi12aa1n02x5               g119(.a(new_n214), .b(new_n213), .c(new_n212), .out0(new_n215));
  160nm_ficinv00aa1n08x5       g120(.clk(new_n215), .clkout(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n210), .c(new_n184), .d(new_n179), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[21] ), .b(\b[20] ), .out0(new_n220));
  xorc02aa1n02x5               g125(.a(\a[22] ), .b(\b[21] ), .out0(new_n221));
  aoi112aa1n02x5               g126(.a(new_n219), .b(new_n221), .c(new_n217), .d(new_n220), .o1(new_n222));
  aoai13aa1n02x5               g127(.a(new_n221), .b(new_n219), .c(new_n217), .d(new_n220), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(\s[22] ));
  160nm_ficinv00aa1n08x5       g129(.clk(\a[21] ), .clkout(new_n225));
  160nm_ficinv00aa1n08x5       g130(.clk(\a[22] ), .clkout(new_n226));
  xroi22aa1d04x5               g131(.a(new_n225), .b(\b[20] ), .c(new_n226), .d(\b[21] ), .out0(new_n227));
  nanp03aa1n02x5               g132(.a(new_n227), .b(new_n192), .c(new_n209), .o1(new_n228));
  160nm_ficinv00aa1n08x5       g133(.clk(\b[21] ), .clkout(new_n229));
  oaoi03aa1n02x5               g134(.a(new_n226), .b(new_n229), .c(new_n219), .o1(new_n230));
  160nm_ficinv00aa1n08x5       g135(.clk(new_n230), .clkout(new_n231));
  aoi012aa1n02x5               g136(.a(new_n231), .b(new_n215), .c(new_n227), .o1(new_n232));
  aoai13aa1n02x5               g137(.a(new_n232), .b(new_n228), .c(new_n184), .d(new_n179), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  xorc02aa1n02x5               g140(.a(\a[23] ), .b(\b[22] ), .out0(new_n236));
  xorc02aa1n02x5               g141(.a(\a[24] ), .b(\b[23] ), .out0(new_n237));
  aoi112aa1n02x5               g142(.a(new_n235), .b(new_n237), .c(new_n233), .d(new_n236), .o1(new_n238));
  aoai13aa1n02x5               g143(.a(new_n237), .b(new_n235), .c(new_n233), .d(new_n236), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n238), .out0(\s[24] ));
  and002aa1n02x5               g145(.a(new_n237), .b(new_n236), .o(new_n241));
  160nm_ficinv00aa1n08x5       g146(.clk(new_n241), .clkout(new_n242));
  nano32aa1n02x4               g147(.a(new_n242), .b(new_n227), .c(new_n192), .d(new_n209), .out0(new_n243));
  aoai13aa1n02x5               g148(.a(new_n227), .b(new_n214), .c(new_n209), .d(new_n194), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n245));
  oab012aa1n02x4               g150(.a(new_n245), .b(\a[24] ), .c(\b[23] ), .out0(new_n246));
  aoai13aa1n02x5               g151(.a(new_n246), .b(new_n242), .c(new_n244), .d(new_n230), .o1(new_n247));
  xorc02aa1n02x5               g152(.a(\a[25] ), .b(\b[24] ), .out0(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n247), .c(new_n185), .d(new_n243), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(new_n248), .b(new_n247), .c(new_n185), .d(new_n243), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n249), .b(new_n250), .out0(\s[25] ));
  norp02aa1n02x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[26] ), .b(\b[25] ), .out0(new_n253));
  nona22aa1n02x4               g158(.a(new_n249), .b(new_n253), .c(new_n252), .out0(new_n254));
  160nm_ficinv00aa1n08x5       g159(.clk(new_n252), .clkout(new_n255));
  aobi12aa1n02x5               g160(.a(new_n253), .b(new_n249), .c(new_n255), .out0(new_n256));
  norb02aa1n02x5               g161(.a(new_n254), .b(new_n256), .out0(\s[26] ));
  and002aa1n02x5               g162(.a(new_n253), .b(new_n248), .o(new_n258));
  nano22aa1n02x4               g163(.a(new_n228), .b(new_n241), .c(new_n258), .out0(new_n259));
  nanp02aa1n02x5               g164(.a(new_n185), .b(new_n259), .o1(new_n260));
  oao003aa1n02x5               g165(.a(\a[26] ), .b(\b[25] ), .c(new_n255), .carry(new_n261));
  aobi12aa1n02x5               g166(.a(new_n261), .b(new_n247), .c(new_n258), .out0(new_n262));
  xorc02aa1n02x5               g167(.a(\a[27] ), .b(\b[26] ), .out0(new_n263));
  xnbna2aa1n03x5               g168(.a(new_n263), .b(new_n260), .c(new_n262), .out0(\s[27] ));
  norp02aa1n02x5               g169(.a(\b[26] ), .b(\a[27] ), .o1(new_n265));
  160nm_ficinv00aa1n08x5       g170(.clk(new_n265), .clkout(new_n266));
  aobi12aa1n02x5               g171(.a(new_n263), .b(new_n260), .c(new_n262), .out0(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[27] ), .b(\a[28] ), .out0(new_n268));
  nano22aa1n02x4               g173(.a(new_n267), .b(new_n266), .c(new_n268), .out0(new_n269));
  160nm_ficinv00aa1n08x5       g174(.clk(new_n259), .clkout(new_n270));
  aoi012aa1n02x5               g175(.a(new_n270), .b(new_n184), .c(new_n179), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n241), .b(new_n231), .c(new_n215), .d(new_n227), .o1(new_n272));
  160nm_ficinv00aa1n08x5       g177(.clk(new_n258), .clkout(new_n273));
  aoai13aa1n02x5               g178(.a(new_n261), .b(new_n273), .c(new_n272), .d(new_n246), .o1(new_n274));
  oai012aa1n02x5               g179(.a(new_n263), .b(new_n274), .c(new_n271), .o1(new_n275));
  aoi012aa1n02x5               g180(.a(new_n268), .b(new_n275), .c(new_n266), .o1(new_n276));
  norp02aa1n02x5               g181(.a(new_n276), .b(new_n269), .o1(\s[28] ));
  norb02aa1n02x5               g182(.a(new_n263), .b(new_n268), .out0(new_n278));
  oai012aa1n02x5               g183(.a(new_n278), .b(new_n274), .c(new_n271), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[28] ), .b(\b[27] ), .c(new_n266), .carry(new_n280));
  xnrc02aa1n02x5               g185(.a(\b[28] ), .b(\a[29] ), .out0(new_n281));
  aoi012aa1n02x5               g186(.a(new_n281), .b(new_n279), .c(new_n280), .o1(new_n282));
  aobi12aa1n02x5               g187(.a(new_n278), .b(new_n260), .c(new_n262), .out0(new_n283));
  nano22aa1n02x4               g188(.a(new_n283), .b(new_n280), .c(new_n281), .out0(new_n284));
  norp02aa1n02x5               g189(.a(new_n282), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g190(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g191(.a(new_n263), .b(new_n281), .c(new_n268), .out0(new_n287));
  oai012aa1n02x5               g192(.a(new_n287), .b(new_n274), .c(new_n271), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n280), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  aobi12aa1n02x5               g196(.a(new_n287), .b(new_n260), .c(new_n262), .out0(new_n292));
  nano22aa1n02x4               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  norp02aa1n02x5               g198(.a(new_n291), .b(new_n293), .o1(\s[30] ));
  norb02aa1n02x5               g199(.a(new_n287), .b(new_n290), .out0(new_n295));
  aobi12aa1n02x5               g200(.a(new_n295), .b(new_n260), .c(new_n262), .out0(new_n296));
  oao003aa1n02x5               g201(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[30] ), .b(\a[31] ), .out0(new_n298));
  nano22aa1n02x4               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  oai012aa1n02x5               g204(.a(new_n295), .b(new_n274), .c(new_n271), .o1(new_n300));
  aoi012aa1n02x5               g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  norp02aa1n02x5               g206(.a(new_n301), .b(new_n299), .o1(\s[31] ));
  xnrb03aa1n02x5               g207(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g208(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n304));
  xorb03aa1n02x5               g209(.a(new_n304), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g210(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g211(.a(new_n122), .b(new_n123), .c(new_n111), .o1(new_n307));
  xnrb03aa1n02x5               g212(.a(new_n307), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g213(.a(\a[6] ), .b(\b[5] ), .c(new_n307), .o1(new_n309));
  xorb03aa1n02x5               g214(.a(new_n309), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g215(.a(new_n115), .b(new_n309), .c(new_n116), .o1(new_n311));
  xnrb03aa1n02x5               g216(.a(new_n311), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g217(.a(new_n146), .b(new_n120), .c(new_n126), .out0(\s[9] ));
endmodule


