// Benchmark "adder" written by ABC on Wed Jul 17 19:31:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n334, new_n335, new_n336, new_n338, new_n340,
    new_n341, new_n342, new_n343, new_n345, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1d36x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  and002aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o(new_n100));
  oaoi03aa1n12x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  xorc02aa1n12x5               g006(.a(\a[3] ), .b(\b[2] ), .out0(new_n102));
  tech160nm_finand02aa1n03p5x5 g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  orn002aa1n02x7               g008(.a(\a[4] ), .b(\b[3] ), .o(new_n104));
  oai112aa1n06x5               g009(.a(new_n104), .b(new_n103), .c(\b[2] ), .d(\a[3] ), .o1(new_n105));
  aoi012aa1d24x5               g010(.a(new_n105), .b(new_n101), .c(new_n102), .o1(new_n106));
  and002aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o(new_n107));
  nand42aa1n03x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand42aa1n06x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nano22aa1n02x4               g014(.a(new_n107), .b(new_n108), .c(new_n109), .out0(new_n110));
  nor022aa1n16x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nor002aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  aoi112aa1n02x5               g017(.a(new_n112), .b(new_n111), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  nor002aa1n04x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nor002aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand42aa1n16x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  norb03aa1n03x4               g021(.a(new_n116), .b(new_n114), .c(new_n115), .out0(new_n117));
  nand23aa1n03x5               g022(.a(new_n110), .b(new_n117), .c(new_n113), .o1(new_n118));
  nona22aa1n02x4               g023(.a(new_n116), .b(new_n115), .c(new_n114), .out0(new_n119));
  inv000aa1n02x5               g024(.a(new_n111), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  nano22aa1n06x5               g026(.a(new_n111), .b(new_n108), .c(new_n116), .out0(new_n122));
  norb02aa1n02x7               g027(.a(new_n109), .b(new_n112), .out0(new_n123));
  aoi013aa1n06x4               g028(.a(new_n121), .b(new_n119), .c(new_n122), .d(new_n123), .o1(new_n124));
  oai012aa1d24x5               g029(.a(new_n124), .b(new_n106), .c(new_n118), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  tech160nm_fixorc02aa1n03p5x5 g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n99), .c(new_n125), .d(new_n126), .o1(new_n128));
  aoi112aa1n02x5               g033(.a(new_n127), .b(new_n99), .c(new_n125), .d(new_n126), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n128), .b(new_n129), .out0(\s[10] ));
  oaoi03aa1n12x5               g035(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nor042aa1n06x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n128), .c(new_n132), .out0(\s[11] ));
  nand02aa1n03x5               g042(.a(new_n128), .b(new_n132), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n138), .b(new_n136), .o1(new_n139));
  inv000aa1n02x5               g044(.a(new_n133), .o1(new_n140));
  aoai13aa1n03x5               g045(.a(new_n140), .b(new_n135), .c(new_n128), .d(new_n132), .o1(new_n141));
  nor042aa1n03x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n04x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  aoib12aa1n02x5               g049(.a(new_n133), .b(new_n143), .c(new_n142), .out0(new_n145));
  aoi022aa1n03x5               g050(.a(new_n141), .b(new_n144), .c(new_n139), .d(new_n145), .o1(\s[12] ));
  nano23aa1d15x5               g051(.a(new_n133), .b(new_n142), .c(new_n143), .d(new_n134), .out0(new_n147));
  inv000aa1n02x5               g052(.a(new_n147), .o1(new_n148));
  nano22aa1n02x4               g053(.a(new_n148), .b(new_n126), .c(new_n127), .out0(new_n149));
  tech160nm_fioaoi03aa1n04x5   g054(.a(\a[12] ), .b(\b[11] ), .c(new_n140), .o1(new_n150));
  aoi012aa1n12x5               g055(.a(new_n150), .b(new_n147), .c(new_n131), .o1(new_n151));
  inv040aa1n03x5               g056(.a(new_n151), .o1(new_n152));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1n08x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  aoai13aa1n03x5               g060(.a(new_n155), .b(new_n152), .c(new_n125), .d(new_n149), .o1(new_n156));
  aoi112aa1n02x5               g061(.a(new_n155), .b(new_n152), .c(new_n125), .d(new_n149), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n156), .b(new_n157), .out0(\s[13] ));
  inv000aa1d42x5               g063(.a(new_n153), .o1(new_n159));
  nor042aa1n04x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n06x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n156), .c(new_n159), .out0(\s[14] ));
  nano23aa1n06x5               g068(.a(new_n153), .b(new_n160), .c(new_n161), .d(new_n154), .out0(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n152), .c(new_n125), .d(new_n149), .o1(new_n165));
  oaoi03aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .c(new_n159), .o1(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  xorc02aa1n12x5               g072(.a(\a[15] ), .b(\b[14] ), .out0(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n165), .c(new_n167), .out0(\s[15] ));
  nand42aa1n02x5               g074(.a(new_n165), .b(new_n167), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(new_n170), .b(new_n168), .o1(new_n171));
  inv000aa1d42x5               g076(.a(\a[15] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(\b[14] ), .o1(new_n173));
  nanp02aa1n02x5               g078(.a(new_n173), .b(new_n172), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n168), .o1(new_n175));
  aoai13aa1n02x7               g080(.a(new_n174), .b(new_n175), .c(new_n165), .d(new_n167), .o1(new_n176));
  xorc02aa1n12x5               g081(.a(\a[16] ), .b(\b[15] ), .out0(new_n177));
  inv000aa1d42x5               g082(.a(\a[16] ), .o1(new_n178));
  inv000aa1d42x5               g083(.a(\b[15] ), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(new_n179), .b(new_n178), .o1(new_n180));
  and002aa1n02x5               g085(.a(\b[15] ), .b(\a[16] ), .o(new_n181));
  aboi22aa1n03x5               g086(.a(new_n181), .b(new_n180), .c(new_n173), .d(new_n172), .out0(new_n182));
  aoi022aa1n02x5               g087(.a(new_n176), .b(new_n177), .c(new_n171), .d(new_n182), .o1(\s[16] ));
  nanp03aa1d12x5               g088(.a(new_n164), .b(new_n168), .c(new_n177), .o1(new_n184));
  nano32aa1n09x5               g089(.a(new_n184), .b(new_n147), .c(new_n127), .d(new_n126), .out0(new_n185));
  nanp02aa1n06x5               g090(.a(new_n125), .b(new_n185), .o1(new_n186));
  nanp02aa1n02x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  oai112aa1n03x5               g092(.a(new_n161), .b(new_n187), .c(new_n160), .d(new_n153), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n180), .b(new_n181), .c(new_n188), .d(new_n174), .o1(new_n189));
  oab012aa1n06x5               g094(.a(new_n189), .b(new_n151), .c(new_n184), .out0(new_n190));
  xorc02aa1n12x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n186), .c(new_n190), .out0(\s[17] ));
  inv040aa1d28x5               g097(.a(\a[17] ), .o1(new_n193));
  inv040aa1d32x5               g098(.a(\b[16] ), .o1(new_n194));
  nanp02aa1n02x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  nand02aa1n02x5               g100(.a(new_n188), .b(new_n174), .o1(new_n196));
  tech160nm_fioaoi03aa1n03p5x5 g101(.a(new_n178), .b(new_n179), .c(new_n196), .o1(new_n197));
  oai012aa1d24x5               g102(.a(new_n197), .b(new_n151), .c(new_n184), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n191), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n199));
  nor002aa1d32x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nand42aa1d28x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  norb02aa1n03x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n199), .c(new_n195), .out0(\s[18] ));
  nanp02aa1n02x5               g108(.a(\b[16] ), .b(\a[17] ), .o1(new_n204));
  nano32aa1n02x4               g109(.a(new_n200), .b(new_n195), .c(new_n201), .d(new_n204), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n206));
  aoai13aa1n12x5               g111(.a(new_n201), .b(new_n200), .c(new_n193), .d(new_n194), .o1(new_n207));
  nor002aa1n16x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nanp02aa1n09x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nanb02aa1n06x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n206), .c(new_n207), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n08x5               g118(.a(new_n186), .b(new_n190), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n207), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n211), .b(new_n215), .c(new_n214), .d(new_n205), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n208), .o1(new_n217));
  aoai13aa1n02x7               g122(.a(new_n217), .b(new_n210), .c(new_n206), .d(new_n207), .o1(new_n218));
  inv000aa1d42x5               g123(.a(\a[20] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(\b[19] ), .o1(new_n220));
  nand22aa1n03x5               g125(.a(new_n220), .b(new_n219), .o1(new_n221));
  nand02aa1n06x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand02aa1n03x5               g127(.a(new_n221), .b(new_n222), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoi012aa1n02x5               g129(.a(new_n208), .b(new_n221), .c(new_n222), .o1(new_n225));
  aoi022aa1n03x5               g130(.a(new_n218), .b(new_n224), .c(new_n216), .d(new_n225), .o1(\s[20] ));
  nor002aa1n03x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nano23aa1n06x5               g132(.a(new_n208), .b(new_n227), .c(new_n222), .d(new_n209), .out0(new_n228));
  nand23aa1n04x5               g133(.a(new_n228), .b(new_n191), .c(new_n202), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n231));
  nona23aa1n09x5               g136(.a(new_n222), .b(new_n209), .c(new_n208), .d(new_n227), .out0(new_n232));
  aob012aa1n02x5               g137(.a(new_n221), .b(new_n208), .c(new_n222), .out0(new_n233));
  oabi12aa1n18x5               g138(.a(new_n233), .b(new_n232), .c(new_n207), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  nor002aa1d32x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  tech160nm_finand02aa1n03p5x5 g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  xnbna2aa1n03x5               g143(.a(new_n238), .b(new_n231), .c(new_n235), .out0(\s[21] ));
  aoai13aa1n03x5               g144(.a(new_n238), .b(new_n234), .c(new_n214), .d(new_n230), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n236), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n238), .o1(new_n242));
  aoai13aa1n02x7               g147(.a(new_n241), .b(new_n242), .c(new_n231), .d(new_n235), .o1(new_n243));
  nor022aa1n06x5               g148(.a(\b[21] ), .b(\a[22] ), .o1(new_n244));
  nand22aa1n04x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  aoib12aa1n02x5               g151(.a(new_n236), .b(new_n245), .c(new_n244), .out0(new_n247));
  aoi022aa1n03x5               g152(.a(new_n243), .b(new_n246), .c(new_n240), .d(new_n247), .o1(\s[22] ));
  nona23aa1d18x5               g153(.a(new_n245), .b(new_n237), .c(new_n236), .d(new_n244), .out0(new_n249));
  nano23aa1n02x4               g154(.a(new_n249), .b(new_n232), .c(new_n191), .d(new_n202), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n249), .o1(new_n252));
  aoi012aa1n02x5               g157(.a(new_n244), .b(new_n236), .c(new_n245), .o1(new_n253));
  aobi12aa1n02x5               g158(.a(new_n253), .b(new_n234), .c(new_n252), .out0(new_n254));
  orn002aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .o(new_n255));
  nand42aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  nanp02aa1n09x5               g161(.a(new_n255), .b(new_n256), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xnbna2aa1n03x5               g163(.a(new_n258), .b(new_n251), .c(new_n254), .out0(\s[23] ));
  nand42aa1n02x5               g164(.a(new_n251), .b(new_n254), .o1(new_n260));
  nand02aa1n02x5               g165(.a(new_n260), .b(new_n258), .o1(new_n261));
  aoai13aa1n02x7               g166(.a(new_n255), .b(new_n257), .c(new_n251), .d(new_n254), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[23] ), .b(\a[24] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  and002aa1n02x5               g169(.a(new_n263), .b(new_n255), .o(new_n265));
  aoi022aa1n03x5               g170(.a(new_n262), .b(new_n264), .c(new_n261), .d(new_n265), .o1(\s[24] ));
  norp02aa1n02x5               g171(.a(new_n263), .b(new_n257), .o1(new_n267));
  nano22aa1n06x5               g172(.a(new_n229), .b(new_n252), .c(new_n267), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n269));
  norp02aa1n02x5               g174(.a(\b[23] ), .b(\a[24] ), .o1(new_n270));
  nor043aa1n02x5               g175(.a(new_n249), .b(new_n257), .c(new_n263), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n256), .b(new_n244), .c(new_n236), .d(new_n245), .o1(new_n272));
  aoi022aa1n02x5               g177(.a(new_n272), .b(new_n255), .c(\a[24] ), .d(\b[23] ), .o1(new_n273));
  aoi112aa1n06x5               g178(.a(new_n270), .b(new_n273), .c(new_n234), .d(new_n271), .o1(new_n274));
  xnrc02aa1n12x5               g179(.a(\b[24] ), .b(\a[25] ), .out0(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n269), .c(new_n274), .out0(\s[25] ));
  norp03aa1n06x5               g182(.a(new_n207), .b(new_n210), .c(new_n223), .o1(new_n278));
  oai012aa1n03x5               g183(.a(new_n271), .b(new_n278), .c(new_n233), .o1(new_n279));
  nona22aa1n03x5               g184(.a(new_n279), .b(new_n273), .c(new_n270), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n276), .b(new_n280), .c(new_n214), .d(new_n268), .o1(new_n281));
  nor042aa1n06x5               g186(.a(\b[24] ), .b(\a[25] ), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  aoai13aa1n02x7               g188(.a(new_n283), .b(new_n275), .c(new_n269), .d(new_n274), .o1(new_n284));
  tech160nm_fixorc02aa1n02p5x5 g189(.a(\a[26] ), .b(\b[25] ), .out0(new_n285));
  norp02aa1n02x5               g190(.a(new_n285), .b(new_n282), .o1(new_n286));
  aoi022aa1n03x5               g191(.a(new_n284), .b(new_n285), .c(new_n281), .d(new_n286), .o1(\s[26] ));
  norb02aa1n06x5               g192(.a(new_n285), .b(new_n275), .out0(new_n288));
  nano22aa1n06x5               g193(.a(new_n229), .b(new_n271), .c(new_n288), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n198), .c(new_n125), .d(new_n185), .o1(new_n290));
  oao003aa1n12x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n283), .carry(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoi012aa1n06x5               g197(.a(new_n292), .b(new_n280), .c(new_n288), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(new_n290), .out0(\s[27] ));
  inv000aa1d42x5               g200(.a(new_n288), .o1(new_n296));
  oaih12aa1n06x5               g201(.a(new_n291), .b(new_n274), .c(new_n296), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n294), .b(new_n297), .c(new_n214), .d(new_n289), .o1(new_n298));
  norp02aa1n02x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  inv000aa1n03x5               g204(.a(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n294), .o1(new_n301));
  aoai13aa1n02x7               g206(.a(new_n300), .b(new_n301), .c(new_n293), .d(new_n290), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(new_n303), .b(new_n299), .o1(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n298), .d(new_n304), .o1(\s[28] ));
  and002aa1n02x5               g210(.a(new_n303), .b(new_n294), .o(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n297), .c(new_n214), .d(new_n289), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n306), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[28] ), .b(\b[27] ), .c(new_n300), .carry(new_n309));
  aoai13aa1n02x7               g214(.a(new_n309), .b(new_n308), .c(new_n293), .d(new_n290), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  norb02aa1n02x5               g216(.a(new_n309), .b(new_n311), .out0(new_n312));
  aoi022aa1n03x5               g217(.a(new_n310), .b(new_n311), .c(new_n307), .d(new_n312), .o1(\s[29] ));
  xnrb03aa1n02x5               g218(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g219(.a(new_n301), .b(new_n303), .c(new_n311), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n297), .c(new_n214), .d(new_n289), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n315), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .carry(new_n318));
  aoai13aa1n02x7               g223(.a(new_n318), .b(new_n317), .c(new_n293), .d(new_n290), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .out0(new_n320));
  norb02aa1n02x5               g225(.a(new_n318), .b(new_n320), .out0(new_n321));
  aoi022aa1n03x5               g226(.a(new_n319), .b(new_n320), .c(new_n316), .d(new_n321), .o1(\s[30] ));
  xorc02aa1n02x5               g227(.a(\a[31] ), .b(\b[30] ), .out0(new_n323));
  nano32aa1n03x7               g228(.a(new_n301), .b(new_n320), .c(new_n303), .d(new_n311), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n297), .c(new_n214), .d(new_n289), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n324), .o1(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n318), .carry(new_n327));
  aoai13aa1n02x7               g232(.a(new_n327), .b(new_n326), .c(new_n293), .d(new_n290), .o1(new_n328));
  and002aa1n02x5               g233(.a(\b[29] ), .b(\a[30] ), .o(new_n329));
  oabi12aa1n02x5               g234(.a(new_n323), .b(\a[30] ), .c(\b[29] ), .out0(new_n330));
  oab012aa1n02x4               g235(.a(new_n330), .b(new_n318), .c(new_n329), .out0(new_n331));
  aoi022aa1n03x5               g236(.a(new_n328), .b(new_n323), .c(new_n325), .d(new_n331), .o1(\s[31] ));
  xorb03aa1n02x5               g237(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g238(.a(new_n106), .o1(new_n334));
  norp02aa1n02x5               g239(.a(\b[2] ), .b(\a[3] ), .o1(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n101), .c(new_n102), .o1(new_n336));
  aoai13aa1n02x5               g241(.a(new_n334), .b(new_n336), .c(new_n104), .d(new_n103), .o1(\s[4] ));
  norp02aa1n02x5               g242(.a(new_n107), .b(new_n114), .o1(new_n338));
  xobna2aa1n03x5               g243(.a(new_n338), .b(new_n334), .c(new_n103), .out0(\s[5] ));
  norb02aa1n02x5               g244(.a(new_n116), .b(new_n115), .out0(new_n340));
  aoi013aa1n02x4               g245(.a(new_n114), .b(new_n334), .c(new_n103), .d(new_n338), .o1(new_n341));
  nanb03aa1n02x5               g246(.a(new_n106), .b(new_n338), .c(new_n103), .out0(new_n342));
  nanp02aa1n03x5               g247(.a(new_n342), .b(new_n117), .o1(new_n343));
  oai012aa1n02x5               g248(.a(new_n343), .b(new_n341), .c(new_n340), .o1(\s[6] ));
  aoi022aa1n02x5               g249(.a(new_n343), .b(new_n116), .c(new_n108), .d(new_n120), .o1(new_n345));
  aoi012aa1n02x5               g250(.a(new_n345), .b(new_n122), .c(new_n343), .o1(\s[7] ));
  nanp02aa1n02x5               g251(.a(new_n343), .b(new_n122), .o1(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n123), .b(new_n347), .c(new_n120), .out0(\s[8] ));
  xorb03aa1n02x5               g253(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


