// Benchmark "adder" written by ABC on Thu Jul 18 13:00:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n131, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n319, new_n322, new_n324, new_n325, new_n326, new_n328,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n03x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  nanp02aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  norp02aa1n24x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nor022aa1n08x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  oai012aa1n02x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n12x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor002aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  tech160nm_fioai012aa1n05x5   g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n02x4               g011(.a(new_n98), .b(new_n106), .c(new_n100), .d(new_n99), .out0(new_n107));
  oai012aa1n04x7               g012(.a(new_n101), .b(new_n107), .c(new_n105), .o1(new_n108));
  nor042aa1n06x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nand42aa1n04x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nor042aa1n06x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nona23aa1n03x5               g017(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n113));
  xnrc02aa1n12x5               g018(.a(\b[7] ), .b(\a[8] ), .out0(new_n114));
  xnrc02aa1n12x5               g019(.a(\b[6] ), .b(\a[7] ), .out0(new_n115));
  nor043aa1n02x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  norp02aa1n02x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  tech160nm_fioai012aa1n03p5x5 g023(.a(new_n117), .b(new_n114), .c(new_n118), .o1(new_n119));
  oaih12aa1n06x5               g024(.a(new_n110), .b(new_n111), .c(new_n109), .o1(new_n120));
  oai013aa1n09x5               g025(.a(new_n119), .b(new_n115), .c(new_n114), .d(new_n120), .o1(new_n121));
  xorc02aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .out0(new_n122));
  aoai13aa1n02x5               g027(.a(new_n122), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n123));
  xorc02aa1n12x5               g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  xnbna2aa1n03x5               g029(.a(new_n124), .b(new_n123), .c(new_n97), .out0(\s[10] ));
  inv000aa1d42x5               g030(.a(new_n124), .o1(new_n126));
  oai022aa1n02x7               g031(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  aob012aa1n03x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n126), .c(new_n123), .d(new_n97), .o1(new_n129));
  xorb03aa1n02x5               g034(.a(new_n129), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1d18x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nand02aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  nor042aa1d18x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  nand02aa1d10x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  aoai13aa1n02x5               g041(.a(new_n136), .b(new_n131), .c(new_n129), .d(new_n133), .o1(new_n137));
  nona22aa1n02x4               g042(.a(new_n135), .b(new_n134), .c(new_n131), .out0(new_n138));
  aoai13aa1n02x5               g043(.a(new_n137), .b(new_n138), .c(new_n133), .d(new_n129), .o1(\s[12] ));
  nona23aa1n09x5               g044(.a(new_n135), .b(new_n132), .c(new_n131), .d(new_n134), .out0(new_n140));
  nano22aa1n02x4               g045(.a(new_n140), .b(new_n122), .c(new_n124), .out0(new_n141));
  aoai13aa1n03x5               g046(.a(new_n141), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n142));
  oai012aa1d24x5               g047(.a(new_n135), .b(new_n134), .c(new_n131), .o1(new_n143));
  tech160nm_fioai012aa1n05x5   g048(.a(new_n143), .b(new_n140), .c(new_n128), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n144), .b(new_n142), .out0(new_n145));
  xorb03aa1n02x5               g050(.a(new_n145), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g051(.a(\b[12] ), .b(\a[13] ), .o1(new_n147));
  nand42aa1d28x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  nanb02aa1n02x5               g053(.a(new_n147), .b(new_n148), .out0(new_n149));
  aoib12aa1n02x5               g054(.a(new_n149), .b(new_n142), .c(new_n144), .out0(new_n150));
  nor002aa1n16x5               g055(.a(\b[13] ), .b(\a[14] ), .o1(new_n151));
  nand42aa1d28x5               g056(.a(\b[13] ), .b(\a[14] ), .o1(new_n152));
  obai22aa1n02x7               g057(.a(new_n152), .b(new_n151), .c(new_n150), .d(new_n147), .out0(new_n153));
  norb03aa1n02x5               g058(.a(new_n152), .b(new_n147), .c(new_n151), .out0(new_n154));
  oaib12aa1n02x5               g059(.a(new_n153), .b(new_n150), .c(new_n154), .out0(\s[14] ));
  nano23aa1d15x5               g060(.a(new_n147), .b(new_n151), .c(new_n152), .d(new_n148), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  oaoi03aa1n03x5               g062(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n158));
  nano23aa1n09x5               g063(.a(new_n131), .b(new_n134), .c(new_n135), .d(new_n132), .out0(new_n159));
  inv000aa1n02x5               g064(.a(new_n143), .o1(new_n160));
  aoai13aa1n06x5               g065(.a(new_n156), .b(new_n160), .c(new_n159), .d(new_n158), .o1(new_n161));
  oai012aa1n12x5               g066(.a(new_n152), .b(new_n151), .c(new_n147), .o1(new_n162));
  oai112aa1n03x5               g067(.a(new_n161), .b(new_n162), .c(new_n142), .d(new_n157), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n09x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand02aa1n02x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  nor042aa1n04x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  nanp02aa1n03x5               g073(.a(\b[15] ), .b(\a[16] ), .o1(new_n169));
  nanb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n171));
  nona22aa1n02x4               g076(.a(new_n169), .b(new_n168), .c(new_n165), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n171), .b(new_n172), .c(new_n167), .d(new_n163), .o1(\s[16] ));
  nano23aa1n06x5               g078(.a(new_n165), .b(new_n168), .c(new_n169), .d(new_n166), .out0(new_n174));
  nand02aa1n02x5               g079(.a(new_n174), .b(new_n156), .o1(new_n175));
  nano32aa1n03x7               g080(.a(new_n175), .b(new_n159), .c(new_n124), .d(new_n122), .out0(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n177));
  inv000aa1n02x5               g082(.a(new_n162), .o1(new_n178));
  aoai13aa1n06x5               g083(.a(new_n174), .b(new_n178), .c(new_n144), .d(new_n156), .o1(new_n179));
  oa0012aa1n06x5               g084(.a(new_n169), .b(new_n168), .c(new_n165), .o(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  nanp03aa1d12x5               g086(.a(new_n177), .b(new_n179), .c(new_n181), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(\a[17] ), .b(new_n184), .out0(new_n185));
  xnrc02aa1n02x5               g090(.a(\b[16] ), .b(\a[17] ), .out0(new_n186));
  nanb02aa1n02x5               g091(.a(new_n186), .b(new_n182), .out0(new_n187));
  xorc02aa1n02x5               g092(.a(\a[18] ), .b(\b[17] ), .out0(new_n188));
  inv000aa1n02x5               g093(.a(new_n174), .o1(new_n189));
  aoai13aa1n12x5               g094(.a(new_n181), .b(new_n189), .c(new_n161), .d(new_n162), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n190), .o1(new_n191));
  oai022aa1n04x7               g096(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n192));
  aoi012aa1n02x5               g097(.a(new_n192), .b(\a[18] ), .c(\b[17] ), .o1(new_n193));
  aoai13aa1n02x5               g098(.a(new_n193), .b(new_n186), .c(new_n191), .d(new_n177), .o1(new_n194));
  aoai13aa1n02x5               g099(.a(new_n194), .b(new_n188), .c(new_n187), .d(new_n185), .o1(\s[18] ));
  nanp02aa1n02x5               g100(.a(new_n108), .b(new_n116), .o1(new_n196));
  nanb02aa1n02x5               g101(.a(new_n121), .b(new_n196), .out0(new_n197));
  inv000aa1d42x5               g102(.a(\b[17] ), .o1(new_n198));
  xroi22aa1d06x4               g103(.a(new_n198), .b(\a[18] ), .c(new_n184), .d(\a[17] ), .out0(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n190), .c(new_n197), .d(new_n176), .o1(new_n200));
  oaib12aa1n09x5               g105(.a(new_n192), .b(new_n198), .c(\a[18] ), .out0(new_n201));
  nor002aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand42aa1n04x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nanb02aa1n02x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  xobna2aa1n03x5               g109(.a(new_n204), .b(new_n200), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n03x5               g111(.a(new_n200), .b(new_n201), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nanp02aa1n04x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n202), .c(new_n207), .d(new_n203), .o1(new_n211));
  norb03aa1n02x5               g116(.a(new_n209), .b(new_n202), .c(new_n208), .out0(new_n212));
  aoai13aa1n02x5               g117(.a(new_n212), .b(new_n204), .c(new_n200), .d(new_n201), .o1(new_n213));
  nanp02aa1n03x5               g118(.a(new_n211), .b(new_n213), .o1(\s[20] ));
  nona23aa1n09x5               g119(.a(new_n209), .b(new_n203), .c(new_n202), .d(new_n208), .out0(new_n215));
  norb03aa1n02x5               g120(.a(new_n188), .b(new_n215), .c(new_n186), .out0(new_n216));
  tech160nm_fioai012aa1n05x5   g121(.a(new_n209), .b(new_n208), .c(new_n202), .o1(new_n217));
  oai012aa1n12x5               g122(.a(new_n217), .b(new_n215), .c(new_n201), .o1(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n09x5               g125(.a(new_n220), .b(new_n218), .c(new_n182), .d(new_n216), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(new_n220), .b(new_n218), .c(new_n182), .d(new_n216), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n221), .b(new_n222), .out0(\s[21] ));
  nor042aa1n06x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  xorc02aa1n02x5               g130(.a(\a[22] ), .b(\b[21] ), .out0(new_n226));
  nanp02aa1n02x5               g131(.a(\b[21] ), .b(\a[22] ), .o1(new_n227));
  oai022aa1n02x5               g132(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n228));
  nanb03aa1n03x5               g133(.a(new_n228), .b(new_n221), .c(new_n227), .out0(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n226), .c(new_n225), .d(new_n221), .o1(\s[22] ));
  nano23aa1n06x5               g135(.a(new_n202), .b(new_n208), .c(new_n209), .d(new_n203), .out0(new_n231));
  orn002aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .o(new_n232));
  nano22aa1n12x5               g137(.a(new_n219), .b(new_n232), .c(new_n227), .out0(new_n233));
  nanp03aa1d12x5               g138(.a(new_n199), .b(new_n233), .c(new_n231), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  oaoi03aa1n02x5               g140(.a(\a[18] ), .b(\b[17] ), .c(new_n185), .o1(new_n236));
  inv000aa1n02x5               g141(.a(new_n217), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n233), .b(new_n237), .c(new_n231), .d(new_n236), .o1(new_n238));
  oaoi03aa1n09x5               g143(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nanp02aa1n02x5               g145(.a(new_n238), .b(new_n240), .o1(new_n241));
  xnrc02aa1n12x5               g146(.a(\b[22] ), .b(\a[23] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n241), .c(new_n182), .d(new_n235), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(new_n243), .b(new_n241), .c(new_n182), .d(new_n235), .o1(new_n245));
  norb02aa1n03x4               g150(.a(new_n244), .b(new_n245), .out0(\s[23] ));
  nor002aa1n03x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  xorc02aa1n02x5               g153(.a(\a[24] ), .b(\b[23] ), .out0(new_n249));
  inv000aa1d42x5               g154(.a(\a[24] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[23] ), .o1(new_n251));
  aoi012aa1n02x5               g156(.a(new_n247), .b(new_n250), .c(new_n251), .o1(new_n252));
  oai112aa1n03x5               g157(.a(new_n244), .b(new_n252), .c(new_n251), .d(new_n250), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n249), .c(new_n248), .d(new_n244), .o1(\s[24] ));
  norb02aa1n09x5               g159(.a(new_n249), .b(new_n242), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  nano32aa1n02x4               g161(.a(new_n256), .b(new_n199), .c(new_n233), .d(new_n231), .out0(new_n257));
  oaoi03aa1n02x5               g162(.a(new_n250), .b(new_n251), .c(new_n247), .o1(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n256), .c(new_n238), .d(new_n240), .o1(new_n259));
  xorc02aa1n12x5               g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n259), .c(new_n182), .d(new_n257), .o1(new_n261));
  aoi112aa1n02x5               g166(.a(new_n260), .b(new_n259), .c(new_n182), .d(new_n257), .o1(new_n262));
  norb02aa1n03x4               g167(.a(new_n261), .b(new_n262), .out0(\s[25] ));
  nor042aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  inv000aa1d42x5               g171(.a(\a[26] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(\b[25] ), .o1(new_n268));
  aoi012aa1n02x5               g173(.a(new_n264), .b(new_n267), .c(new_n268), .o1(new_n269));
  oai112aa1n03x5               g174(.a(new_n261), .b(new_n269), .c(new_n268), .d(new_n267), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n266), .c(new_n265), .d(new_n261), .o1(\s[26] ));
  and002aa1n06x5               g176(.a(new_n266), .b(new_n260), .o(new_n272));
  nano22aa1d15x5               g177(.a(new_n234), .b(new_n272), .c(new_n255), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n190), .c(new_n197), .d(new_n176), .o1(new_n274));
  oaoi03aa1n02x5               g179(.a(new_n267), .b(new_n268), .c(new_n264), .o1(new_n275));
  aobi12aa1n06x5               g180(.a(new_n275), .b(new_n259), .c(new_n272), .out0(new_n276));
  xorc02aa1n02x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n274), .c(new_n276), .out0(\s[27] ));
  xorc02aa1n02x5               g183(.a(\a[28] ), .b(\b[27] ), .out0(new_n279));
  inv020aa1n03x5               g184(.a(new_n273), .o1(new_n280));
  aoi013aa1n02x4               g185(.a(new_n280), .b(new_n177), .c(new_n179), .d(new_n181), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n255), .b(new_n239), .c(new_n218), .d(new_n233), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n272), .o1(new_n283));
  aoai13aa1n12x5               g188(.a(new_n275), .b(new_n283), .c(new_n282), .d(new_n258), .o1(new_n284));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  oaoi13aa1n02x5               g190(.a(new_n285), .b(new_n277), .c(new_n281), .d(new_n284), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n277), .b(new_n284), .c(new_n182), .d(new_n273), .o1(new_n287));
  oai112aa1n03x5               g192(.a(new_n287), .b(new_n279), .c(\b[26] ), .d(\a[27] ), .o1(new_n288));
  oai012aa1n03x5               g193(.a(new_n288), .b(new_n286), .c(new_n279), .o1(\s[28] ));
  and002aa1n02x5               g194(.a(new_n279), .b(new_n277), .o(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n284), .c(new_n182), .d(new_n273), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .out0(new_n292));
  inv000aa1d42x5               g197(.a(\a[28] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  aoi112aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n295));
  aoi112aa1n02x5               g200(.a(new_n292), .b(new_n295), .c(new_n293), .d(new_n294), .o1(new_n296));
  aoi012aa1n02x5               g201(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n297));
  nanp02aa1n03x5               g202(.a(new_n291), .b(new_n297), .o1(new_n298));
  aoi022aa1n02x7               g203(.a(new_n298), .b(new_n292), .c(new_n291), .d(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g205(.a(new_n277), .b(new_n292), .c(new_n279), .o(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n284), .c(new_n182), .d(new_n273), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .o1(new_n304));
  aoi012aa1n02x5               g209(.a(new_n297), .b(\a[29] ), .c(\b[28] ), .o1(new_n305));
  norp03aa1n02x5               g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n307));
  nanp02aa1n03x5               g212(.a(new_n302), .b(new_n307), .o1(new_n308));
  aoi022aa1n02x7               g213(.a(new_n308), .b(new_n303), .c(new_n302), .d(new_n306), .o1(\s[30] ));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  and003aa1n02x5               g215(.a(new_n290), .b(new_n303), .c(new_n292), .o(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n284), .c(new_n182), .d(new_n273), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n313));
  aoi012aa1n03x5               g218(.a(new_n310), .b(new_n312), .c(new_n313), .o1(new_n314));
  aobi12aa1n03x5               g219(.a(new_n311), .b(new_n274), .c(new_n276), .out0(new_n315));
  nano22aa1n03x5               g220(.a(new_n315), .b(new_n310), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[31] ));
  xnrb03aa1n02x5               g222(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g223(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g225(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g226(.a(new_n111), .b(new_n108), .c(new_n112), .o1(new_n322));
  xnrb03aa1n02x5               g227(.a(new_n322), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g228(.a(new_n109), .b(new_n110), .out0(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n115), .b(new_n120), .c(new_n322), .d(new_n324), .o1(new_n325));
  oai112aa1n02x5               g230(.a(new_n120), .b(new_n115), .c(new_n322), .d(new_n324), .o1(new_n326));
  norb02aa1n02x5               g231(.a(new_n326), .b(new_n325), .out0(\s[7] ));
  oabi12aa1n02x5               g232(.a(new_n114), .b(\a[7] ), .c(\b[6] ), .out0(new_n328));
  oai012aa1n02x5               g233(.a(new_n114), .b(new_n325), .c(new_n118), .o1(new_n329));
  oai012aa1n02x5               g234(.a(new_n329), .b(new_n325), .c(new_n328), .o1(\s[8] ));
  xorb03aa1n02x5               g235(.a(new_n197), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


