// Benchmark "adder" written by ABC on Wed Jul 17 18:10:07 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n131, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n295, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n316,
    new_n318, new_n319, new_n320, new_n321, new_n323, new_n324, new_n326,
    new_n327, new_n329, new_n330, new_n332, new_n334, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n09x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  oai112aa1n06x5               g002(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n98));
  nand42aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  norp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  aoi113aa1n09x5               g007(.a(new_n102), .b(new_n100), .c(new_n98), .d(new_n101), .e(new_n99), .o1(new_n103));
  and002aa1n03x5               g008(.a(\b[4] ), .b(\a[5] ), .o(new_n104));
  nor042aa1n06x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  aoi112aa1n03x5               g010(.a(new_n104), .b(new_n105), .c(\a[4] ), .d(\b[3] ), .o1(new_n106));
  tech160nm_fixorc02aa1n02p5x5 g011(.a(\a[8] ), .b(\b[7] ), .out0(new_n107));
  nor002aa1n16x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand42aa1n03x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nano23aa1n02x4               g016(.a(new_n108), .b(new_n110), .c(new_n111), .d(new_n109), .out0(new_n112));
  nand23aa1n03x5               g017(.a(new_n112), .b(new_n106), .c(new_n107), .o1(new_n113));
  norb02aa1n02x7               g018(.a(new_n109), .b(new_n108), .out0(new_n114));
  inv000aa1n09x5               g019(.a(new_n105), .o1(new_n115));
  oaoi03aa1n12x5               g020(.a(\a[6] ), .b(\b[5] ), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(new_n108), .o1(new_n117));
  oaoi03aa1n02x5               g022(.a(\a[8] ), .b(\b[7] ), .c(new_n117), .o1(new_n118));
  aoi013aa1n06x4               g023(.a(new_n118), .b(new_n116), .c(new_n107), .d(new_n114), .o1(new_n119));
  oai012aa1d24x5               g024(.a(new_n119), .b(new_n113), .c(new_n103), .o1(new_n120));
  xorc02aa1n02x5               g025(.a(\a[9] ), .b(\b[8] ), .out0(new_n121));
  xorc02aa1n02x5               g026(.a(\a[10] ), .b(\b[9] ), .out0(new_n122));
  aoai13aa1n04x5               g027(.a(new_n122), .b(new_n97), .c(new_n120), .d(new_n121), .o1(new_n123));
  aoi112aa1n02x5               g028(.a(new_n122), .b(new_n97), .c(new_n120), .d(new_n121), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n123), .b(new_n124), .out0(\s[10] ));
  inv040aa1n03x5               g030(.a(new_n97), .o1(new_n126));
  oaoi03aa1n12x5               g031(.a(\a[10] ), .b(\b[9] ), .c(new_n126), .o1(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[11] ), .b(\b[10] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n123), .c(new_n128), .out0(\s[11] ));
  aob012aa1n03x5               g035(.a(new_n129), .b(new_n123), .c(new_n128), .out0(new_n131));
  xorc02aa1n02x5               g036(.a(\a[12] ), .b(\b[11] ), .out0(new_n132));
  nor042aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norp02aa1n02x5               g038(.a(new_n132), .b(new_n133), .o1(new_n134));
  inv040aa1n03x5               g039(.a(new_n133), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n129), .o1(new_n136));
  aoai13aa1n02x5               g041(.a(new_n135), .b(new_n136), .c(new_n123), .d(new_n128), .o1(new_n137));
  aoi022aa1n02x5               g042(.a(new_n137), .b(new_n132), .c(new_n131), .d(new_n134), .o1(\s[12] ));
  nano32aa1n02x4               g043(.a(new_n136), .b(new_n132), .c(new_n121), .d(new_n122), .out0(new_n139));
  nanp02aa1n02x5               g044(.a(new_n120), .b(new_n139), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  xnrc02aa1n02x5               g046(.a(\b[11] ), .b(\a[12] ), .out0(new_n142));
  nano22aa1n02x4               g047(.a(new_n142), .b(new_n135), .c(new_n141), .out0(new_n143));
  oao003aa1n02x5               g048(.a(\a[12] ), .b(\b[11] ), .c(new_n135), .carry(new_n144));
  inv000aa1n02x5               g049(.a(new_n144), .o1(new_n145));
  tech160nm_fiaoi012aa1n05x5   g050(.a(new_n145), .b(new_n143), .c(new_n127), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(new_n140), .b(new_n146), .o1(new_n147));
  xnrc02aa1n12x5               g052(.a(\b[12] ), .b(\a[13] ), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoi112aa1n02x5               g054(.a(new_n145), .b(new_n149), .c(new_n143), .d(new_n127), .o1(new_n150));
  aoi022aa1n02x5               g055(.a(new_n147), .b(new_n149), .c(new_n140), .d(new_n150), .o1(\s[13] ));
  nor042aa1n03x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  inv000aa1n03x5               g057(.a(new_n152), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n146), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n149), .b(new_n154), .c(new_n120), .d(new_n139), .o1(new_n155));
  xorc02aa1n12x5               g060(.a(\a[14] ), .b(\b[13] ), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n155), .c(new_n153), .out0(\s[14] ));
  norb02aa1n02x5               g062(.a(new_n156), .b(new_n148), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n154), .c(new_n120), .d(new_n139), .o1(new_n159));
  oaoi03aa1n09x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n153), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  xorc02aa1n02x5               g066(.a(\a[15] ), .b(\b[14] ), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n159), .c(new_n161), .out0(\s[15] ));
  aoai13aa1n04x5               g068(.a(new_n162), .b(new_n160), .c(new_n147), .d(new_n158), .o1(new_n164));
  tech160nm_fixorc02aa1n04x5   g069(.a(\a[16] ), .b(\b[15] ), .out0(new_n165));
  nor042aa1n03x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  norp02aa1n02x5               g071(.a(new_n165), .b(new_n166), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n166), .o1(new_n168));
  xnrc02aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n168), .b(new_n169), .c(new_n159), .d(new_n161), .o1(new_n170));
  aoi022aa1n03x5               g075(.a(new_n170), .b(new_n165), .c(new_n164), .d(new_n167), .o1(\s[16] ));
  nona23aa1n09x5               g076(.a(new_n165), .b(new_n156), .c(new_n148), .d(new_n169), .out0(new_n172));
  nano32aa1n03x7               g077(.a(new_n172), .b(new_n143), .c(new_n122), .d(new_n121), .out0(new_n173));
  nanp02aa1n06x5               g078(.a(new_n173), .b(new_n120), .o1(new_n174));
  nanp03aa1n02x5               g079(.a(new_n127), .b(new_n129), .c(new_n132), .o1(new_n175));
  oaoi03aa1n02x5               g080(.a(\a[16] ), .b(\b[15] ), .c(new_n168), .o1(new_n176));
  aoi013aa1n02x4               g081(.a(new_n176), .b(new_n160), .c(new_n162), .d(new_n165), .o1(new_n177));
  aoai13aa1n12x5               g082(.a(new_n177), .b(new_n172), .c(new_n175), .d(new_n144), .o1(new_n178));
  nanb02aa1n06x5               g083(.a(new_n178), .b(new_n174), .out0(new_n179));
  tech160nm_fixorc02aa1n04x5   g084(.a(\a[17] ), .b(\b[16] ), .out0(new_n180));
  aoi113aa1n02x5               g085(.a(new_n176), .b(new_n180), .c(new_n160), .d(new_n162), .e(new_n165), .o1(new_n181));
  oa0012aa1n02x5               g086(.a(new_n181), .b(new_n146), .c(new_n172), .o(new_n182));
  aoi022aa1n02x5               g087(.a(new_n179), .b(new_n180), .c(new_n174), .d(new_n182), .o1(\s[17] ));
  inv000aa1d42x5               g088(.a(\a[17] ), .o1(new_n184));
  nanb02aa1n12x5               g089(.a(\b[16] ), .b(new_n184), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n180), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n186));
  tech160nm_fixorc02aa1n02p5x5 g091(.a(\a[18] ), .b(\b[17] ), .out0(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n186), .c(new_n185), .out0(\s[18] ));
  and002aa1n02x5               g093(.a(new_n187), .b(new_n180), .o(new_n189));
  aoai13aa1n03x5               g094(.a(new_n189), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n190));
  oaoi03aa1n12x5               g095(.a(\a[18] ), .b(\b[17] ), .c(new_n185), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  nor002aa1d32x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nanp02aa1n04x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n190), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n02x7               g102(.a(new_n195), .b(new_n191), .c(new_n179), .d(new_n189), .o1(new_n198));
  nor042aa1n02x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanp02aa1n04x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1n02x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  aoib12aa1n02x5               g106(.a(new_n193), .b(new_n200), .c(new_n199), .out0(new_n202));
  inv030aa1n02x5               g107(.a(new_n193), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n195), .o1(new_n204));
  aoai13aa1n02x5               g109(.a(new_n203), .b(new_n204), .c(new_n190), .d(new_n192), .o1(new_n205));
  aoi022aa1n03x5               g110(.a(new_n205), .b(new_n201), .c(new_n198), .d(new_n202), .o1(\s[20] ));
  nano23aa1d15x5               g111(.a(new_n193), .b(new_n199), .c(new_n200), .d(new_n194), .out0(new_n207));
  nand23aa1n09x5               g112(.a(new_n207), .b(new_n180), .c(new_n187), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n210));
  oaoi03aa1n12x5               g115(.a(\a[20] ), .b(\b[19] ), .c(new_n203), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aob012aa1n02x5               g117(.a(new_n212), .b(new_n207), .c(new_n191), .out0(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  xnrc02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .out0(new_n215));
  aoi012aa1n02x5               g120(.a(new_n215), .b(new_n210), .c(new_n214), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n207), .o1(new_n217));
  oai112aa1n02x5               g122(.a(new_n212), .b(new_n215), .c(new_n217), .d(new_n192), .o1(new_n218));
  aoib12aa1n02x5               g123(.a(new_n216), .b(new_n210), .c(new_n218), .out0(\s[21] ));
  xnrc02aa1n12x5               g124(.a(\b[21] ), .b(\a[22] ), .out0(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  nor042aa1n03x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n220), .b(new_n222), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n222), .o1(new_n224));
  aoai13aa1n02x5               g129(.a(new_n224), .b(new_n215), .c(new_n210), .d(new_n214), .o1(new_n225));
  aboi22aa1n03x5               g130(.a(new_n216), .b(new_n223), .c(new_n225), .d(new_n221), .out0(\s[22] ));
  norp02aa1n04x5               g131(.a(new_n220), .b(new_n215), .o1(new_n227));
  norb02aa1n03x5               g132(.a(new_n227), .b(new_n208), .out0(new_n228));
  aoai13aa1n02x5               g133(.a(new_n228), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n229));
  aoai13aa1n12x5               g134(.a(new_n227), .b(new_n211), .c(new_n207), .d(new_n191), .o1(new_n230));
  oao003aa1n02x5               g135(.a(\a[22] ), .b(\b[21] ), .c(new_n224), .carry(new_n231));
  nand42aa1n03x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  xorc02aa1n12x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  aoai13aa1n04x5               g138(.a(new_n233), .b(new_n232), .c(new_n179), .d(new_n228), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n233), .o1(new_n235));
  and003aa1n02x5               g140(.a(new_n230), .b(new_n235), .c(new_n231), .o(new_n236));
  aobi12aa1n03x7               g141(.a(new_n234), .b(new_n236), .c(new_n229), .out0(\s[23] ));
  xorc02aa1n02x5               g142(.a(\a[24] ), .b(\b[23] ), .out0(new_n238));
  nor042aa1n03x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  norp02aa1n02x5               g144(.a(new_n238), .b(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n232), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n239), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n235), .c(new_n229), .d(new_n241), .o1(new_n243));
  aoi022aa1n03x5               g148(.a(new_n243), .b(new_n238), .c(new_n234), .d(new_n240), .o1(\s[24] ));
  nano32aa1n06x5               g149(.a(new_n208), .b(new_n238), .c(new_n227), .d(new_n233), .out0(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n246));
  and002aa1n02x5               g151(.a(new_n238), .b(new_n233), .o(new_n247));
  inv020aa1n02x5               g152(.a(new_n247), .o1(new_n248));
  oao003aa1n02x5               g153(.a(\a[24] ), .b(\b[23] ), .c(new_n242), .carry(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n248), .c(new_n230), .d(new_n231), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[25] ), .b(\b[24] ), .out0(new_n251));
  aoai13aa1n04x5               g156(.a(new_n251), .b(new_n250), .c(new_n179), .d(new_n245), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n251), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n249), .b(new_n253), .o1(new_n254));
  aoi012aa1n02x5               g159(.a(new_n254), .b(new_n232), .c(new_n247), .o1(new_n255));
  aobi12aa1n03x7               g160(.a(new_n252), .b(new_n255), .c(new_n246), .out0(\s[25] ));
  xorc02aa1n02x5               g161(.a(\a[26] ), .b(\b[25] ), .out0(new_n257));
  norp02aa1n02x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  norp02aa1n02x5               g163(.a(new_n257), .b(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n250), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n258), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n253), .c(new_n246), .d(new_n260), .o1(new_n262));
  aoi022aa1n03x5               g167(.a(new_n262), .b(new_n257), .c(new_n252), .d(new_n259), .o1(\s[26] ));
  and002aa1n02x5               g168(.a(new_n257), .b(new_n251), .o(new_n264));
  nano23aa1n03x7               g169(.a(new_n248), .b(new_n208), .c(new_n264), .d(new_n227), .out0(new_n265));
  aoai13aa1n12x5               g170(.a(new_n265), .b(new_n178), .c(new_n173), .d(new_n120), .o1(new_n266));
  nand02aa1d04x5               g171(.a(new_n250), .b(new_n264), .o1(new_n267));
  nanp02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .o1(new_n268));
  oai022aa1n02x5               g173(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(new_n269), .b(new_n268), .o1(new_n270));
  nand23aa1n06x5               g175(.a(new_n266), .b(new_n267), .c(new_n270), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[27] ), .b(\b[26] ), .out0(new_n272));
  aoi122aa1n02x5               g177(.a(new_n272), .b(new_n268), .c(new_n269), .d(new_n250), .e(new_n264), .o1(new_n273));
  aoi022aa1n02x5               g178(.a(new_n273), .b(new_n266), .c(new_n271), .d(new_n272), .o1(\s[27] ));
  nand42aa1n04x5               g179(.a(new_n271), .b(new_n272), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[28] ), .b(\b[27] ), .out0(new_n276));
  norp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  norp02aa1n02x5               g182(.a(new_n276), .b(new_n277), .o1(new_n278));
  aoi022aa1n06x5               g183(.a(new_n250), .b(new_n264), .c(new_n268), .d(new_n269), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n277), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n272), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n280), .b(new_n281), .c(new_n279), .d(new_n266), .o1(new_n282));
  aoi022aa1n03x5               g187(.a(new_n282), .b(new_n276), .c(new_n275), .d(new_n278), .o1(\s[28] ));
  and002aa1n02x5               g188(.a(new_n276), .b(new_n272), .o(new_n284));
  nand42aa1n02x5               g189(.a(new_n271), .b(new_n284), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[29] ), .b(\b[28] ), .out0(new_n286));
  inv000aa1d42x5               g191(.a(\a[28] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[27] ), .o1(new_n288));
  aoi112aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n289));
  aoi112aa1n02x5               g194(.a(new_n286), .b(new_n289), .c(new_n287), .d(new_n288), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n284), .o1(new_n291));
  aoi012aa1n02x5               g196(.a(new_n289), .b(new_n287), .c(new_n288), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n291), .c(new_n279), .d(new_n266), .o1(new_n293));
  aoi022aa1n03x5               g198(.a(new_n293), .b(new_n286), .c(new_n285), .d(new_n290), .o1(\s[29] ));
  nanp02aa1n02x5               g199(.a(\b[0] ), .b(\a[1] ), .o1(new_n295));
  xorb03aa1n02x5               g200(.a(new_n295), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g201(.a(new_n281), .b(new_n276), .c(new_n286), .out0(new_n297));
  nanp02aa1n03x5               g202(.a(new_n271), .b(new_n297), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .out0(new_n299));
  tech160nm_fiao0012aa1n02p5x5 g204(.a(new_n292), .b(\a[29] ), .c(\b[28] ), .o(new_n300));
  oabi12aa1n02x5               g205(.a(new_n299), .b(\a[29] ), .c(\b[28] ), .out0(new_n301));
  norb02aa1n02x5               g206(.a(new_n300), .b(new_n301), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n297), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[29] ), .b(\b[28] ), .c(new_n292), .carry(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n303), .c(new_n279), .d(new_n266), .o1(new_n305));
  aoi022aa1n03x5               g210(.a(new_n305), .b(new_n299), .c(new_n298), .d(new_n302), .o1(\s[30] ));
  nano32aa1n02x4               g211(.a(new_n281), .b(new_n299), .c(new_n276), .d(new_n286), .out0(new_n307));
  nand42aa1n02x5               g212(.a(new_n271), .b(new_n307), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[31] ), .b(\b[30] ), .out0(new_n309));
  oa0022aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(\a[29] ), .d(\b[28] ), .o(new_n310));
  ao0022aa1n03x5               g215(.a(new_n300), .b(new_n310), .c(\a[30] ), .d(\b[29] ), .o(new_n311));
  norb02aa1n02x5               g216(.a(new_n311), .b(new_n309), .out0(new_n312));
  inv000aa1n02x5               g217(.a(new_n307), .o1(new_n313));
  aoai13aa1n03x5               g218(.a(new_n311), .b(new_n313), .c(new_n279), .d(new_n266), .o1(new_n314));
  aoi022aa1n03x5               g219(.a(new_n314), .b(new_n309), .c(new_n308), .d(new_n312), .o1(\s[31] ));
  nanb02aa1n02x5               g220(.a(new_n100), .b(new_n101), .out0(new_n316));
  xnbna2aa1n03x5               g221(.a(new_n316), .b(new_n98), .c(new_n99), .out0(\s[3] ));
  inv000aa1d42x5               g222(.a(new_n103), .o1(new_n318));
  and002aa1n02x5               g223(.a(\b[3] ), .b(\a[4] ), .o(new_n319));
  norp02aa1n02x5               g224(.a(new_n319), .b(new_n102), .o1(new_n320));
  aoi113aa1n02x5               g225(.a(new_n320), .b(new_n100), .c(new_n98), .d(new_n101), .e(new_n99), .o1(new_n321));
  aoi012aa1n02x5               g226(.a(new_n321), .b(new_n318), .c(new_n320), .o1(\s[4] ));
  norb02aa1n02x5               g227(.a(new_n106), .b(new_n103), .out0(new_n323));
  xnrc02aa1n02x5               g228(.a(\b[4] ), .b(\a[5] ), .out0(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n323), .b(new_n324), .c(new_n103), .d(new_n319), .o1(\s[5] ));
  norb02aa1n02x5               g230(.a(new_n111), .b(new_n110), .out0(new_n326));
  inv000aa1n03x5               g231(.a(new_n323), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n326), .b(new_n327), .c(new_n115), .out0(\s[6] ));
  inv000aa1d42x5               g233(.a(new_n116), .o1(new_n329));
  nanb03aa1n02x5               g234(.a(new_n103), .b(new_n326), .c(new_n106), .out0(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n114), .b(new_n330), .c(new_n329), .out0(\s[7] ));
  aob012aa1n02x5               g236(.a(new_n114), .b(new_n330), .c(new_n329), .out0(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n107), .b(new_n332), .c(new_n117), .out0(\s[8] ));
  nanb02aa1n02x5               g238(.a(new_n113), .b(new_n318), .out0(new_n334));
  aoi113aa1n02x5               g239(.a(new_n121), .b(new_n118), .c(new_n116), .d(new_n107), .e(new_n114), .o1(new_n335));
  aoi022aa1n02x5               g240(.a(new_n334), .b(new_n335), .c(new_n120), .d(new_n121), .o1(\s[9] ));
endmodule


