// Benchmark "adder" written by ABC on Thu Jul 18 11:56:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n319, new_n320, new_n322, new_n323, new_n325, new_n326,
    new_n327, new_n328, new_n330, new_n332, new_n333, new_n334, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv030aa1n06x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  oab012aa1n06x5               g004(.a(new_n99), .b(\a[4] ), .c(\b[3] ), .out0(new_n100));
  nanp02aa1n02x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nanb02aa1n06x5               g006(.a(new_n99), .b(new_n101), .out0(new_n102));
  nanp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n06x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nor002aa1n03x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  oai012aa1n06x5               g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  oaih12aa1n06x5               g011(.a(new_n100), .b(new_n106), .c(new_n102), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[7] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[6] ), .o1(new_n109));
  nand02aa1n06x5               g014(.a(new_n109), .b(new_n108), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  oai112aa1n02x5               g016(.a(new_n110), .b(new_n111), .c(\b[5] ), .d(\a[6] ), .o1(new_n112));
  tech160nm_fixnrc02aa1n04x5   g017(.a(\b[4] ), .b(\a[5] ), .out0(new_n113));
  aoi022aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n114));
  inv040aa1d32x5               g019(.a(\a[8] ), .o1(new_n115));
  inv000aa1d42x5               g020(.a(\b[7] ), .o1(new_n116));
  nand42aa1n02x5               g021(.a(new_n116), .b(new_n115), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanp03aa1n02x5               g023(.a(new_n114), .b(new_n117), .c(new_n118), .o1(new_n119));
  nor043aa1n03x5               g024(.a(new_n119), .b(new_n112), .c(new_n113), .o1(new_n120));
  oai022aa1n02x5               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  nanp02aa1n03x5               g026(.a(new_n121), .b(new_n118), .o1(new_n122));
  aoi022aa1n06x5               g027(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n123));
  inv000aa1n02x5               g028(.a(new_n123), .o1(new_n124));
  aoai13aa1n06x5               g029(.a(new_n117), .b(new_n124), .c(new_n122), .d(new_n110), .o1(new_n125));
  xnrc02aa1n12x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  inv000aa1d42x5               g031(.a(new_n126), .o1(new_n127));
  aoai13aa1n03x5               g032(.a(new_n127), .b(new_n125), .c(new_n120), .d(new_n107), .o1(new_n128));
  tech160nm_fixnrc02aa1n04x5   g033(.a(\b[9] ), .b(\a[10] ), .out0(new_n129));
  xobna2aa1n03x5               g034(.a(new_n129), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  oaoi03aa1n12x5               g035(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  aoai13aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n128), .d(new_n98), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nand22aa1n06x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  norb02aa1n06x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  nor042aa1n06x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nanp02aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  aoi012aa1n03x5               g044(.a(new_n138), .b(new_n133), .c(new_n139), .o1(new_n140));
  xnrc02aa1n02x5               g045(.a(new_n140), .b(new_n137), .out0(\s[12] ));
  nona23aa1n03x5               g046(.a(new_n136), .b(new_n139), .c(new_n138), .d(new_n135), .out0(new_n142));
  norp03aa1n02x5               g047(.a(new_n142), .b(new_n129), .c(new_n126), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n125), .c(new_n120), .d(new_n107), .o1(new_n144));
  norp02aa1n02x5               g049(.a(\b[9] ), .b(\a[10] ), .o1(new_n145));
  aoi112aa1n03x5               g050(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n146));
  norb02aa1n03x4               g051(.a(new_n139), .b(new_n138), .out0(new_n147));
  oai112aa1n03x5               g052(.a(new_n147), .b(new_n137), .c(new_n146), .d(new_n145), .o1(new_n148));
  oa0012aa1n03x5               g053(.a(new_n136), .b(new_n135), .c(new_n138), .o(new_n149));
  inv040aa1n02x5               g054(.a(new_n149), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n148), .b(new_n150), .o1(new_n151));
  inv000aa1n02x5               g056(.a(new_n151), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(new_n144), .b(new_n152), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n155), .b(new_n153), .c(new_n156), .o1(new_n157));
  xnrb03aa1n02x5               g062(.a(new_n157), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nanp02aa1n04x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nona23aa1n09x5               g065(.a(new_n160), .b(new_n156), .c(new_n155), .d(new_n159), .out0(new_n161));
  oai012aa1n12x5               g066(.a(new_n160), .b(new_n159), .c(new_n155), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n161), .c(new_n144), .d(new_n152), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand02aa1n03x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  aoi012aa1n03x5               g071(.a(new_n165), .b(new_n163), .c(new_n166), .o1(new_n167));
  xnrb03aa1n03x5               g072(.a(new_n167), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  tech160nm_fiaoi012aa1n03p5x5 g073(.a(new_n125), .b(new_n120), .c(new_n107), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand22aa1n04x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nona23aa1d18x5               g076(.a(new_n171), .b(new_n166), .c(new_n165), .d(new_n170), .out0(new_n172));
  nor042aa1n06x5               g077(.a(new_n172), .b(new_n161), .o1(new_n173));
  nona32aa1n09x5               g078(.a(new_n173), .b(new_n142), .c(new_n129), .d(new_n126), .out0(new_n174));
  inv030aa1n02x5               g079(.a(new_n172), .o1(new_n175));
  aoai13aa1n06x5               g080(.a(new_n162), .b(new_n161), .c(new_n150), .d(new_n148), .o1(new_n176));
  nand42aa1n04x5               g081(.a(new_n176), .b(new_n175), .o1(new_n177));
  aoi012aa1d18x5               g082(.a(new_n170), .b(new_n165), .c(new_n171), .o1(new_n178));
  oai112aa1n06x5               g083(.a(new_n177), .b(new_n178), .c(new_n174), .d(new_n169), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g085(.a(\a[17] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\b[16] ), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(new_n182), .b(new_n181), .o1(new_n183));
  nanp02aa1n06x5               g088(.a(new_n120), .b(new_n107), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n122), .b(new_n110), .o1(new_n185));
  aoi022aa1n09x5               g090(.a(new_n185), .b(new_n123), .c(new_n116), .d(new_n115), .o1(new_n186));
  aoi012aa1d18x5               g091(.a(new_n174), .b(new_n184), .c(new_n186), .o1(new_n187));
  nano23aa1n02x4               g092(.a(new_n138), .b(new_n135), .c(new_n136), .d(new_n139), .out0(new_n188));
  inv040aa1n02x5               g093(.a(new_n161), .o1(new_n189));
  aoai13aa1n04x5               g094(.a(new_n189), .b(new_n149), .c(new_n188), .d(new_n131), .o1(new_n190));
  aoai13aa1n12x5               g095(.a(new_n178), .b(new_n172), .c(new_n190), .d(new_n162), .o1(new_n191));
  xorc02aa1n12x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  oaih12aa1n02x5               g097(.a(new_n192), .b(new_n191), .c(new_n187), .o1(new_n193));
  nor002aa1n03x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  nand22aa1n06x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nanb02aa1n09x5               g100(.a(new_n194), .b(new_n195), .out0(new_n196));
  xobna2aa1n03x5               g101(.a(new_n196), .b(new_n193), .c(new_n183), .out0(\s[18] ));
  norb02aa1n02x5               g102(.a(new_n192), .b(new_n196), .out0(new_n198));
  tech160nm_fioai012aa1n05x5   g103(.a(new_n198), .b(new_n191), .c(new_n187), .o1(new_n199));
  aoi013aa1n09x5               g104(.a(new_n194), .b(new_n195), .c(new_n181), .d(new_n182), .o1(new_n200));
  nor002aa1d32x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nand42aa1n04x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  xnbna2aa1n03x5               g108(.a(new_n203), .b(new_n199), .c(new_n200), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g110(.a(new_n199), .b(new_n200), .o1(new_n206));
  nor002aa1d32x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nand22aa1n09x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nanb02aa1n02x5               g113(.a(new_n207), .b(new_n208), .out0(new_n209));
  aoai13aa1n02x5               g114(.a(new_n209), .b(new_n201), .c(new_n206), .d(new_n203), .o1(new_n210));
  oaoi03aa1n02x5               g115(.a(\a[18] ), .b(\b[17] ), .c(new_n183), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n203), .b(new_n211), .c(new_n179), .d(new_n198), .o1(new_n212));
  nona22aa1n02x5               g117(.a(new_n212), .b(new_n209), .c(new_n201), .out0(new_n213));
  nanp02aa1n03x5               g118(.a(new_n210), .b(new_n213), .o1(\s[20] ));
  inv000aa1d42x5               g119(.a(new_n178), .o1(new_n215));
  aoi112aa1n06x5               g120(.a(new_n187), .b(new_n215), .c(new_n175), .d(new_n176), .o1(new_n216));
  nona23aa1d18x5               g121(.a(new_n208), .b(new_n202), .c(new_n201), .d(new_n207), .out0(new_n217));
  norb03aa1n06x5               g122(.a(new_n192), .b(new_n217), .c(new_n196), .out0(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  oa0012aa1n03x5               g124(.a(new_n208), .b(new_n207), .c(new_n201), .o(new_n220));
  oabi12aa1n18x5               g125(.a(new_n220), .b(new_n200), .c(new_n217), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oai012aa1n04x7               g127(.a(new_n222), .b(new_n216), .c(new_n219), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  tech160nm_fixnrc02aa1n05x5   g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  aoai13aa1n03x5               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n227), .b(new_n221), .c(new_n179), .d(new_n218), .o1(new_n230));
  nona22aa1n02x5               g135(.a(new_n230), .b(new_n228), .c(new_n225), .out0(new_n231));
  nanp02aa1n03x5               g136(.a(new_n229), .b(new_n231), .o1(\s[22] ));
  nor042aa1n09x5               g137(.a(new_n228), .b(new_n226), .o1(new_n233));
  nona23aa1d24x5               g138(.a(new_n233), .b(new_n192), .c(new_n217), .d(new_n196), .out0(new_n234));
  inv000aa1d42x5               g139(.a(\a[22] ), .o1(new_n235));
  inv000aa1d42x5               g140(.a(\b[21] ), .o1(new_n236));
  oaoi03aa1n09x5               g141(.a(new_n235), .b(new_n236), .c(new_n225), .o1(new_n237));
  inv040aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1d24x5               g143(.a(new_n238), .b(new_n221), .c(new_n233), .o1(new_n239));
  oai012aa1n06x5               g144(.a(new_n239), .b(new_n216), .c(new_n234), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  xorc02aa1n12x5               g147(.a(\a[23] ), .b(\b[22] ), .out0(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[23] ), .b(\a[24] ), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n242), .c(new_n240), .d(new_n243), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n234), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n239), .o1(new_n247));
  aoai13aa1n03x5               g152(.a(new_n243), .b(new_n247), .c(new_n179), .d(new_n246), .o1(new_n248));
  nona22aa1n02x5               g153(.a(new_n248), .b(new_n244), .c(new_n242), .out0(new_n249));
  nanp02aa1n03x5               g154(.a(new_n245), .b(new_n249), .o1(\s[24] ));
  norb02aa1n03x5               g155(.a(new_n243), .b(new_n244), .out0(new_n251));
  inv030aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  nor042aa1n04x5               g157(.a(new_n234), .b(new_n252), .o1(new_n253));
  oai012aa1n06x5               g158(.a(new_n253), .b(new_n191), .c(new_n187), .o1(new_n254));
  nano23aa1n02x5               g159(.a(new_n201), .b(new_n207), .c(new_n208), .d(new_n202), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n233), .b(new_n220), .c(new_n255), .d(new_n211), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n257));
  oab012aa1n02x4               g162(.a(new_n257), .b(\a[24] ), .c(\b[23] ), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n252), .c(new_n256), .d(new_n237), .o1(new_n259));
  inv030aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  xorc02aa1n12x5               g165(.a(\a[25] ), .b(\b[24] ), .out0(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n254), .c(new_n260), .out0(\s[25] ));
  nanp02aa1n06x5               g167(.a(new_n254), .b(new_n260), .o1(new_n263));
  norp02aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  tech160nm_fixnrc02aa1n02p5x5 g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n264), .c(new_n263), .d(new_n261), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n261), .b(new_n259), .c(new_n179), .d(new_n253), .o1(new_n267));
  nona22aa1n02x5               g172(.a(new_n267), .b(new_n265), .c(new_n264), .out0(new_n268));
  nanp02aa1n03x5               g173(.a(new_n266), .b(new_n268), .o1(\s[26] ));
  norb02aa1n06x4               g174(.a(new_n261), .b(new_n265), .out0(new_n270));
  nano22aa1n12x5               g175(.a(new_n234), .b(new_n251), .c(new_n270), .out0(new_n271));
  tech160nm_fioai012aa1n04x5   g176(.a(new_n271), .b(new_n191), .c(new_n187), .o1(new_n272));
  inv000aa1d42x5               g177(.a(\a[26] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\b[25] ), .o1(new_n274));
  tech160nm_fioaoi03aa1n03p5x5 g179(.a(new_n273), .b(new_n274), .c(new_n264), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoi012aa1n09x5               g181(.a(new_n276), .b(new_n259), .c(new_n270), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n277), .c(new_n272), .out0(\s[27] ));
  inv020aa1n03x5               g184(.a(new_n271), .o1(new_n280));
  oai012aa1n06x5               g185(.a(new_n277), .b(new_n216), .c(new_n280), .o1(new_n281));
  norp02aa1n02x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  norp02aa1n04x5               g187(.a(\b[27] ), .b(\a[28] ), .o1(new_n283));
  nanp02aa1n04x5               g188(.a(\b[27] ), .b(\a[28] ), .o1(new_n284));
  nanb02aa1n06x5               g189(.a(new_n283), .b(new_n284), .out0(new_n285));
  aoai13aa1n04x5               g190(.a(new_n285), .b(new_n282), .c(new_n281), .d(new_n278), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n251), .b(new_n238), .c(new_n221), .d(new_n233), .o1(new_n287));
  inv000aa1n02x5               g192(.a(new_n270), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n275), .b(new_n288), .c(new_n287), .d(new_n258), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n278), .b(new_n289), .c(new_n179), .d(new_n271), .o1(new_n290));
  nona22aa1n02x5               g195(.a(new_n290), .b(new_n285), .c(new_n282), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n286), .b(new_n291), .o1(\s[28] ));
  norb02aa1n03x5               g197(.a(new_n278), .b(new_n285), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n179), .d(new_n271), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n293), .o1(new_n295));
  oai012aa1n02x5               g200(.a(new_n284), .b(new_n283), .c(new_n282), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n295), .c(new_n277), .d(new_n272), .o1(new_n297));
  xorc02aa1n12x5               g202(.a(\a[29] ), .b(\b[28] ), .out0(new_n298));
  norb02aa1n02x5               g203(.a(new_n296), .b(new_n298), .out0(new_n299));
  aoi022aa1n02x7               g204(.a(new_n297), .b(new_n298), .c(new_n294), .d(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g206(.a(new_n285), .b(new_n278), .c(new_n298), .out0(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n289), .c(new_n179), .d(new_n271), .o1(new_n303));
  inv000aa1n02x5               g208(.a(new_n302), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n305));
  aoai13aa1n02x7               g210(.a(new_n305), .b(new_n304), .c(new_n277), .d(new_n272), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[30] ));
  nand03aa1n02x5               g214(.a(new_n293), .b(new_n298), .c(new_n307), .o1(new_n310));
  nanb02aa1n03x5               g215(.a(new_n310), .b(new_n281), .out0(new_n311));
  oao003aa1n02x5               g216(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n312));
  aoai13aa1n02x7               g217(.a(new_n312), .b(new_n310), .c(new_n277), .d(new_n272), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[31] ), .b(\b[30] ), .out0(new_n314));
  norb02aa1n02x5               g219(.a(new_n312), .b(new_n314), .out0(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n311), .d(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g221(.a(new_n106), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  orn002aa1n02x5               g222(.a(new_n106), .b(new_n102), .o(new_n318));
  xorc02aa1n02x5               g223(.a(\a[4] ), .b(\b[3] ), .out0(new_n319));
  norp02aa1n02x5               g224(.a(new_n319), .b(new_n99), .o1(new_n320));
  aoi022aa1n02x5               g225(.a(new_n318), .b(new_n320), .c(new_n107), .d(new_n319), .o1(\s[4] ));
  and002aa1n02x5               g226(.a(\b[3] ), .b(\a[4] ), .o(new_n322));
  inv000aa1d42x5               g227(.a(new_n322), .o1(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n113), .b(new_n107), .c(new_n323), .out0(\s[5] ));
  nona22aa1n02x4               g229(.a(new_n107), .b(new_n113), .c(new_n322), .out0(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[5] ), .b(\a[6] ), .out0(new_n326));
  oaoi13aa1n02x5               g231(.a(new_n326), .b(new_n325), .c(\a[5] ), .d(\b[4] ), .o1(new_n327));
  oai112aa1n02x5               g232(.a(new_n325), .b(new_n326), .c(\b[4] ), .d(\a[5] ), .o1(new_n328));
  norb02aa1n02x5               g233(.a(new_n328), .b(new_n327), .out0(\s[6] ));
  nanb02aa1n02x5               g234(.a(new_n327), .b(new_n122), .out0(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp03aa1n02x5               g236(.a(new_n330), .b(new_n110), .c(new_n111), .o1(new_n332));
  aob012aa1n02x5               g237(.a(new_n110), .b(new_n330), .c(new_n111), .out0(new_n333));
  xorc02aa1n02x5               g238(.a(\a[8] ), .b(\b[7] ), .out0(new_n334));
  norb02aa1n02x5               g239(.a(new_n110), .b(new_n334), .out0(new_n335));
  aoi022aa1n02x5               g240(.a(new_n333), .b(new_n334), .c(new_n332), .d(new_n335), .o1(\s[8] ));
  xnbna2aa1n03x5               g241(.a(new_n127), .b(new_n184), .c(new_n186), .out0(\s[9] ));
endmodule


