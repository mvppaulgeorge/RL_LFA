// Benchmark "adder" written by ABC on Thu Jul 18 08:49:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n306, new_n307, new_n308, new_n311, new_n313,
    new_n315;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  nor002aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n03x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor002aa1d32x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1n08x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n02x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor002aa1n12x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n02x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nanb03aa1n03x5               g013(.a(new_n102), .b(new_n108), .c(new_n105), .out0(new_n109));
  tech160nm_fiaoi012aa1n03p5x5 g014(.a(new_n103), .b(new_n106), .c(new_n104), .o1(new_n110));
  nor042aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand02aa1n04x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1n10x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand22aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nano23aa1n03x7               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nona22aa1n02x4               g022(.a(new_n115), .b(new_n116), .c(new_n117), .out0(new_n118));
  inv040aa1d32x5               g023(.a(\a[5] ), .o1(new_n119));
  inv040aa1d28x5               g024(.a(\b[4] ), .o1(new_n120));
  tech160nm_finand02aa1n03p5x5 g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  tech160nm_fiaoi012aa1n03p5x5 g027(.a(new_n111), .b(new_n113), .c(new_n112), .o1(new_n123));
  aobi12aa1n06x5               g028(.a(new_n123), .b(new_n115), .c(new_n122), .out0(new_n124));
  aoai13aa1n04x5               g029(.a(new_n124), .b(new_n118), .c(new_n109), .d(new_n110), .o1(new_n125));
  tech160nm_fixorc02aa1n03p5x5 g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoi012aa1n02x5               g031(.a(new_n98), .b(new_n125), .c(new_n126), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  tech160nm_fixorc02aa1n02p5x5 g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  inv000aa1d42x5               g034(.a(\b[9] ), .o1(new_n130));
  oao003aa1n02x5               g035(.a(new_n97), .b(new_n130), .c(new_n98), .carry(new_n131));
  aoi013aa1n03x5               g036(.a(new_n131), .b(new_n125), .c(new_n126), .d(new_n129), .o1(new_n132));
  xnrb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  oaoi03aa1n02x5               g038(.a(\a[11] ), .b(\b[10] ), .c(new_n132), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nona23aa1n09x5               g040(.a(new_n107), .b(new_n104), .c(new_n103), .d(new_n106), .out0(new_n136));
  oaih12aa1n06x5               g041(.a(new_n110), .b(new_n136), .c(new_n102), .o1(new_n137));
  nona23aa1n09x5               g042(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n138));
  nor043aa1n03x5               g043(.a(new_n138), .b(new_n116), .c(new_n117), .o1(new_n139));
  oaib12aa1n06x5               g044(.a(new_n123), .b(new_n138), .c(new_n122), .out0(new_n140));
  nor022aa1n16x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  tech160nm_finand02aa1n03p5x5 g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n04x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nona23aa1n02x4               g049(.a(new_n144), .b(new_n142), .c(new_n141), .d(new_n143), .out0(new_n145));
  nano22aa1n02x4               g050(.a(new_n145), .b(new_n129), .c(new_n126), .out0(new_n146));
  aoai13aa1n06x5               g051(.a(new_n146), .b(new_n140), .c(new_n137), .d(new_n139), .o1(new_n147));
  nano23aa1n03x7               g052(.a(new_n141), .b(new_n143), .c(new_n144), .d(new_n142), .out0(new_n148));
  tech160nm_fiaoi012aa1n03p5x5 g053(.a(new_n143), .b(new_n141), .c(new_n144), .o1(new_n149));
  aobi12aa1n06x5               g054(.a(new_n149), .b(new_n148), .c(new_n131), .out0(new_n150));
  xorc02aa1n12x5               g055(.a(\a[13] ), .b(\b[12] ), .out0(new_n151));
  xnbna2aa1n03x5               g056(.a(new_n151), .b(new_n147), .c(new_n150), .out0(\s[13] ));
  orn002aa1n24x5               g057(.a(\a[13] ), .b(\b[12] ), .o(new_n153));
  oaoi03aa1n02x5               g058(.a(new_n97), .b(new_n130), .c(new_n98), .o1(new_n154));
  oaih12aa1n06x5               g059(.a(new_n149), .b(new_n145), .c(new_n154), .o1(new_n155));
  aoai13aa1n02x5               g060(.a(new_n151), .b(new_n155), .c(new_n125), .d(new_n146), .o1(new_n156));
  xorc02aa1n12x5               g061(.a(\a[14] ), .b(\b[13] ), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n156), .c(new_n153), .out0(\s[14] ));
  nanp02aa1n02x5               g063(.a(new_n157), .b(new_n151), .o1(new_n159));
  oaoi03aa1n12x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n153), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n04x5               g066(.a(new_n161), .b(new_n159), .c(new_n147), .d(new_n150), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand02aa1d24x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  norp02aa1n06x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand02aa1d16x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n164), .b(new_n168), .c(new_n162), .d(new_n165), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nano23aa1n06x5               g076(.a(new_n164), .b(new_n166), .c(new_n167), .d(new_n165), .out0(new_n172));
  nand23aa1n02x5               g077(.a(new_n172), .b(new_n151), .c(new_n157), .o1(new_n173));
  nano32aa1n03x7               g078(.a(new_n173), .b(new_n148), .c(new_n126), .d(new_n129), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n140), .c(new_n137), .d(new_n139), .o1(new_n175));
  tech160nm_fiao0012aa1n02p5x5 g080(.a(new_n166), .b(new_n164), .c(new_n167), .o(new_n176));
  tech160nm_fiao0012aa1n03p5x5 g081(.a(new_n176), .b(new_n172), .c(new_n160), .o(new_n177));
  aoib12aa1n12x5               g082(.a(new_n177), .b(new_n155), .c(new_n173), .out0(new_n178));
  nanp02aa1n09x5               g083(.a(new_n175), .b(new_n178), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  xroi22aa1d06x4               g090(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n186));
  oai022aa1d24x5               g091(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n187));
  oaib12aa1n18x5               g092(.a(new_n187), .b(new_n181), .c(\b[17] ), .out0(new_n188));
  inv040aa1n08x5               g093(.a(new_n188), .o1(new_n189));
  aoi012aa1n09x5               g094(.a(new_n189), .b(new_n179), .c(new_n186), .o1(new_n190));
  nor002aa1d32x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  nand02aa1n08x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n190), .b(new_n193), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g100(.a(new_n191), .b(new_n193), .out0(new_n196));
  nor042aa1n06x5               g101(.a(\b[19] ), .b(\a[20] ), .o1(new_n197));
  nand02aa1d16x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nanb02aa1n02x5               g103(.a(new_n197), .b(new_n198), .out0(new_n199));
  oaoi13aa1n02x7               g104(.a(new_n199), .b(new_n192), .c(new_n190), .d(new_n196), .o1(new_n200));
  nor042aa1n02x5               g105(.a(new_n190), .b(new_n196), .o1(new_n201));
  nano22aa1n03x7               g106(.a(new_n201), .b(new_n192), .c(new_n199), .out0(new_n202));
  norp02aa1n03x5               g107(.a(new_n200), .b(new_n202), .o1(\s[20] ));
  nano23aa1n09x5               g108(.a(new_n191), .b(new_n197), .c(new_n198), .d(new_n193), .out0(new_n204));
  nanp02aa1n02x5               g109(.a(new_n186), .b(new_n204), .o1(new_n205));
  nona23aa1n09x5               g110(.a(new_n198), .b(new_n193), .c(new_n191), .d(new_n197), .out0(new_n206));
  aoi012aa1n09x5               g111(.a(new_n197), .b(new_n191), .c(new_n198), .o1(new_n207));
  oai012aa1n18x5               g112(.a(new_n207), .b(new_n206), .c(new_n188), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n205), .c(new_n175), .d(new_n178), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g116(.a(\b[20] ), .b(\a[21] ), .o1(new_n212));
  xorc02aa1n02x5               g117(.a(\a[21] ), .b(\b[20] ), .out0(new_n213));
  xorc02aa1n02x5               g118(.a(\a[22] ), .b(\b[21] ), .out0(new_n214));
  aoai13aa1n03x5               g119(.a(new_n214), .b(new_n212), .c(new_n210), .d(new_n213), .o1(new_n215));
  aoi112aa1n02x5               g120(.a(new_n212), .b(new_n214), .c(new_n210), .d(new_n213), .o1(new_n216));
  norb02aa1n03x4               g121(.a(new_n215), .b(new_n216), .out0(\s[22] ));
  inv000aa1d42x5               g122(.a(\a[21] ), .o1(new_n218));
  inv040aa1d32x5               g123(.a(\a[22] ), .o1(new_n219));
  xroi22aa1d06x4               g124(.a(new_n218), .b(\b[20] ), .c(new_n219), .d(\b[21] ), .out0(new_n220));
  nand03aa1n02x5               g125(.a(new_n220), .b(new_n186), .c(new_n204), .o1(new_n221));
  inv000aa1d42x5               g126(.a(\b[21] ), .o1(new_n222));
  oao003aa1n02x5               g127(.a(new_n219), .b(new_n222), .c(new_n212), .carry(new_n223));
  aoi012aa1n02x5               g128(.a(new_n223), .b(new_n208), .c(new_n220), .o1(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n221), .c(new_n175), .d(new_n178), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g131(.a(\b[22] ), .b(\a[23] ), .o1(new_n227));
  xorc02aa1n12x5               g132(.a(\a[23] ), .b(\b[22] ), .out0(new_n228));
  tech160nm_fixorc02aa1n05x5   g133(.a(\a[24] ), .b(\b[23] ), .out0(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n227), .c(new_n225), .d(new_n228), .o1(new_n230));
  aoi112aa1n03x5               g135(.a(new_n227), .b(new_n229), .c(new_n225), .d(new_n228), .o1(new_n231));
  norb02aa1n03x4               g136(.a(new_n230), .b(new_n231), .out0(\s[24] ));
  aoi012aa1n02x5               g137(.a(new_n176), .b(new_n172), .c(new_n160), .o1(new_n233));
  oaih12aa1n02x5               g138(.a(new_n233), .b(new_n150), .c(new_n173), .o1(new_n234));
  and002aa1n03x5               g139(.a(new_n229), .b(new_n228), .o(new_n235));
  inv000aa1n03x5               g140(.a(new_n235), .o1(new_n236));
  nano32aa1n03x7               g141(.a(new_n236), .b(new_n220), .c(new_n186), .d(new_n204), .out0(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n125), .d(new_n174), .o1(new_n238));
  inv020aa1n03x5               g143(.a(new_n207), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n220), .b(new_n239), .c(new_n204), .d(new_n189), .o1(new_n240));
  inv000aa1n02x5               g145(.a(new_n223), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n242));
  oab012aa1n02x4               g147(.a(new_n242), .b(\a[24] ), .c(\b[23] ), .out0(new_n243));
  aoai13aa1n12x5               g148(.a(new_n243), .b(new_n236), .c(new_n240), .d(new_n241), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[24] ), .b(\a[25] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xnbna2aa1n03x5               g152(.a(new_n247), .b(new_n238), .c(new_n245), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n247), .b(new_n244), .c(new_n179), .d(new_n237), .o1(new_n251));
  xnrc02aa1n12x5               g156(.a(\b[25] ), .b(\a[26] ), .out0(new_n252));
  aoi012aa1n02x7               g157(.a(new_n252), .b(new_n251), .c(new_n250), .o1(new_n253));
  nand23aa1n03x5               g158(.a(new_n251), .b(new_n250), .c(new_n252), .o1(new_n254));
  norb02aa1n02x7               g159(.a(new_n254), .b(new_n253), .out0(\s[26] ));
  nor042aa1n06x5               g160(.a(new_n252), .b(new_n246), .o1(new_n256));
  nano22aa1n06x5               g161(.a(new_n221), .b(new_n235), .c(new_n256), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n234), .c(new_n125), .d(new_n174), .o1(new_n258));
  nanp02aa1n09x5               g163(.a(new_n244), .b(new_n256), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .c(new_n250), .carry(new_n260));
  xorc02aa1n12x5               g165(.a(\a[27] ), .b(\b[26] ), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoi013aa1n06x4               g167(.a(new_n262), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n263));
  aobi12aa1n06x5               g168(.a(new_n257), .b(new_n175), .c(new_n178), .out0(new_n264));
  aoai13aa1n03x5               g169(.a(new_n235), .b(new_n223), .c(new_n208), .d(new_n220), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n256), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n260), .b(new_n266), .c(new_n265), .d(new_n243), .o1(new_n267));
  norp03aa1n02x5               g172(.a(new_n267), .b(new_n264), .c(new_n261), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n263), .b(new_n268), .o1(\s[27] ));
  nor042aa1n03x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  oaih12aa1n02x5               g176(.a(new_n261), .b(new_n267), .c(new_n264), .o1(new_n272));
  xnrc02aa1n12x5               g177(.a(\b[27] ), .b(\a[28] ), .out0(new_n273));
  aoi012aa1n03x5               g178(.a(new_n273), .b(new_n272), .c(new_n271), .o1(new_n274));
  nano22aa1n03x5               g179(.a(new_n263), .b(new_n271), .c(new_n273), .out0(new_n275));
  norp02aa1n03x5               g180(.a(new_n274), .b(new_n275), .o1(\s[28] ));
  norb02aa1n02x5               g181(.a(new_n261), .b(new_n273), .out0(new_n277));
  tech160nm_fioai012aa1n03p5x5 g182(.a(new_n277), .b(new_n267), .c(new_n264), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[28] ), .b(\b[27] ), .c(new_n271), .carry(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[28] ), .b(\a[29] ), .out0(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n278), .c(new_n279), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n277), .o1(new_n282));
  aoi013aa1n03x5               g187(.a(new_n282), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n283));
  nano22aa1n03x5               g188(.a(new_n283), .b(new_n279), .c(new_n280), .out0(new_n284));
  norp02aa1n03x5               g189(.a(new_n281), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g190(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g191(.a(new_n261), .b(new_n280), .c(new_n273), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n267), .c(new_n264), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n279), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  aoi012aa1n03x5               g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n287), .o1(new_n292));
  aoi013aa1n03x5               g197(.a(new_n292), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n290), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n291), .b(new_n294), .o1(\s[30] ));
  norb02aa1n02x5               g200(.a(new_n287), .b(new_n290), .out0(new_n296));
  inv000aa1n02x5               g201(.a(new_n296), .o1(new_n297));
  aoi013aa1n03x5               g202(.a(new_n297), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n300), .out0(new_n301));
  oaih12aa1n02x5               g206(.a(new_n296), .b(new_n267), .c(new_n264), .o1(new_n302));
  aoi012aa1n03x5               g207(.a(new_n300), .b(new_n302), .c(new_n299), .o1(new_n303));
  norp02aa1n03x5               g208(.a(new_n303), .b(new_n301), .o1(\s[31] ));
  xnrb03aa1n02x5               g209(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g210(.a(new_n103), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n108), .b(new_n99), .c(new_n101), .d(new_n100), .o1(new_n307));
  aoi012aa1n02x5               g212(.a(new_n106), .b(new_n306), .c(new_n104), .o1(new_n308));
  aoi022aa1n02x5               g213(.a(new_n137), .b(new_n306), .c(new_n307), .d(new_n308), .o1(\s[4] ));
  xorb03aa1n02x5               g214(.a(new_n137), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g215(.a(new_n119), .b(new_n120), .c(new_n137), .o1(new_n311));
  xnrb03aa1n02x5               g216(.a(new_n311), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g217(.a(\a[6] ), .b(\b[5] ), .c(new_n311), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g219(.a(new_n113), .b(new_n313), .c(new_n114), .o1(new_n315));
  xnrb03aa1n02x5               g220(.a(new_n315), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g221(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


