// Benchmark "adder" written by ABC on Wed Jul 17 19:25:46 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n162, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n363, new_n364, new_n366, new_n367,
    new_n368, new_n369, new_n371, new_n373, new_n374, new_n375, new_n377;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[2] ), .b(\b[1] ), .o(new_n97));
  nand02aa1n08x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  aob012aa1d18x5               g003(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(new_n99));
  norp02aa1n24x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1n08x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nanb02aa1n06x5               g006(.a(new_n100), .b(new_n101), .out0(new_n102));
  nand42aa1d28x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb03aa1n06x5               g009(.a(new_n103), .b(new_n100), .c(new_n104), .out0(new_n105));
  aoai13aa1n12x5               g010(.a(new_n105), .b(new_n102), .c(new_n97), .d(new_n99), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nor043aa1n09x5               g014(.a(new_n109), .b(new_n108), .c(new_n107), .o1(new_n110));
  tech160nm_fioai012aa1n04x5   g015(.a(new_n103), .b(\b[7] ), .c(\a[8] ), .o1(new_n111));
  nand42aa1n16x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  aob012aa1d18x5               g017(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .out0(new_n113));
  aoi022aa1d24x5               g018(.a(\b[7] ), .b(\a[8] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n114));
  norb03aa1n03x5               g019(.a(new_n114), .b(new_n113), .c(new_n111), .out0(new_n115));
  inv000aa1d42x5               g020(.a(new_n108), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[7] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\b[6] ), .o1(new_n118));
  nor022aa1n08x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nand42aa1n16x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  aoai13aa1n09x5               g025(.a(new_n120), .b(new_n119), .c(new_n117), .d(new_n118), .o1(new_n121));
  norb02aa1n02x7               g026(.a(new_n112), .b(new_n109), .out0(new_n122));
  aoi022aa1d24x5               g027(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n123));
  nona23aa1n03x5               g028(.a(new_n123), .b(new_n120), .c(new_n119), .d(new_n107), .out0(new_n124));
  aoai13aa1n03x5               g029(.a(new_n121), .b(new_n124), .c(new_n122), .d(new_n116), .o1(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n106), .c(new_n110), .d(new_n115), .o1(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[9] ), .b(\b[8] ), .c(new_n126), .o1(new_n127));
  nor042aa1n09x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  and002aa1n12x5               g033(.a(\b[9] ), .b(\a[10] ), .o(new_n129));
  nor042aa1n06x5               g034(.a(new_n129), .b(new_n128), .o1(new_n130));
  norp02aa1n24x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nand02aa1n08x5               g036(.a(new_n99), .b(new_n97), .o1(new_n132));
  norb02aa1n06x5               g037(.a(new_n101), .b(new_n100), .out0(new_n133));
  nona22aa1n03x5               g038(.a(new_n103), .b(new_n104), .c(new_n100), .out0(new_n134));
  aoi012aa1n12x5               g039(.a(new_n134), .b(new_n132), .c(new_n133), .o1(new_n135));
  nona23aa1d18x5               g040(.a(new_n110), .b(new_n114), .c(new_n113), .d(new_n111), .out0(new_n136));
  inv000aa1n02x5               g041(.a(new_n121), .o1(new_n137));
  inv040aa1n03x5               g042(.a(new_n109), .o1(new_n138));
  oai112aa1n06x5               g043(.a(new_n138), .b(new_n112), .c(\b[4] ), .d(\a[5] ), .o1(new_n139));
  nor002aa1n04x5               g044(.a(new_n113), .b(new_n107), .o1(new_n140));
  norb02aa1n06x4               g045(.a(new_n120), .b(new_n119), .out0(new_n141));
  aoi013aa1n06x4               g046(.a(new_n137), .b(new_n140), .c(new_n139), .d(new_n141), .o1(new_n142));
  oai012aa1d24x5               g047(.a(new_n142), .b(new_n135), .c(new_n136), .o1(new_n143));
  xorc02aa1n12x5               g048(.a(\a[9] ), .b(\b[8] ), .out0(new_n144));
  aoi112aa1n02x5               g049(.a(new_n130), .b(new_n131), .c(new_n143), .d(new_n144), .o1(new_n145));
  aoi012aa1n02x5               g050(.a(new_n145), .b(new_n127), .c(new_n130), .o1(\s[10] ));
  aoai13aa1n06x5               g051(.a(new_n130), .b(new_n131), .c(new_n143), .d(new_n144), .o1(new_n147));
  oabi12aa1n18x5               g052(.a(new_n129), .b(new_n131), .c(new_n128), .out0(new_n148));
  nor002aa1d32x5               g053(.a(\b[10] ), .b(\a[11] ), .o1(new_n149));
  nand02aa1d28x5               g054(.a(\b[10] ), .b(\a[11] ), .o1(new_n150));
  nanb02aa1n02x5               g055(.a(new_n149), .b(new_n150), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n147), .c(new_n148), .out0(\s[11] ));
  oab012aa1n06x5               g058(.a(new_n129), .b(new_n131), .c(new_n128), .out0(new_n154));
  aoai13aa1n02x5               g059(.a(new_n152), .b(new_n154), .c(new_n127), .d(new_n130), .o1(new_n155));
  inv040aa1n02x5               g060(.a(new_n149), .o1(new_n156));
  aoai13aa1n03x5               g061(.a(new_n156), .b(new_n151), .c(new_n147), .d(new_n148), .o1(new_n157));
  nor022aa1n12x5               g062(.a(\b[11] ), .b(\a[12] ), .o1(new_n158));
  nand42aa1n10x5               g063(.a(\b[11] ), .b(\a[12] ), .o1(new_n159));
  nanb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoib12aa1n02x5               g066(.a(new_n149), .b(new_n159), .c(new_n158), .out0(new_n162));
  aoi022aa1n03x5               g067(.a(new_n157), .b(new_n161), .c(new_n155), .d(new_n162), .o1(\s[12] ));
  nano23aa1n09x5               g068(.a(new_n149), .b(new_n158), .c(new_n159), .d(new_n150), .out0(new_n164));
  nand23aa1n03x5               g069(.a(new_n164), .b(new_n144), .c(new_n130), .o1(new_n165));
  oaoi03aa1n12x5               g070(.a(\a[12] ), .b(\b[11] ), .c(new_n156), .o1(new_n166));
  tech160nm_fiaoi012aa1n05x5   g071(.a(new_n166), .b(new_n164), .c(new_n154), .o1(new_n167));
  tech160nm_fioai012aa1n02p5x5 g072(.a(new_n167), .b(new_n126), .c(new_n165), .o1(new_n168));
  nor002aa1n20x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nand02aa1d24x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  norb02aa1n03x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  nona23aa1d18x5               g076(.a(new_n159), .b(new_n150), .c(new_n149), .d(new_n158), .out0(new_n172));
  nano22aa1n03x7               g077(.a(new_n172), .b(new_n144), .c(new_n130), .out0(new_n173));
  oabi12aa1n18x5               g078(.a(new_n166), .b(new_n172), .c(new_n148), .out0(new_n174));
  aoi112aa1n02x5               g079(.a(new_n171), .b(new_n174), .c(new_n143), .d(new_n173), .o1(new_n175));
  aoi012aa1n02x5               g080(.a(new_n175), .b(new_n168), .c(new_n171), .o1(\s[13] ));
  inv000aa1d42x5               g081(.a(new_n169), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n171), .b(new_n174), .c(new_n143), .d(new_n173), .o1(new_n178));
  nor002aa1n03x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nand02aa1d12x5               g084(.a(\b[13] ), .b(\a[14] ), .o1(new_n180));
  norb02aa1n03x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n178), .c(new_n177), .out0(\s[14] ));
  nano23aa1n06x5               g087(.a(new_n169), .b(new_n179), .c(new_n180), .d(new_n170), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n174), .c(new_n143), .d(new_n173), .o1(new_n184));
  tech160nm_fioaoi03aa1n03p5x5 g089(.a(\a[14] ), .b(\b[13] ), .c(new_n177), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  xorc02aa1n12x5               g091(.a(\a[15] ), .b(\b[14] ), .out0(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n184), .c(new_n186), .out0(\s[15] ));
  aoai13aa1n02x5               g093(.a(new_n187), .b(new_n185), .c(new_n168), .d(new_n183), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[15] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[14] ), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(new_n191), .b(new_n190), .o1(new_n192));
  inv030aa1n02x5               g097(.a(new_n187), .o1(new_n193));
  aoai13aa1n02x7               g098(.a(new_n192), .b(new_n193), .c(new_n184), .d(new_n186), .o1(new_n194));
  xorc02aa1n12x5               g099(.a(\a[16] ), .b(\b[15] ), .out0(new_n195));
  inv000aa1d42x5               g100(.a(\a[16] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[15] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  and002aa1n02x5               g103(.a(\b[15] ), .b(\a[16] ), .o(new_n199));
  aboi22aa1n03x5               g104(.a(new_n199), .b(new_n198), .c(new_n191), .d(new_n190), .out0(new_n200));
  aoi022aa1n02x5               g105(.a(new_n194), .b(new_n195), .c(new_n189), .d(new_n200), .o1(\s[16] ));
  nand23aa1n03x5               g106(.a(new_n183), .b(new_n187), .c(new_n195), .o1(new_n202));
  nor042aa1n04x5               g107(.a(new_n202), .b(new_n165), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n143), .b(new_n203), .o1(new_n204));
  nano32aa1n03x7               g109(.a(new_n193), .b(new_n195), .c(new_n171), .d(new_n181), .out0(new_n205));
  nand02aa1n02x5               g110(.a(new_n205), .b(new_n173), .o1(new_n206));
  oai022aa1n03x5               g111(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(\b[14] ), .b(\a[15] ), .o1(new_n208));
  nanp03aa1n03x5               g113(.a(new_n207), .b(new_n180), .c(new_n208), .o1(new_n209));
  aoai13aa1n02x5               g114(.a(new_n198), .b(new_n199), .c(new_n209), .d(new_n192), .o1(new_n210));
  aoi012aa1n06x5               g115(.a(new_n210), .b(new_n205), .c(new_n174), .o1(new_n211));
  oai012aa1n12x5               g116(.a(new_n211), .b(new_n126), .c(new_n206), .o1(new_n212));
  xorc02aa1n02x5               g117(.a(\a[17] ), .b(\b[16] ), .out0(new_n213));
  aoi112aa1n02x5               g118(.a(new_n210), .b(new_n213), .c(new_n205), .d(new_n174), .o1(new_n214));
  aoi022aa1n02x5               g119(.a(new_n212), .b(new_n213), .c(new_n204), .d(new_n214), .o1(\s[17] ));
  inv040aa1d32x5               g120(.a(\a[17] ), .o1(new_n216));
  inv000aa1d42x5               g121(.a(\b[16] ), .o1(new_n217));
  nand02aa1d08x5               g122(.a(new_n217), .b(new_n216), .o1(new_n218));
  nanp02aa1n02x5               g123(.a(new_n209), .b(new_n192), .o1(new_n219));
  tech160nm_fioaoi03aa1n02p5x5 g124(.a(new_n196), .b(new_n197), .c(new_n219), .o1(new_n220));
  oai012aa1n12x5               g125(.a(new_n220), .b(new_n167), .c(new_n202), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n213), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[18] ), .b(\b[17] ), .out0(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n222), .c(new_n218), .out0(\s[18] ));
  inv040aa1d32x5               g129(.a(\a[18] ), .o1(new_n225));
  xroi22aa1d06x4               g130(.a(new_n216), .b(\b[16] ), .c(new_n225), .d(\b[17] ), .out0(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n227));
  oaoi03aa1n12x5               g132(.a(\a[18] ), .b(\b[17] ), .c(new_n218), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  nor002aa1d32x5               g134(.a(\b[18] ), .b(\a[19] ), .o1(new_n230));
  nand42aa1n06x5               g135(.a(\b[18] ), .b(\a[19] ), .o1(new_n231));
  norb02aa1n09x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  xnbna2aa1n03x5               g137(.a(new_n232), .b(new_n227), .c(new_n229), .out0(\s[19] ));
  xnrc02aa1n02x5               g138(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g139(.a(new_n232), .b(new_n228), .c(new_n212), .d(new_n226), .o1(new_n235));
  inv040aa1n02x5               g140(.a(new_n230), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n232), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n237), .c(new_n227), .d(new_n229), .o1(new_n238));
  xorc02aa1n02x5               g143(.a(\a[20] ), .b(\b[19] ), .out0(new_n239));
  inv040aa1d32x5               g144(.a(\a[20] ), .o1(new_n240));
  inv040aa1d28x5               g145(.a(\b[19] ), .o1(new_n241));
  nand42aa1n08x5               g146(.a(new_n241), .b(new_n240), .o1(new_n242));
  nand02aa1d16x5               g147(.a(\b[19] ), .b(\a[20] ), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n230), .b(new_n242), .c(new_n243), .o1(new_n244));
  aoi022aa1n03x5               g149(.a(new_n238), .b(new_n239), .c(new_n235), .d(new_n244), .o1(\s[20] ));
  nano32aa1n03x7               g150(.a(new_n237), .b(new_n239), .c(new_n213), .d(new_n223), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n247));
  nanp03aa1n06x5               g152(.a(new_n242), .b(new_n231), .c(new_n243), .o1(new_n248));
  nand42aa1n02x5               g153(.a(\b[17] ), .b(\a[18] ), .o1(new_n249));
  oai022aa1d18x5               g154(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n250));
  oai112aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(\b[18] ), .d(\a[19] ), .o1(new_n251));
  oaoi03aa1n12x5               g156(.a(new_n240), .b(new_n241), .c(new_n230), .o1(new_n252));
  oaih12aa1n12x5               g157(.a(new_n252), .b(new_n251), .c(new_n248), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  nor002aa1d24x5               g159(.a(\b[20] ), .b(\a[21] ), .o1(new_n255));
  nand42aa1n16x5               g160(.a(\b[20] ), .b(\a[21] ), .o1(new_n256));
  norb02aa1n02x7               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  xnbna2aa1n03x5               g162(.a(new_n257), .b(new_n247), .c(new_n254), .out0(\s[21] ));
  aoai13aa1n03x5               g163(.a(new_n257), .b(new_n253), .c(new_n212), .d(new_n246), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n255), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n257), .o1(new_n261));
  aoai13aa1n02x7               g166(.a(new_n260), .b(new_n261), .c(new_n247), .d(new_n254), .o1(new_n262));
  nor042aa1n04x5               g167(.a(\b[21] ), .b(\a[22] ), .o1(new_n263));
  nand42aa1n20x5               g168(.a(\b[21] ), .b(\a[22] ), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n264), .b(new_n263), .out0(new_n265));
  aoib12aa1n02x5               g170(.a(new_n255), .b(new_n264), .c(new_n263), .out0(new_n266));
  aoi022aa1n02x7               g171(.a(new_n262), .b(new_n265), .c(new_n259), .d(new_n266), .o1(\s[22] ));
  inv000aa1d42x5               g172(.a(new_n243), .o1(new_n268));
  nano32aa1n02x5               g173(.a(new_n268), .b(new_n236), .c(new_n242), .d(new_n231), .out0(new_n269));
  nano23aa1d15x5               g174(.a(new_n255), .b(new_n263), .c(new_n264), .d(new_n256), .out0(new_n270));
  and003aa1n03x5               g175(.a(new_n226), .b(new_n270), .c(new_n269), .o(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n272));
  oai012aa1n02x5               g177(.a(new_n264), .b(new_n263), .c(new_n255), .o1(new_n273));
  aobi12aa1n06x5               g178(.a(new_n273), .b(new_n253), .c(new_n270), .out0(new_n274));
  inv040aa1d32x5               g179(.a(\a[23] ), .o1(new_n275));
  inv040aa1d28x5               g180(.a(\b[22] ), .o1(new_n276));
  nand22aa1n12x5               g181(.a(new_n276), .b(new_n275), .o1(new_n277));
  nand22aa1n09x5               g182(.a(\b[22] ), .b(\a[23] ), .o1(new_n278));
  nand22aa1n09x5               g183(.a(new_n277), .b(new_n278), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  xnbna2aa1n03x5               g185(.a(new_n280), .b(new_n272), .c(new_n274), .out0(\s[23] ));
  inv000aa1n02x5               g186(.a(new_n274), .o1(new_n282));
  aoai13aa1n03x5               g187(.a(new_n280), .b(new_n282), .c(new_n212), .d(new_n271), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n277), .b(new_n279), .c(new_n272), .d(new_n274), .o1(new_n284));
  nor002aa1n20x5               g189(.a(\b[23] ), .b(\a[24] ), .o1(new_n285));
  nand42aa1n16x5               g190(.a(\b[23] ), .b(\a[24] ), .o1(new_n286));
  norb02aa1n02x5               g191(.a(new_n286), .b(new_n285), .out0(new_n287));
  aboi22aa1n03x5               g192(.a(new_n285), .b(new_n286), .c(new_n275), .d(new_n276), .out0(new_n288));
  aoi022aa1n03x5               g193(.a(new_n284), .b(new_n287), .c(new_n283), .d(new_n288), .o1(\s[24] ));
  nanb02aa1n03x5               g194(.a(new_n285), .b(new_n286), .out0(new_n290));
  nona22aa1n09x5               g195(.a(new_n270), .b(new_n290), .c(new_n279), .out0(new_n291));
  nano22aa1n03x7               g196(.a(new_n291), .b(new_n226), .c(new_n269), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n293));
  inv000aa1n06x5               g198(.a(new_n291), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n285), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n286), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n278), .b(new_n263), .c(new_n255), .d(new_n264), .o1(new_n297));
  aoai13aa1n06x5               g202(.a(new_n295), .b(new_n296), .c(new_n297), .d(new_n277), .o1(new_n298));
  aoi012aa1n02x5               g203(.a(new_n298), .b(new_n294), .c(new_n253), .o1(new_n299));
  inv000aa1n03x5               g204(.a(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[25] ), .b(\b[24] ), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n300), .c(new_n212), .d(new_n292), .o1(new_n302));
  oai012aa1n02x5               g207(.a(new_n231), .b(\b[19] ), .c(\a[20] ), .o1(new_n303));
  nona32aa1n02x4               g208(.a(new_n228), .b(new_n303), .c(new_n268), .d(new_n230), .out0(new_n304));
  tech160nm_fiaoi012aa1n04x5   g209(.a(new_n291), .b(new_n304), .c(new_n252), .o1(new_n305));
  norp03aa1n02x5               g210(.a(new_n305), .b(new_n298), .c(new_n301), .o1(new_n306));
  aobi12aa1n02x7               g211(.a(new_n302), .b(new_n306), .c(new_n293), .out0(\s[25] ));
  nor042aa1n03x5               g212(.a(\b[24] ), .b(\a[25] ), .o1(new_n308));
  inv000aa1n03x5               g213(.a(new_n308), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n301), .o1(new_n310));
  aoai13aa1n02x5               g215(.a(new_n309), .b(new_n310), .c(new_n293), .d(new_n299), .o1(new_n311));
  tech160nm_fixorc02aa1n02p5x5 g216(.a(\a[26] ), .b(\b[25] ), .out0(new_n312));
  norp02aa1n02x5               g217(.a(new_n312), .b(new_n308), .o1(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n302), .d(new_n313), .o1(\s[26] ));
  nanp02aa1n04x5               g219(.a(new_n312), .b(new_n301), .o1(new_n315));
  nano23aa1n06x5               g220(.a(new_n315), .b(new_n291), .c(new_n226), .d(new_n269), .out0(new_n316));
  inv020aa1n02x5               g221(.a(new_n315), .o1(new_n317));
  aoai13aa1n06x5               g222(.a(new_n317), .b(new_n298), .c(new_n294), .d(new_n253), .o1(new_n318));
  oaoi03aa1n12x5               g223(.a(\a[26] ), .b(\b[25] ), .c(new_n309), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n319), .o1(new_n320));
  nand42aa1n03x5               g225(.a(new_n318), .b(new_n320), .o1(new_n321));
  xorc02aa1n12x5               g226(.a(\a[27] ), .b(\b[26] ), .out0(new_n322));
  aoai13aa1n04x5               g227(.a(new_n322), .b(new_n321), .c(new_n212), .d(new_n316), .o1(new_n323));
  aoai13aa1n06x5               g228(.a(new_n316), .b(new_n221), .c(new_n143), .d(new_n203), .o1(new_n324));
  nano32aa1n03x7               g229(.a(new_n322), .b(new_n324), .c(new_n318), .d(new_n320), .out0(new_n325));
  norb02aa1n03x4               g230(.a(new_n323), .b(new_n325), .out0(\s[27] ));
  oaoi13aa1n09x5               g231(.a(new_n319), .b(new_n317), .c(new_n305), .d(new_n298), .o1(new_n327));
  norp02aa1n02x5               g232(.a(\b[26] ), .b(\a[27] ), .o1(new_n328));
  inv000aa1n03x5               g233(.a(new_n328), .o1(new_n329));
  inv000aa1n02x5               g234(.a(new_n322), .o1(new_n330));
  aoai13aa1n03x5               g235(.a(new_n329), .b(new_n330), .c(new_n324), .d(new_n327), .o1(new_n331));
  tech160nm_fixorc02aa1n03p5x5 g236(.a(\a[28] ), .b(\b[27] ), .out0(new_n332));
  norp02aa1n02x5               g237(.a(new_n332), .b(new_n328), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n331), .b(new_n332), .c(new_n323), .d(new_n333), .o1(\s[28] ));
  and002aa1n02x5               g239(.a(new_n332), .b(new_n322), .o(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n321), .c(new_n212), .d(new_n316), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n335), .o1(new_n337));
  oao003aa1n02x5               g242(.a(\a[28] ), .b(\b[27] ), .c(new_n329), .carry(new_n338));
  aoai13aa1n03x5               g243(.a(new_n338), .b(new_n337), .c(new_n324), .d(new_n327), .o1(new_n339));
  tech160nm_fixorc02aa1n03p5x5 g244(.a(\a[29] ), .b(\b[28] ), .out0(new_n340));
  norb02aa1n02x5               g245(.a(new_n338), .b(new_n340), .out0(new_n341));
  aoi022aa1n03x5               g246(.a(new_n339), .b(new_n340), .c(new_n336), .d(new_n341), .o1(\s[29] ));
  xorb03aa1n02x5               g247(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g248(.a(new_n330), .b(new_n332), .c(new_n340), .out0(new_n344));
  aoai13aa1n03x5               g249(.a(new_n344), .b(new_n321), .c(new_n212), .d(new_n316), .o1(new_n345));
  inv000aa1d42x5               g250(.a(new_n344), .o1(new_n346));
  oao003aa1n02x5               g251(.a(\a[29] ), .b(\b[28] ), .c(new_n338), .carry(new_n347));
  aoai13aa1n03x5               g252(.a(new_n347), .b(new_n346), .c(new_n324), .d(new_n327), .o1(new_n348));
  xorc02aa1n02x5               g253(.a(\a[30] ), .b(\b[29] ), .out0(new_n349));
  norb02aa1n02x5               g254(.a(new_n347), .b(new_n349), .out0(new_n350));
  aoi022aa1n03x5               g255(.a(new_n348), .b(new_n349), .c(new_n345), .d(new_n350), .o1(\s[30] ));
  nano32aa1n06x5               g256(.a(new_n330), .b(new_n349), .c(new_n332), .d(new_n340), .out0(new_n352));
  aoai13aa1n02x7               g257(.a(new_n352), .b(new_n321), .c(new_n212), .d(new_n316), .o1(new_n353));
  xorc02aa1n02x5               g258(.a(\a[31] ), .b(\b[30] ), .out0(new_n354));
  and002aa1n02x5               g259(.a(\b[29] ), .b(\a[30] ), .o(new_n355));
  oabi12aa1n02x5               g260(.a(new_n354), .b(\a[30] ), .c(\b[29] ), .out0(new_n356));
  oab012aa1n02x4               g261(.a(new_n356), .b(new_n347), .c(new_n355), .out0(new_n357));
  inv000aa1d42x5               g262(.a(new_n352), .o1(new_n358));
  oao003aa1n02x5               g263(.a(\a[30] ), .b(\b[29] ), .c(new_n347), .carry(new_n359));
  aoai13aa1n03x5               g264(.a(new_n359), .b(new_n358), .c(new_n324), .d(new_n327), .o1(new_n360));
  aoi022aa1n03x5               g265(.a(new_n360), .b(new_n354), .c(new_n353), .d(new_n357), .o1(\s[31] ));
  xnbna2aa1n03x5               g266(.a(new_n133), .b(new_n99), .c(new_n97), .out0(\s[3] ));
  norb02aa1n02x5               g267(.a(new_n103), .b(new_n104), .out0(new_n363));
  aoi012aa1n02x5               g268(.a(new_n100), .b(new_n132), .c(new_n133), .o1(new_n364));
  oai012aa1n02x5               g269(.a(new_n106), .b(new_n364), .c(new_n363), .o1(\s[4] ));
  xnrc02aa1n02x5               g270(.a(\b[4] ), .b(\a[5] ), .out0(new_n366));
  aoai13aa1n02x5               g271(.a(new_n103), .b(new_n134), .c(new_n132), .d(new_n133), .o1(new_n367));
  and002aa1n02x5               g272(.a(\b[4] ), .b(\a[5] ), .o(new_n368));
  aoi112aa1n02x5               g273(.a(new_n368), .b(new_n108), .c(\a[4] ), .d(\b[3] ), .o1(new_n369));
  aoi022aa1n02x5               g274(.a(new_n367), .b(new_n366), .c(new_n106), .d(new_n369), .o1(\s[5] ));
  aoai13aa1n02x5               g275(.a(new_n369), .b(new_n134), .c(new_n132), .d(new_n133), .o1(new_n371));
  xnbna2aa1n03x5               g276(.a(new_n122), .b(new_n371), .c(new_n116), .out0(\s[6] ));
  nanb02aa1n02x5               g277(.a(new_n139), .b(new_n371), .out0(new_n373));
  xnrc02aa1n02x5               g278(.a(\b[6] ), .b(\a[7] ), .out0(new_n374));
  aoai13aa1n02x5               g279(.a(new_n112), .b(new_n139), .c(new_n106), .d(new_n369), .o1(new_n375));
  aoi022aa1n02x5               g280(.a(new_n375), .b(new_n374), .c(new_n373), .d(new_n140), .o1(\s[7] ));
  aoi022aa1n02x5               g281(.a(new_n373), .b(new_n123), .c(new_n117), .d(new_n118), .o1(new_n377));
  xnrc02aa1n02x5               g282(.a(new_n377), .b(new_n141), .out0(\s[8] ));
  xorb03aa1n02x5               g283(.a(new_n143), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


