// Benchmark "adder" written by ABC on Wed Jul 17 19:11:34 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n345,
    new_n346, new_n349, new_n351, new_n352, new_n353, new_n355, new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d30x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  and002aa1n24x5               g004(.a(\b[3] ), .b(\a[4] ), .o(new_n100));
  inv020aa1n12x5               g005(.a(\a[3] ), .o1(new_n101));
  inv040aa1n08x5               g006(.a(\b[2] ), .o1(new_n102));
  nor042aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  aoi112aa1n09x5               g008(.a(new_n100), .b(new_n103), .c(new_n101), .d(new_n102), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(new_n102), .b(new_n101), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n03x5               g011(.a(new_n105), .b(new_n106), .o1(new_n107));
  nor042aa1n02x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nand02aa1n04x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  nanp02aa1n04x5               g014(.a(\b[1] ), .b(\a[2] ), .o1(new_n110));
  aoi012aa1n12x5               g015(.a(new_n108), .b(new_n109), .c(new_n110), .o1(new_n111));
  oaoi13aa1n12x5               g016(.a(new_n100), .b(new_n104), .c(new_n111), .d(new_n107), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[4] ), .o1(new_n114));
  nanb02aa1d24x5               g019(.a(\a[5] ), .b(new_n114), .out0(new_n115));
  nor002aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  norb02aa1n02x5               g022(.a(new_n117), .b(new_n116), .out0(new_n118));
  nanp02aa1n04x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nor022aa1n06x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nand42aa1n04x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nor002aa1d24x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  nona23aa1n03x5               g027(.a(new_n121), .b(new_n119), .c(new_n122), .d(new_n120), .out0(new_n123));
  nano32aa1n03x7               g028(.a(new_n123), .b(new_n118), .c(new_n115), .d(new_n113), .out0(new_n124));
  oai012aa1n02x5               g029(.a(new_n121), .b(new_n122), .c(new_n120), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[6] ), .b(\b[5] ), .c(new_n115), .o1(new_n126));
  oaib12aa1n06x5               g031(.a(new_n125), .b(new_n123), .c(new_n126), .out0(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n129));
  nor002aa1d32x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1d28x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g038(.a(new_n130), .o1(new_n134));
  inv000aa1n02x5               g039(.a(new_n131), .o1(new_n135));
  nor002aa1n16x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand42aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x7               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  aoi113aa1n03x7               g044(.a(new_n139), .b(new_n135), .c(new_n129), .d(new_n134), .e(new_n99), .o1(new_n140));
  nanp02aa1n03x5               g045(.a(new_n129), .b(new_n99), .o1(new_n141));
  aoai13aa1n12x5               g046(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  aoi112aa1n02x5               g048(.a(new_n143), .b(new_n138), .c(new_n141), .d(new_n132), .o1(new_n144));
  norp02aa1n02x5               g049(.a(new_n144), .b(new_n140), .o1(\s[11] ));
  inv000aa1d42x5               g050(.a(new_n136), .o1(new_n146));
  nor042aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand42aa1n04x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nano22aa1n02x4               g055(.a(new_n140), .b(new_n146), .c(new_n150), .out0(new_n151));
  aoai13aa1n03x5               g056(.a(new_n138), .b(new_n143), .c(new_n141), .d(new_n132), .o1(new_n152));
  aoi012aa1n03x5               g057(.a(new_n150), .b(new_n152), .c(new_n146), .o1(new_n153));
  nor002aa1n02x5               g058(.a(new_n153), .b(new_n151), .o1(\s[12] ));
  and002aa1n06x5               g059(.a(\b[8] ), .b(\a[9] ), .o(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nona23aa1n09x5               g061(.a(new_n148), .b(new_n137), .c(new_n136), .d(new_n147), .out0(new_n157));
  nano32aa1n02x4               g062(.a(new_n157), .b(new_n132), .c(new_n156), .d(new_n99), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n159));
  tech160nm_fioai012aa1n03p5x5 g064(.a(new_n148), .b(new_n147), .c(new_n136), .o1(new_n160));
  oai012aa1d24x5               g065(.a(new_n160), .b(new_n157), .c(new_n142), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(new_n159), .b(new_n162), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g069(.a(\a[13] ), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[12] ), .o1(new_n166));
  oaoi03aa1n02x5               g071(.a(new_n165), .b(new_n166), .c(new_n163), .o1(new_n167));
  xnrb03aa1n02x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n06x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  tech160nm_finand02aa1n03p5x5 g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n169), .c(new_n165), .d(new_n166), .o1(new_n171));
  norp02aa1n02x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  nand42aa1n02x5               g077(.a(\b[12] ), .b(\a[13] ), .o1(new_n173));
  nona23aa1n03x5               g078(.a(new_n170), .b(new_n173), .c(new_n172), .d(new_n169), .out0(new_n174));
  aoai13aa1n04x5               g079(.a(new_n171), .b(new_n174), .c(new_n159), .d(new_n162), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanp02aa1n04x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nor022aa1n16x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand42aa1n03x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  aoi112aa1n02x5               g087(.a(new_n182), .b(new_n177), .c(new_n175), .d(new_n178), .o1(new_n183));
  aoai13aa1n03x5               g088(.a(new_n182), .b(new_n177), .c(new_n175), .d(new_n178), .o1(new_n184));
  norb02aa1n03x4               g089(.a(new_n184), .b(new_n183), .out0(\s[16] ));
  aoi112aa1n02x5               g090(.a(new_n135), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n186));
  nano23aa1n02x4               g091(.a(new_n136), .b(new_n147), .c(new_n148), .d(new_n137), .out0(new_n187));
  nano23aa1n02x5               g092(.a(new_n172), .b(new_n169), .c(new_n170), .d(new_n173), .out0(new_n188));
  nano23aa1n02x5               g093(.a(new_n177), .b(new_n179), .c(new_n180), .d(new_n178), .out0(new_n189));
  nanp02aa1n02x5               g094(.a(new_n189), .b(new_n188), .o1(new_n190));
  nano32aa1n03x7               g095(.a(new_n190), .b(new_n187), .c(new_n186), .d(new_n156), .out0(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n192));
  nona23aa1n02x4               g097(.a(new_n180), .b(new_n178), .c(new_n177), .d(new_n179), .out0(new_n193));
  nor002aa1n03x5               g098(.a(new_n193), .b(new_n174), .o1(new_n194));
  oa0012aa1n02x5               g099(.a(new_n180), .b(new_n179), .c(new_n177), .o(new_n195));
  norp02aa1n03x5               g100(.a(new_n193), .b(new_n171), .o1(new_n196));
  aoi112aa1n09x5               g101(.a(new_n196), .b(new_n195), .c(new_n161), .d(new_n194), .o1(new_n197));
  nand02aa1d08x5               g102(.a(new_n192), .b(new_n197), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g104(.a(\a[17] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[16] ), .o1(new_n201));
  oaoi03aa1n03x5               g106(.a(new_n200), .b(new_n201), .c(new_n198), .o1(new_n202));
  xnrb03aa1n03x5               g107(.a(new_n202), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n02x5               g108(.a(new_n201), .b(new_n200), .o1(new_n204));
  nanp02aa1n02x5               g109(.a(\b[16] ), .b(\a[17] ), .o1(new_n205));
  nor022aa1n06x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand42aa1n03x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nanb02aa1n02x5               g112(.a(new_n206), .b(new_n207), .out0(new_n208));
  nano22aa1n12x5               g113(.a(new_n208), .b(new_n204), .c(new_n205), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n207), .b(new_n206), .c(new_n200), .d(new_n201), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n210), .c(new_n192), .d(new_n197), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nanp02aa1n02x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  nor042aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoi112aa1n02x7               g125(.a(new_n215), .b(new_n220), .c(new_n212), .d(new_n216), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n215), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n216), .b(new_n215), .out0(new_n223));
  nanp02aa1n03x5               g128(.a(new_n212), .b(new_n223), .o1(new_n224));
  aoi012aa1n03x5               g129(.a(new_n219), .b(new_n224), .c(new_n222), .o1(new_n225));
  nor002aa1n02x5               g130(.a(new_n225), .b(new_n221), .o1(\s[20] ));
  nano23aa1n03x7               g131(.a(new_n215), .b(new_n217), .c(new_n218), .d(new_n216), .out0(new_n227));
  nanp02aa1n02x5               g132(.a(new_n209), .b(new_n227), .o1(new_n228));
  inv000aa1n02x5               g133(.a(new_n211), .o1(new_n229));
  tech160nm_fioai012aa1n04x5   g134(.a(new_n218), .b(new_n217), .c(new_n215), .o1(new_n230));
  aobi12aa1n06x5               g135(.a(new_n230), .b(new_n227), .c(new_n229), .out0(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n228), .c(new_n192), .d(new_n197), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  nand42aa1n02x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  xorc02aa1n02x5               g140(.a(\a[22] ), .b(\b[21] ), .out0(new_n236));
  aoi112aa1n03x4               g141(.a(new_n234), .b(new_n236), .c(new_n232), .d(new_n235), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n234), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n235), .b(new_n234), .out0(new_n239));
  nanp02aa1n02x5               g144(.a(new_n232), .b(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n236), .o1(new_n241));
  tech160nm_fiaoi012aa1n04x5   g146(.a(new_n241), .b(new_n240), .c(new_n238), .o1(new_n242));
  norp02aa1n03x5               g147(.a(new_n242), .b(new_n237), .o1(\s[22] ));
  norp02aa1n02x5               g148(.a(\b[21] ), .b(\a[22] ), .o1(new_n244));
  nanp02aa1n02x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  nano23aa1n03x7               g150(.a(new_n234), .b(new_n244), .c(new_n245), .d(new_n235), .out0(new_n246));
  nand23aa1n02x5               g151(.a(new_n209), .b(new_n227), .c(new_n246), .o1(new_n247));
  nona23aa1n03x5               g152(.a(new_n218), .b(new_n216), .c(new_n215), .d(new_n217), .out0(new_n248));
  tech160nm_fioai012aa1n05x5   g153(.a(new_n230), .b(new_n248), .c(new_n211), .o1(new_n249));
  oaoi03aa1n02x5               g154(.a(\a[22] ), .b(\b[21] ), .c(new_n238), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n250), .b(new_n249), .c(new_n246), .o1(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n247), .c(new_n192), .d(new_n197), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  nor042aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nand42aa1n02x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  norb02aa1n02x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  aoi112aa1n03x4               g163(.a(new_n254), .b(new_n258), .c(new_n252), .d(new_n255), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n254), .o1(new_n260));
  norb02aa1n02x5               g165(.a(new_n255), .b(new_n254), .out0(new_n261));
  nand02aa1n02x5               g166(.a(new_n252), .b(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n258), .o1(new_n263));
  aoi012aa1n02x5               g168(.a(new_n263), .b(new_n262), .c(new_n260), .o1(new_n264));
  nor002aa1n02x5               g169(.a(new_n264), .b(new_n259), .o1(\s[24] ));
  nano23aa1n06x5               g170(.a(new_n254), .b(new_n256), .c(new_n257), .d(new_n255), .out0(new_n266));
  nanb03aa1n02x5               g171(.a(new_n228), .b(new_n266), .c(new_n246), .out0(new_n267));
  nona22aa1n02x4               g172(.a(new_n257), .b(new_n256), .c(new_n254), .out0(new_n268));
  aoi022aa1n03x5               g173(.a(new_n266), .b(new_n250), .c(new_n268), .d(new_n257), .o1(new_n269));
  inv020aa1n03x5               g174(.a(new_n269), .o1(new_n270));
  aoi013aa1n02x4               g175(.a(new_n270), .b(new_n249), .c(new_n246), .d(new_n266), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n267), .c(new_n192), .d(new_n197), .o1(new_n272));
  xorb03aa1n02x5               g177(.a(new_n272), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xnrc02aa1n12x5               g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoi112aa1n02x7               g182(.a(new_n274), .b(new_n277), .c(new_n272), .d(new_n275), .o1(new_n278));
  inv020aa1n02x5               g183(.a(new_n274), .o1(new_n279));
  norb02aa1n02x5               g184(.a(new_n275), .b(new_n274), .out0(new_n280));
  nand42aa1n02x5               g185(.a(new_n272), .b(new_n280), .o1(new_n281));
  aoi012aa1n03x5               g186(.a(new_n276), .b(new_n281), .c(new_n279), .o1(new_n282));
  norp02aa1n03x5               g187(.a(new_n282), .b(new_n278), .o1(\s[26] ));
  inv000aa1d42x5               g188(.a(new_n100), .o1(new_n284));
  oaih12aa1n02x5               g189(.a(new_n104), .b(new_n111), .c(new_n107), .o1(new_n285));
  nanp02aa1n03x5               g190(.a(new_n285), .b(new_n284), .o1(new_n286));
  nano22aa1n02x4               g191(.a(new_n116), .b(new_n115), .c(new_n117), .out0(new_n287));
  nano23aa1n02x4               g192(.a(new_n122), .b(new_n120), .c(new_n119), .d(new_n121), .out0(new_n288));
  nanp03aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n113), .o1(new_n289));
  aobi12aa1n02x5               g194(.a(new_n125), .b(new_n288), .c(new_n126), .out0(new_n290));
  oai012aa1n02x7               g195(.a(new_n290), .b(new_n286), .c(new_n289), .o1(new_n291));
  nand42aa1n02x5               g196(.a(new_n161), .b(new_n194), .o1(new_n292));
  nona22aa1n03x5               g197(.a(new_n292), .b(new_n196), .c(new_n195), .out0(new_n293));
  nano22aa1n06x5               g198(.a(new_n276), .b(new_n279), .c(new_n275), .out0(new_n294));
  nano22aa1n03x7               g199(.a(new_n247), .b(new_n266), .c(new_n294), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n293), .c(new_n291), .d(new_n191), .o1(new_n296));
  nano22aa1n03x7               g201(.a(new_n231), .b(new_n246), .c(new_n266), .out0(new_n297));
  oaoi03aa1n02x5               g202(.a(\a[26] ), .b(\b[25] ), .c(new_n279), .o1(new_n298));
  oaoi13aa1n09x5               g203(.a(new_n298), .b(new_n294), .c(new_n297), .d(new_n270), .o1(new_n299));
  norp02aa1n04x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  nand42aa1n03x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  norb02aa1n02x5               g206(.a(new_n301), .b(new_n300), .out0(new_n302));
  xnbna2aa1n03x5               g207(.a(new_n302), .b(new_n296), .c(new_n299), .out0(\s[27] ));
  inv040aa1n02x5               g208(.a(new_n300), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n302), .o1(new_n305));
  aoi012aa1n02x5               g210(.a(new_n305), .b(new_n296), .c(new_n299), .o1(new_n306));
  xnrc02aa1n12x5               g211(.a(\b[27] ), .b(\a[28] ), .out0(new_n307));
  nano22aa1n02x4               g212(.a(new_n306), .b(new_n304), .c(new_n307), .out0(new_n308));
  nanp03aa1n03x5               g213(.a(new_n249), .b(new_n246), .c(new_n266), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n294), .o1(new_n310));
  inv000aa1n02x5               g215(.a(new_n298), .o1(new_n311));
  aoai13aa1n06x5               g216(.a(new_n311), .b(new_n310), .c(new_n309), .d(new_n269), .o1(new_n312));
  aoai13aa1n06x5               g217(.a(new_n302), .b(new_n312), .c(new_n198), .d(new_n295), .o1(new_n313));
  tech160nm_fiaoi012aa1n05x5   g218(.a(new_n307), .b(new_n313), .c(new_n304), .o1(new_n314));
  norp02aa1n03x5               g219(.a(new_n314), .b(new_n308), .o1(\s[28] ));
  xnrc02aa1n12x5               g220(.a(\b[28] ), .b(\a[29] ), .out0(new_n316));
  nano22aa1n03x7               g221(.a(new_n307), .b(new_n304), .c(new_n301), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n312), .c(new_n198), .d(new_n295), .o1(new_n318));
  oao003aa1n02x5               g223(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n319));
  aoi012aa1n03x5               g224(.a(new_n316), .b(new_n318), .c(new_n319), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n317), .o1(new_n321));
  tech160nm_fiaoi012aa1n02p5x5 g226(.a(new_n321), .b(new_n296), .c(new_n299), .o1(new_n322));
  nano22aa1n02x4               g227(.a(new_n322), .b(new_n316), .c(new_n319), .out0(new_n323));
  norp02aa1n03x5               g228(.a(new_n320), .b(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1d15x5               g230(.a(new_n316), .b(new_n307), .c(new_n301), .d(new_n304), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n312), .c(new_n198), .d(new_n295), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .c(new_n319), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[29] ), .b(\a[30] ), .out0(new_n329));
  aoi012aa1n03x5               g234(.a(new_n329), .b(new_n327), .c(new_n328), .o1(new_n330));
  inv000aa1d42x5               g235(.a(new_n326), .o1(new_n331));
  tech160nm_fiaoi012aa1n02p5x5 g236(.a(new_n331), .b(new_n296), .c(new_n299), .o1(new_n332));
  nano22aa1n03x5               g237(.a(new_n332), .b(new_n328), .c(new_n329), .out0(new_n333));
  norp02aa1n03x5               g238(.a(new_n330), .b(new_n333), .o1(\s[30] ));
  norb03aa1d15x5               g239(.a(new_n317), .b(new_n316), .c(new_n329), .out0(new_n335));
  inv000aa1d42x5               g240(.a(new_n335), .o1(new_n336));
  tech160nm_fiaoi012aa1n02p5x5 g241(.a(new_n336), .b(new_n296), .c(new_n299), .o1(new_n337));
  oao003aa1n02x5               g242(.a(\a[30] ), .b(\b[29] ), .c(new_n328), .carry(new_n338));
  xnrc02aa1n02x5               g243(.a(\b[30] ), .b(\a[31] ), .out0(new_n339));
  nano22aa1n02x4               g244(.a(new_n337), .b(new_n338), .c(new_n339), .out0(new_n340));
  aoai13aa1n03x5               g245(.a(new_n335), .b(new_n312), .c(new_n198), .d(new_n295), .o1(new_n341));
  aoi012aa1n03x5               g246(.a(new_n339), .b(new_n341), .c(new_n338), .o1(new_n342));
  nor002aa1n02x5               g247(.a(new_n342), .b(new_n340), .o1(\s[31] ));
  xnbna2aa1n03x5               g248(.a(new_n111), .b(new_n105), .c(new_n106), .out0(\s[3] ));
  xnrc02aa1n02x5               g249(.a(\b[3] ), .b(\a[4] ), .out0(new_n345));
  oaoi03aa1n02x5               g250(.a(\a[3] ), .b(\b[2] ), .c(new_n111), .o1(new_n346));
  aob012aa1n02x5               g251(.a(new_n285), .b(new_n346), .c(new_n345), .out0(\s[4] ));
  xorb03aa1n02x5               g252(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g253(.a(\a[5] ), .b(\b[4] ), .c(new_n286), .o1(new_n349));
  xorb03aa1n02x5               g254(.a(new_n349), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g255(.a(new_n119), .b(new_n122), .out0(new_n351));
  oai112aa1n02x5               g256(.a(new_n351), .b(new_n117), .c(new_n349), .d(new_n116), .o1(new_n352));
  oaoi13aa1n02x5               g257(.a(new_n351), .b(new_n117), .c(new_n349), .d(new_n116), .o1(new_n353));
  norb02aa1n02x5               g258(.a(new_n352), .b(new_n353), .out0(\s[7] ));
  norb02aa1n02x5               g259(.a(new_n121), .b(new_n120), .out0(new_n355));
  inv000aa1d42x5               g260(.a(new_n122), .o1(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n355), .b(new_n352), .c(new_n356), .out0(\s[8] ));
  xorb03aa1n02x5               g262(.a(new_n291), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


