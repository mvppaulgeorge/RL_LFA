// Benchmark "adder" written by ABC on Wed Jul 17 17:22:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n356, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n364, new_n366, new_n367, new_n369, new_n370,
    new_n371, new_n373;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv030aa1n02x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n08x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norb03aa1n03x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  tech160nm_fixnrc02aa1n04x5   g007(.a(\b[3] ), .b(\a[4] ), .out0(new_n103));
  nand42aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nor022aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb03aa1n02x5               g010(.a(new_n105), .b(new_n100), .c(new_n104), .out0(new_n106));
  norp02aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  aob012aa1n06x5               g012(.a(new_n105), .b(\b[3] ), .c(\a[4] ), .out0(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  oai013aa1n03x5               g014(.a(new_n109), .b(new_n102), .c(new_n106), .d(new_n103), .o1(new_n110));
  xorc02aa1n02x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  nanp02aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  oai012aa1n02x5               g017(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .o1(new_n113));
  aoi022aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n114));
  oai122aa1n02x7               g019(.a(new_n114), .b(\a[6] ), .c(\b[5] ), .d(\a[5] ), .e(\b[4] ), .o1(new_n115));
  norb03aa1n03x5               g020(.a(new_n111), .b(new_n115), .c(new_n113), .out0(new_n116));
  oai022aa1n02x5               g021(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n117));
  aob012aa1n02x5               g022(.a(new_n117), .b(\b[7] ), .c(\a[8] ), .out0(new_n118));
  oai122aa1n02x7               g023(.a(new_n112), .b(\a[8] ), .c(\b[7] ), .d(\a[7] ), .e(\b[6] ), .o1(new_n119));
  oai022aa1n02x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  aoi022aa1n02x5               g025(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n120), .b(new_n121), .o1(new_n122));
  tech160nm_fioai012aa1n05x5   g027(.a(new_n118), .b(new_n122), .c(new_n119), .o1(new_n123));
  xnrc02aa1n12x5               g028(.a(\b[8] ), .b(\a[9] ), .out0(new_n124));
  inv000aa1d42x5               g029(.a(new_n124), .o1(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n123), .c(new_n110), .d(new_n116), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n127), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g033(.a(new_n127), .o1(new_n129));
  aoi012aa1n02x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .o1(new_n130));
  aoi112aa1n02x5               g035(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n131));
  tech160nm_fioaoi03aa1n03p5x5 g036(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n132));
  nand42aa1n03x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb02aa1n03x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  oai012aa1n02x5               g040(.a(new_n135), .b(new_n130), .c(new_n132), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n134), .o1(new_n137));
  oai112aa1n02x5               g042(.a(new_n137), .b(new_n133), .c(\b[9] ), .d(\a[10] ), .o1(new_n138));
  oai013aa1n02x4               g043(.a(new_n136), .b(new_n131), .c(new_n130), .d(new_n138), .o1(\s[11] ));
  norp02aa1n02x5               g044(.a(\b[9] ), .b(\a[10] ), .o1(new_n140));
  norp03aa1n02x5               g045(.a(new_n131), .b(new_n134), .c(new_n140), .o1(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n129), .c(new_n126), .d(new_n98), .o1(new_n142));
  xorc02aa1n12x5               g047(.a(\a[12] ), .b(\b[11] ), .out0(new_n143));
  xobna2aa1n03x5               g048(.a(new_n143), .b(new_n142), .c(new_n133), .out0(\s[12] ));
  nona22aa1n06x5               g049(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n145));
  nano22aa1n03x7               g050(.a(new_n105), .b(new_n100), .c(new_n104), .out0(new_n146));
  nanb03aa1n03x5               g051(.a(new_n103), .b(new_n146), .c(new_n145), .out0(new_n147));
  nona23aa1n02x4               g052(.a(new_n111), .b(new_n114), .c(new_n113), .d(new_n120), .out0(new_n148));
  inv000aa1n02x5               g053(.a(new_n123), .o1(new_n149));
  aoai13aa1n04x5               g054(.a(new_n149), .b(new_n148), .c(new_n147), .d(new_n109), .o1(new_n150));
  nona23aa1d18x5               g055(.a(new_n143), .b(new_n127), .c(new_n124), .d(new_n135), .out0(new_n151));
  nanb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  nanp02aa1n02x5               g057(.a(new_n110), .b(new_n116), .o1(new_n153));
  nanb03aa1n06x5               g058(.a(new_n135), .b(new_n132), .c(new_n143), .out0(new_n154));
  oao003aa1n02x5               g059(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .carry(new_n155));
  nanp02aa1n02x5               g060(.a(new_n154), .b(new_n155), .o1(new_n156));
  inv040aa1n03x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n04x5               g062(.a(new_n157), .b(new_n151), .c(new_n153), .d(new_n149), .o1(new_n158));
  xorc02aa1n12x5               g063(.a(\a[13] ), .b(\b[12] ), .out0(new_n159));
  nano22aa1n02x4               g064(.a(new_n159), .b(new_n154), .c(new_n155), .out0(new_n160));
  aoi022aa1n02x5               g065(.a(new_n158), .b(new_n159), .c(new_n152), .d(new_n160), .o1(\s[13] ));
  nor042aa1d18x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  inv040aa1n08x5               g067(.a(new_n162), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(new_n158), .b(new_n159), .o1(new_n164));
  xorc02aa1n12x5               g069(.a(\a[14] ), .b(\b[13] ), .out0(new_n165));
  inv000aa1d42x5               g070(.a(\a[14] ), .o1(new_n166));
  inv000aa1d42x5               g071(.a(\b[13] ), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n162), .b(new_n166), .c(new_n167), .o1(new_n168));
  oai112aa1n02x5               g073(.a(new_n164), .b(new_n168), .c(new_n167), .d(new_n166), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n165), .c(new_n163), .d(new_n164), .o1(\s[14] ));
  inv000aa1d42x5               g075(.a(\a[13] ), .o1(new_n171));
  xroi22aa1d04x5               g076(.a(new_n171), .b(\b[12] ), .c(new_n166), .d(\b[13] ), .out0(new_n172));
  oaoi03aa1n12x5               g077(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n173));
  xorc02aa1n02x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  aoai13aa1n04x5               g079(.a(new_n174), .b(new_n173), .c(new_n158), .d(new_n172), .o1(new_n175));
  aoi112aa1n02x5               g080(.a(new_n174), .b(new_n173), .c(new_n158), .d(new_n172), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(\s[15] ));
  nor042aa1n12x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  nor042aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nand42aa1n20x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n181), .b(new_n180), .out0(new_n182));
  norb03aa1n02x5               g087(.a(new_n181), .b(new_n178), .c(new_n180), .out0(new_n183));
  nand42aa1n03x5               g088(.a(new_n175), .b(new_n183), .o1(new_n184));
  aoai13aa1n03x5               g089(.a(new_n184), .b(new_n182), .c(new_n179), .d(new_n175), .o1(\s[16] ));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  nand42aa1d28x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  nano23aa1d12x5               g092(.a(new_n180), .b(new_n178), .c(new_n181), .d(new_n187), .out0(new_n188));
  nand23aa1n09x5               g093(.a(new_n188), .b(new_n159), .c(new_n165), .o1(new_n189));
  nor042aa1n09x5               g094(.a(new_n151), .b(new_n189), .o1(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n123), .c(new_n110), .d(new_n116), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  aoi112aa1n02x5               g097(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n193));
  aoi112aa1n06x5               g098(.a(new_n193), .b(new_n180), .c(new_n188), .d(new_n173), .o1(new_n194));
  aoai13aa1n12x5               g099(.a(new_n194), .b(new_n189), .c(new_n154), .d(new_n155), .o1(new_n195));
  inv040aa1d30x5               g100(.a(new_n195), .o1(new_n196));
  nanp02aa1n12x5               g101(.a(new_n191), .b(new_n196), .o1(new_n197));
  inv000aa1d42x5               g102(.a(new_n189), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(new_n156), .b(new_n198), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n173), .o1(new_n200));
  nano22aa1n02x4               g105(.a(new_n200), .b(new_n174), .c(new_n182), .out0(new_n201));
  inv000aa1d42x5               g106(.a(\a[17] ), .o1(new_n202));
  inv000aa1d42x5               g107(.a(\b[16] ), .o1(new_n203));
  oai022aa1n02x5               g108(.a(\a[16] ), .b(\b[15] ), .c(\b[16] ), .d(\a[17] ), .o1(new_n204));
  oabi12aa1n02x5               g109(.a(new_n204), .b(new_n202), .c(new_n203), .out0(new_n205));
  nona32aa1n02x4               g110(.a(new_n199), .b(new_n205), .c(new_n193), .d(new_n201), .out0(new_n206));
  obai22aa1n02x7               g111(.a(new_n197), .b(new_n186), .c(new_n206), .d(new_n192), .out0(\s[17] ));
  xnrc02aa1n02x5               g112(.a(\b[17] ), .b(\a[18] ), .out0(new_n208));
  nona32aa1n02x4               g113(.a(new_n199), .b(new_n204), .c(new_n193), .d(new_n201), .out0(new_n209));
  nanb02aa1n02x5               g114(.a(new_n209), .b(new_n191), .out0(new_n210));
  obai22aa1n02x5               g115(.a(new_n191), .b(new_n209), .c(new_n202), .d(new_n203), .out0(new_n211));
  oai022aa1n02x5               g116(.a(new_n202), .b(new_n203), .c(\b[17] ), .d(\a[18] ), .o1(new_n212));
  aoi012aa1n02x5               g117(.a(new_n212), .b(\a[18] ), .c(\b[17] ), .o1(new_n213));
  aoi022aa1n02x5               g118(.a(new_n211), .b(new_n208), .c(new_n210), .d(new_n213), .o1(\s[18] ));
  inv000aa1d42x5               g119(.a(\a[18] ), .o1(new_n215));
  xroi22aa1d04x5               g120(.a(new_n202), .b(\b[16] ), .c(new_n215), .d(\b[17] ), .out0(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n195), .c(new_n150), .d(new_n190), .o1(new_n217));
  aoi112aa1n03x5               g122(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n218));
  aoib12aa1n06x5               g123(.a(new_n218), .b(new_n215), .c(\b[17] ), .out0(new_n219));
  nand22aa1n06x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nor002aa1d32x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n220), .b(new_n221), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n217), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n08x5               g129(.a(new_n221), .o1(new_n225));
  nor042aa1n06x5               g130(.a(\b[16] ), .b(\a[17] ), .o1(new_n226));
  aob012aa1n02x5               g131(.a(new_n226), .b(\b[17] ), .c(\a[18] ), .out0(new_n227));
  oaib12aa1n09x5               g132(.a(new_n227), .b(\b[17] ), .c(new_n215), .out0(new_n228));
  aoai13aa1n03x5               g133(.a(new_n222), .b(new_n228), .c(new_n197), .d(new_n216), .o1(new_n229));
  nor042aa1n06x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nand02aa1n06x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n222), .o1(new_n233));
  norb03aa1n02x5               g138(.a(new_n231), .b(new_n221), .c(new_n230), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n233), .c(new_n217), .d(new_n219), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n232), .c(new_n229), .d(new_n225), .o1(\s[20] ));
  nona23aa1n09x5               g141(.a(new_n220), .b(new_n231), .c(new_n230), .d(new_n221), .out0(new_n237));
  norb03aa1n03x5               g142(.a(new_n186), .b(new_n237), .c(new_n208), .out0(new_n238));
  aoai13aa1n02x5               g143(.a(new_n238), .b(new_n195), .c(new_n150), .d(new_n190), .o1(new_n239));
  oaoi03aa1n12x5               g144(.a(\a[20] ), .b(\b[19] ), .c(new_n225), .o1(new_n240));
  inv040aa1n02x5               g145(.a(new_n240), .o1(new_n241));
  oai012aa1n12x5               g146(.a(new_n241), .b(new_n237), .c(new_n219), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[20] ), .b(\a[21] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n242), .c(new_n197), .d(new_n238), .o1(new_n245));
  nano23aa1d12x5               g150(.a(new_n230), .b(new_n221), .c(new_n231), .d(new_n220), .out0(new_n246));
  aoi112aa1n02x5               g151(.a(new_n240), .b(new_n244), .c(new_n246), .d(new_n228), .o1(new_n247));
  aobi12aa1n03x7               g152(.a(new_n245), .b(new_n247), .c(new_n239), .out0(\s[21] ));
  nor042aa1n06x5               g153(.a(\b[20] ), .b(\a[21] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  xnrc02aa1n12x5               g155(.a(\b[21] ), .b(\a[22] ), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n242), .o1(new_n253));
  oai022aa1n02x5               g158(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n254));
  aoi012aa1n02x5               g159(.a(new_n254), .b(\a[22] ), .c(\b[21] ), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n243), .c(new_n239), .d(new_n253), .o1(new_n256));
  aoai13aa1n03x5               g161(.a(new_n256), .b(new_n252), .c(new_n245), .d(new_n250), .o1(\s[22] ));
  nor042aa1n06x5               g162(.a(new_n251), .b(new_n243), .o1(new_n258));
  and003aa1n02x5               g163(.a(new_n216), .b(new_n258), .c(new_n246), .o(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n195), .c(new_n150), .d(new_n190), .o1(new_n260));
  aoai13aa1n12x5               g165(.a(new_n258), .b(new_n240), .c(new_n246), .d(new_n228), .o1(new_n261));
  oaoi03aa1n12x5               g166(.a(\a[22] ), .b(\b[21] ), .c(new_n250), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(new_n261), .b(new_n263), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  nor042aa1n02x5               g170(.a(\b[22] ), .b(\a[23] ), .o1(new_n266));
  nand42aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .o1(new_n267));
  norb02aa1n02x5               g172(.a(new_n267), .b(new_n266), .out0(new_n268));
  inv000aa1d42x5               g173(.a(new_n261), .o1(new_n269));
  nona23aa1n02x4               g174(.a(new_n260), .b(new_n268), .c(new_n262), .d(new_n269), .out0(new_n270));
  aoai13aa1n02x5               g175(.a(new_n270), .b(new_n268), .c(new_n260), .d(new_n265), .o1(\s[23] ));
  nor042aa1n03x5               g176(.a(\b[23] ), .b(\a[24] ), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(\b[23] ), .b(\a[24] ), .o1(new_n273));
  nanb02aa1n02x5               g178(.a(new_n272), .b(new_n273), .out0(new_n274));
  nona32aa1n02x4               g179(.a(new_n260), .b(new_n266), .c(new_n262), .d(new_n269), .out0(new_n275));
  nanp02aa1n02x5               g180(.a(new_n275), .b(new_n267), .o1(new_n276));
  nano22aa1n02x4               g181(.a(new_n272), .b(new_n267), .c(new_n273), .out0(new_n277));
  aoi022aa1n02x7               g182(.a(new_n276), .b(new_n274), .c(new_n275), .d(new_n277), .o1(\s[24] ));
  nano23aa1d12x5               g183(.a(new_n266), .b(new_n272), .c(new_n273), .d(new_n267), .out0(new_n279));
  inv040aa1n02x5               g184(.a(new_n279), .o1(new_n280));
  nano32aa1n02x4               g185(.a(new_n280), .b(new_n216), .c(new_n258), .d(new_n246), .out0(new_n281));
  aoai13aa1n02x5               g186(.a(new_n281), .b(new_n195), .c(new_n150), .d(new_n190), .o1(new_n282));
  oai012aa1n02x5               g187(.a(new_n273), .b(new_n272), .c(new_n266), .o1(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n280), .c(new_n261), .d(new_n263), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n284), .c(new_n197), .d(new_n281), .o1(new_n286));
  aoai13aa1n02x5               g191(.a(new_n279), .b(new_n262), .c(new_n242), .d(new_n258), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  and003aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n283), .o(new_n289));
  aobi12aa1n03x7               g194(.a(new_n286), .b(new_n289), .c(new_n282), .out0(\s[25] ));
  norp02aa1n02x5               g195(.a(\b[24] ), .b(\a[25] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .out0(new_n293));
  inv000aa1n02x5               g198(.a(new_n284), .o1(new_n294));
  nanp02aa1n02x5               g199(.a(\b[25] ), .b(\a[26] ), .o1(new_n295));
  oai022aa1n02x5               g200(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n296));
  norb02aa1n02x5               g201(.a(new_n295), .b(new_n296), .out0(new_n297));
  aoai13aa1n02x7               g202(.a(new_n297), .b(new_n288), .c(new_n282), .d(new_n294), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n293), .c(new_n286), .d(new_n292), .o1(\s[26] ));
  and002aa1n06x5               g204(.a(new_n293), .b(new_n285), .o(new_n300));
  inv000aa1n02x5               g205(.a(new_n300), .o1(new_n301));
  nano32aa1n03x7               g206(.a(new_n301), .b(new_n238), .c(new_n258), .d(new_n279), .out0(new_n302));
  aoai13aa1n04x5               g207(.a(new_n302), .b(new_n195), .c(new_n150), .d(new_n190), .o1(new_n303));
  aoi022aa1n12x5               g208(.a(new_n284), .b(new_n300), .c(new_n295), .d(new_n296), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[27] ), .b(\b[26] ), .out0(new_n305));
  nand22aa1n03x5               g210(.a(new_n284), .b(new_n300), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(new_n296), .b(new_n295), .o1(new_n307));
  and002aa1n02x5               g212(.a(new_n305), .b(new_n307), .o(new_n308));
  nanp03aa1n02x5               g213(.a(new_n303), .b(new_n306), .c(new_n308), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n303), .d(new_n304), .o1(\s[27] ));
  xnrc02aa1n02x5               g215(.a(\b[27] ), .b(\a[28] ), .out0(new_n311));
  inv040aa1d30x5               g216(.a(\a[27] ), .o1(new_n312));
  inv000aa1d42x5               g217(.a(\b[26] ), .o1(new_n313));
  aoi022aa1n02x5               g218(.a(new_n296), .b(new_n295), .c(new_n312), .d(new_n313), .o1(new_n314));
  nanp03aa1n03x5               g219(.a(new_n303), .b(new_n306), .c(new_n314), .o1(new_n315));
  oaib12aa1n06x5               g220(.a(new_n315), .b(new_n313), .c(\a[27] ), .out0(new_n316));
  oai022aa1n02x5               g221(.a(new_n312), .b(new_n313), .c(\b[27] ), .d(\a[28] ), .o1(new_n317));
  aoi012aa1n02x5               g222(.a(new_n317), .b(\a[28] ), .c(\b[27] ), .o1(new_n318));
  aoi022aa1n02x7               g223(.a(new_n316), .b(new_n311), .c(new_n315), .d(new_n318), .o1(\s[28] ));
  aoai13aa1n02x5               g224(.a(new_n307), .b(new_n301), .c(new_n287), .d(new_n283), .o1(new_n320));
  inv040aa1d32x5               g225(.a(\a[28] ), .o1(new_n321));
  xroi22aa1d06x4               g226(.a(new_n312), .b(\b[26] ), .c(new_n321), .d(\b[27] ), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n322), .b(new_n320), .c(new_n197), .d(new_n302), .o1(new_n323));
  inv000aa1n02x5               g228(.a(new_n322), .o1(new_n324));
  nanp02aa1n06x5               g229(.a(new_n313), .b(new_n312), .o1(new_n325));
  oao003aa1n03x5               g230(.a(\a[28] ), .b(\b[27] ), .c(new_n325), .carry(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n324), .c(new_n304), .d(new_n303), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .out0(new_n328));
  norb02aa1n02x5               g233(.a(new_n326), .b(new_n328), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n323), .d(new_n329), .o1(\s[29] ));
  xorb03aa1n02x5               g235(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g236(.a(new_n311), .b(new_n305), .c(new_n328), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n320), .c(new_n197), .d(new_n302), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n332), .o1(new_n334));
  oaoi03aa1n02x5               g239(.a(\a[29] ), .b(\b[28] ), .c(new_n326), .o1(new_n335));
  inv000aa1d42x5               g240(.a(new_n335), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n334), .c(new_n304), .d(new_n303), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[30] ), .b(\b[29] ), .out0(new_n338));
  aoi012aa1n02x5               g243(.a(new_n326), .b(\a[29] ), .c(\b[28] ), .o1(new_n339));
  oabi12aa1n02x5               g244(.a(new_n338), .b(\a[29] ), .c(\b[28] ), .out0(new_n340));
  norp02aa1n02x5               g245(.a(new_n339), .b(new_n340), .o1(new_n341));
  aoi022aa1n02x7               g246(.a(new_n337), .b(new_n338), .c(new_n333), .d(new_n341), .o1(\s[30] ));
  nano22aa1n02x5               g247(.a(new_n324), .b(new_n328), .c(new_n338), .out0(new_n343));
  aoai13aa1n02x5               g248(.a(new_n343), .b(new_n320), .c(new_n197), .d(new_n302), .o1(new_n344));
  inv000aa1d42x5               g249(.a(new_n343), .o1(new_n345));
  inv000aa1d42x5               g250(.a(\a[30] ), .o1(new_n346));
  inv000aa1d42x5               g251(.a(\b[29] ), .o1(new_n347));
  oaoi03aa1n02x5               g252(.a(new_n346), .b(new_n347), .c(new_n335), .o1(new_n348));
  aoai13aa1n03x5               g253(.a(new_n348), .b(new_n345), .c(new_n304), .d(new_n303), .o1(new_n349));
  xorc02aa1n02x5               g254(.a(\a[31] ), .b(\b[30] ), .out0(new_n350));
  oabi12aa1n02x5               g255(.a(new_n350), .b(\a[30] ), .c(\b[29] ), .out0(new_n351));
  oaoi13aa1n02x5               g256(.a(new_n351), .b(new_n335), .c(new_n346), .d(new_n347), .o1(new_n352));
  aoi022aa1n03x5               g257(.a(new_n349), .b(new_n350), .c(new_n344), .d(new_n352), .o1(\s[31] ));
  norb02aa1n02x5               g258(.a(new_n104), .b(new_n105), .out0(new_n354));
  xobna2aa1n03x5               g259(.a(new_n354), .b(new_n145), .c(new_n100), .out0(\s[3] ));
  aoai13aa1n02x5               g260(.a(new_n354), .b(new_n102), .c(\a[2] ), .d(\b[1] ), .o1(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n103), .b(new_n356), .c(new_n104), .out0(\s[4] ));
  norp02aa1n02x5               g262(.a(\b[4] ), .b(\a[5] ), .o1(new_n358));
  nanp02aa1n02x5               g263(.a(\b[4] ), .b(\a[5] ), .o1(new_n359));
  norb02aa1n02x5               g264(.a(new_n359), .b(new_n358), .out0(new_n360));
  nano23aa1n02x4               g265(.a(new_n107), .b(new_n358), .c(new_n108), .d(new_n359), .out0(new_n361));
  oai013aa1n02x4               g266(.a(new_n361), .b(new_n103), .c(new_n102), .d(new_n106), .o1(new_n362));
  aoai13aa1n02x5               g267(.a(new_n362), .b(new_n360), .c(new_n147), .d(new_n109), .o1(\s[5] ));
  xorc02aa1n02x5               g268(.a(\a[6] ), .b(\b[5] ), .out0(new_n364));
  xobna2aa1n03x5               g269(.a(new_n364), .b(new_n362), .c(new_n359), .out0(\s[6] ));
  aob012aa1n03x5               g270(.a(new_n364), .b(new_n362), .c(new_n359), .out0(new_n366));
  xorc02aa1n02x5               g271(.a(\a[7] ), .b(\b[6] ), .out0(new_n367));
  xobna2aa1n03x5               g272(.a(new_n367), .b(new_n366), .c(new_n112), .out0(\s[7] ));
  aob012aa1n02x5               g273(.a(new_n367), .b(new_n366), .c(new_n112), .out0(new_n369));
  aob012aa1n02x5               g274(.a(new_n369), .b(\b[6] ), .c(\a[7] ), .out0(new_n370));
  oa0012aa1n02x5               g275(.a(new_n121), .b(\b[7] ), .c(\a[8] ), .o(new_n371));
  aboi22aa1n03x5               g276(.a(new_n111), .b(new_n370), .c(new_n371), .d(new_n369), .out0(\s[8] ));
  oai112aa1n02x5               g277(.a(new_n118), .b(new_n124), .c(new_n122), .d(new_n119), .o1(new_n373));
  aboi22aa1n03x5               g278(.a(new_n373), .b(new_n153), .c(new_n150), .d(new_n125), .out0(\s[9] ));
endmodule


