// Benchmark "adder" written by ABC on Thu Jul 18 05:06:13 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n283, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n304, new_n305, new_n306, new_n308, new_n310, new_n312, new_n313,
    new_n314, new_n315, new_n317;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n04x5   g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\a[9] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\b[8] ), .b(new_n98), .out0(new_n99));
  oai022aa1n02x5               g004(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nand22aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  norb02aa1n06x5               g007(.a(new_n102), .b(new_n101), .out0(new_n103));
  nanp02aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oai112aa1n06x5               g009(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n105));
  aoi013aa1n09x5               g010(.a(new_n100), .b(new_n103), .c(new_n105), .d(new_n104), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor042aa1n04x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  norb03aa1n02x5               g014(.a(new_n107), .b(new_n109), .c(new_n108), .out0(new_n110));
  xorc02aa1n02x5               g015(.a(\a[6] ), .b(\b[5] ), .out0(new_n111));
  nanp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano32aa1n02x4               g020(.a(new_n114), .b(new_n115), .c(new_n112), .d(new_n113), .out0(new_n116));
  nanp03aa1n02x5               g021(.a(new_n116), .b(new_n110), .c(new_n111), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\a[6] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[5] ), .o1(new_n119));
  oao003aa1n02x5               g024(.a(new_n118), .b(new_n119), .c(new_n114), .carry(new_n120));
  nano23aa1n02x4               g025(.a(new_n109), .b(new_n108), .c(new_n112), .d(new_n107), .out0(new_n121));
  inv000aa1d42x5               g026(.a(new_n109), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  tech160nm_fiaoi012aa1n02p5x5 g028(.a(new_n123), .b(new_n121), .c(new_n120), .o1(new_n124));
  oai012aa1n12x5               g029(.a(new_n124), .b(new_n117), .c(new_n106), .o1(new_n125));
  oaib12aa1n06x5               g030(.a(new_n125), .b(new_n98), .c(\b[8] ), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  oai022aa1d24x5               g032(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  aoi022aa1n03x5               g034(.a(new_n126), .b(new_n129), .c(\b[9] ), .d(\a[10] ), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nanp02aa1n02x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norp02aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  aoi012aa1n03x5               g038(.a(new_n133), .b(new_n130), .c(new_n132), .o1(new_n134));
  xnrb03aa1n02x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv000aa1d42x5               g040(.a(\a[13] ), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanb02aa1n02x5               g042(.a(new_n133), .b(new_n132), .out0(new_n138));
  norp02aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n139), .b(new_n137), .out0(new_n140));
  xorc02aa1n02x5               g045(.a(\a[9] ), .b(\b[8] ), .out0(new_n141));
  nona23aa1n08x5               g046(.a(new_n97), .b(new_n141), .c(new_n140), .d(new_n138), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  norp02aa1n02x5               g048(.a(new_n139), .b(new_n133), .o1(new_n144));
  aoi022aa1n02x5               g049(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n145));
  aob012aa1n02x5               g050(.a(new_n144), .b(new_n128), .c(new_n145), .out0(new_n146));
  aoi022aa1n06x5               g051(.a(new_n125), .b(new_n143), .c(new_n137), .d(new_n146), .o1(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[12] ), .c(new_n136), .out0(\s[13] ));
  oaoi03aa1n02x5               g053(.a(\a[13] ), .b(\b[12] ), .c(new_n147), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xnrc02aa1n02x5               g055(.a(\b[12] ), .b(\a[13] ), .out0(new_n151));
  norp02aa1n02x5               g056(.a(\b[13] ), .b(\a[14] ), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nanb02aa1n02x5               g058(.a(new_n152), .b(new_n153), .out0(new_n154));
  norp02aa1n02x5               g059(.a(new_n151), .b(new_n154), .o1(new_n155));
  inv000aa1d42x5               g060(.a(\b[12] ), .o1(new_n156));
  aoai13aa1n02x5               g061(.a(new_n153), .b(new_n152), .c(new_n136), .d(new_n156), .o1(new_n157));
  oaib12aa1n06x5               g062(.a(new_n157), .b(new_n147), .c(new_n155), .out0(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv000aa1d42x5               g064(.a(\a[15] ), .o1(new_n160));
  inv000aa1d42x5               g065(.a(\b[14] ), .o1(new_n161));
  nand02aa1n04x5               g066(.a(new_n161), .b(new_n160), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nor002aa1n12x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n163), .c(new_n158), .d(new_n164), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n163), .b(new_n167), .c(new_n158), .d(new_n164), .o1(new_n169));
  nanb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(\s[16] ));
  nano22aa1n02x4               g075(.a(new_n167), .b(new_n162), .c(new_n164), .out0(new_n171));
  nano22aa1n12x5               g076(.a(new_n142), .b(new_n155), .c(new_n171), .out0(new_n172));
  nanp02aa1n02x5               g077(.a(new_n125), .b(new_n172), .o1(new_n173));
  oai012aa1n02x5               g078(.a(new_n137), .b(\b[12] ), .c(\a[13] ), .o1(new_n174));
  oai022aa1n02x5               g079(.a(new_n136), .b(new_n156), .c(\b[14] ), .d(\a[15] ), .o1(new_n175));
  norp03aa1n02x5               g080(.a(new_n154), .b(new_n174), .c(new_n175), .o1(new_n176));
  nano22aa1n02x4               g081(.a(new_n165), .b(new_n164), .c(new_n166), .out0(new_n177));
  nanp03aa1n02x5               g082(.a(new_n176), .b(new_n146), .c(new_n177), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n165), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(new_n166), .b(new_n164), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n179), .b(new_n180), .c(new_n157), .d(new_n162), .o1(new_n181));
  nanb02aa1n12x5               g086(.a(new_n181), .b(new_n178), .out0(new_n182));
  inv000aa1d42x5               g087(.a(new_n182), .o1(new_n183));
  xorc02aa1n02x5               g088(.a(\a[17] ), .b(\b[16] ), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n173), .c(new_n183), .out0(\s[17] ));
  orn002aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .o(new_n186));
  aoai13aa1n02x5               g091(.a(new_n184), .b(new_n182), .c(new_n125), .d(new_n172), .o1(new_n187));
  xorc02aa1n02x5               g092(.a(\a[18] ), .b(\b[17] ), .out0(new_n188));
  xnbna2aa1n03x5               g093(.a(new_n188), .b(new_n187), .c(new_n186), .out0(\s[18] ));
  norp02aa1n02x5               g094(.a(\b[17] ), .b(\a[18] ), .o1(new_n190));
  and002aa1n02x5               g095(.a(new_n188), .b(new_n184), .o(new_n191));
  aoai13aa1n02x5               g096(.a(new_n191), .b(new_n182), .c(new_n125), .d(new_n172), .o1(new_n192));
  aoi112aa1n03x5               g097(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n193));
  nona22aa1n03x5               g098(.a(new_n192), .b(new_n193), .c(new_n190), .out0(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n04x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nor042aa1n04x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1d16x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1n12x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  aoai13aa1n02x5               g107(.a(new_n202), .b(new_n197), .c(new_n194), .d(new_n198), .o1(new_n203));
  aoi112aa1n02x5               g108(.a(new_n197), .b(new_n202), .c(new_n194), .d(new_n198), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n204), .b(new_n203), .out0(\s[20] ));
  nano23aa1n02x4               g110(.a(new_n197), .b(new_n199), .c(new_n200), .d(new_n198), .out0(new_n206));
  nand03aa1n02x5               g111(.a(new_n206), .b(new_n184), .c(new_n188), .o1(new_n207));
  norb02aa1n06x4               g112(.a(new_n198), .b(new_n197), .out0(new_n208));
  oai112aa1n06x5               g113(.a(new_n208), .b(new_n201), .c(new_n193), .d(new_n190), .o1(new_n209));
  oai012aa1n02x7               g114(.a(new_n200), .b(new_n199), .c(new_n197), .o1(new_n210));
  nanp02aa1n02x5               g115(.a(new_n209), .b(new_n210), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n207), .c(new_n173), .d(new_n183), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  tech160nm_fixorc02aa1n02p5x5 g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  nor042aa1n04x5               g121(.a(\b[21] ), .b(\a[22] ), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(\b[21] ), .b(\a[22] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n215), .c(new_n213), .d(new_n216), .o1(new_n220));
  aoi112aa1n02x5               g125(.a(new_n215), .b(new_n219), .c(new_n213), .d(new_n216), .o1(new_n221));
  nanb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(\s[22] ));
  nanb02aa1n09x5               g127(.a(new_n219), .b(new_n216), .out0(new_n223));
  nano32aa1n02x4               g128(.a(new_n223), .b(new_n206), .c(new_n188), .d(new_n184), .out0(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n182), .c(new_n125), .d(new_n172), .o1(new_n225));
  oai012aa1n02x5               g130(.a(new_n218), .b(new_n217), .c(new_n215), .o1(new_n226));
  aoai13aa1n12x5               g131(.a(new_n226), .b(new_n223), .c(new_n209), .d(new_n210), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  xorc02aa1n02x5               g133(.a(\a[23] ), .b(\b[22] ), .out0(new_n229));
  xnbna2aa1n03x5               g134(.a(new_n229), .b(new_n225), .c(new_n228), .out0(\s[23] ));
  nand22aa1n03x5               g135(.a(new_n225), .b(new_n228), .o1(new_n231));
  norp02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[24] ), .b(\b[23] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n232), .c(new_n231), .d(new_n229), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n232), .b(new_n234), .c(new_n231), .d(new_n229), .o1(new_n236));
  nanb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(\s[24] ));
  inv000aa1d42x5               g142(.a(\a[23] ), .o1(new_n238));
  inv000aa1d42x5               g143(.a(\a[24] ), .o1(new_n239));
  xroi22aa1d04x5               g144(.a(new_n238), .b(\b[22] ), .c(new_n239), .d(\b[23] ), .out0(new_n240));
  norb03aa1n02x5               g145(.a(new_n240), .b(new_n207), .c(new_n223), .out0(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n182), .c(new_n125), .d(new_n172), .o1(new_n242));
  inv000aa1d42x5               g147(.a(\b[23] ), .o1(new_n243));
  oao003aa1n02x5               g148(.a(new_n239), .b(new_n243), .c(new_n232), .carry(new_n244));
  tech160nm_fiao0012aa1n02p5x5 g149(.a(new_n244), .b(new_n227), .c(new_n240), .o(new_n245));
  nanb02aa1n03x5               g150(.a(new_n245), .b(new_n242), .out0(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g152(.a(\b[24] ), .b(\a[25] ), .o1(new_n248));
  xorc02aa1n02x5               g153(.a(\a[25] ), .b(\b[24] ), .out0(new_n249));
  xorc02aa1n12x5               g154(.a(\a[26] ), .b(\b[25] ), .out0(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n248), .c(new_n246), .d(new_n249), .o1(new_n252));
  oaib12aa1n02x5               g157(.a(new_n249), .b(new_n245), .c(new_n242), .out0(new_n253));
  nona22aa1n02x4               g158(.a(new_n253), .b(new_n251), .c(new_n248), .out0(new_n254));
  nanp02aa1n03x5               g159(.a(new_n252), .b(new_n254), .o1(\s[26] ));
  norb02aa1n02x5               g160(.a(new_n216), .b(new_n219), .out0(new_n256));
  and002aa1n02x5               g161(.a(new_n250), .b(new_n249), .o(new_n257));
  nano32aa1n02x4               g162(.a(new_n207), .b(new_n257), .c(new_n256), .d(new_n240), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n182), .c(new_n125), .d(new_n172), .o1(new_n259));
  aoai13aa1n09x5               g164(.a(new_n257), .b(new_n244), .c(new_n227), .d(new_n240), .o1(new_n260));
  oai022aa1n02x5               g165(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n261));
  aob012aa1n02x5               g166(.a(new_n261), .b(\b[25] ), .c(\a[26] ), .out0(new_n262));
  nanp03aa1d12x5               g167(.a(new_n259), .b(new_n260), .c(new_n262), .o1(new_n263));
  xorb03aa1n02x5               g168(.a(new_n263), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n09x5               g169(.a(\b[26] ), .b(\a[27] ), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[27] ), .b(\b[26] ), .out0(new_n266));
  tech160nm_fixorc02aa1n02p5x5 g171(.a(\a[28] ), .b(\b[27] ), .out0(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n02x5               g173(.a(new_n268), .b(new_n265), .c(new_n263), .d(new_n266), .o1(new_n269));
  aoi112aa1n03x5               g174(.a(new_n265), .b(new_n268), .c(new_n263), .d(new_n266), .o1(new_n270));
  nanb02aa1n03x5               g175(.a(new_n270), .b(new_n269), .out0(\s[28] ));
  and002aa1n02x5               g176(.a(new_n267), .b(new_n266), .o(new_n272));
  nanp02aa1n03x5               g177(.a(new_n263), .b(new_n272), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\a[28] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(\b[27] ), .o1(new_n275));
  oaoi03aa1n12x5               g180(.a(new_n274), .b(new_n275), .c(new_n265), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[29] ), .b(\b[28] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  aoi012aa1n03x5               g183(.a(new_n278), .b(new_n273), .c(new_n276), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n276), .o1(new_n280));
  aoi112aa1n02x7               g185(.a(new_n277), .b(new_n280), .c(new_n263), .d(new_n272), .o1(new_n281));
  norp02aa1n03x5               g186(.a(new_n279), .b(new_n281), .o1(\s[29] ));
  nanp02aa1n02x5               g187(.a(\b[0] ), .b(\a[1] ), .o1(new_n283));
  xorb03aa1n02x5               g188(.a(new_n283), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xorc02aa1n02x5               g189(.a(\a[30] ), .b(\b[29] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  nano22aa1n02x4               g191(.a(new_n278), .b(new_n266), .c(new_n267), .out0(new_n287));
  nand02aa1n02x5               g192(.a(new_n263), .b(new_n287), .o1(new_n288));
  oao003aa1n09x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n276), .carry(new_n289));
  aoi012aa1n03x5               g194(.a(new_n286), .b(new_n288), .c(new_n289), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n289), .o1(new_n291));
  aoi112aa1n03x4               g196(.a(new_n285), .b(new_n291), .c(new_n263), .d(new_n287), .o1(new_n292));
  nor002aa1n02x5               g197(.a(new_n290), .b(new_n292), .o1(\s[30] ));
  xorc02aa1n02x5               g198(.a(\a[31] ), .b(\b[30] ), .out0(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  nano32aa1n02x4               g200(.a(new_n286), .b(new_n277), .c(new_n267), .d(new_n266), .out0(new_n296));
  nanp02aa1n02x5               g201(.a(new_n263), .b(new_n296), .o1(new_n297));
  tech160nm_fioaoi03aa1n03p5x5 g202(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n298), .o1(new_n299));
  aoi012aa1n03x5               g204(.a(new_n295), .b(new_n297), .c(new_n299), .o1(new_n300));
  aoi112aa1n03x4               g205(.a(new_n294), .b(new_n298), .c(new_n263), .d(new_n296), .o1(new_n301));
  nor002aa1n02x5               g206(.a(new_n300), .b(new_n301), .o1(\s[31] ));
  xobna2aa1n03x5               g207(.a(new_n103), .b(new_n105), .c(new_n104), .out0(\s[3] ));
  inv000aa1d42x5               g208(.a(new_n106), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[4] ), .b(\b[3] ), .out0(new_n305));
  aoi113aa1n02x5               g210(.a(new_n305), .b(new_n101), .c(new_n105), .d(new_n102), .e(new_n104), .o1(new_n306));
  aoi012aa1n02x5               g211(.a(new_n306), .b(new_n304), .c(new_n305), .o1(\s[4] ));
  norb02aa1n02x5               g212(.a(new_n115), .b(new_n114), .out0(new_n308));
  xobna2aa1n03x5               g213(.a(new_n308), .b(new_n304), .c(new_n113), .out0(\s[5] ));
  aoi013aa1n02x4               g214(.a(new_n114), .b(new_n304), .c(new_n113), .d(new_n115), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[5] ), .c(new_n118), .out0(\s[6] ));
  norb02aa1n02x5               g216(.a(new_n107), .b(new_n109), .out0(new_n312));
  nanp02aa1n02x5               g217(.a(new_n310), .b(new_n111), .o1(new_n313));
  oaoi13aa1n02x5               g218(.a(new_n312), .b(new_n313), .c(new_n118), .d(new_n119), .o1(new_n314));
  oai112aa1n02x5               g219(.a(new_n313), .b(new_n312), .c(new_n119), .d(new_n118), .o1(new_n315));
  norb02aa1n02x5               g220(.a(new_n315), .b(new_n314), .out0(\s[7] ));
  norb02aa1n02x5               g221(.a(new_n112), .b(new_n108), .out0(new_n317));
  xnbna2aa1n03x5               g222(.a(new_n317), .b(new_n315), .c(new_n122), .out0(\s[8] ));
  xorb03aa1n02x5               g223(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


