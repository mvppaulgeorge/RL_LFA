// Benchmark "adder" written by ABC on Thu Jul 18 00:02:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n308, new_n310,
    new_n311, new_n314, new_n315, new_n317, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  orn002aa1n02x5               g002(.a(\a[3] ), .b(\b[2] ), .o(new_n98));
  oao003aa1n02x5               g003(.a(\a[4] ), .b(\b[3] ), .c(new_n98), .carry(new_n99));
  tech160nm_fixorc02aa1n04x5   g004(.a(\a[4] ), .b(\b[3] ), .out0(new_n100));
  nand22aa1n06x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand42aa1n08x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  norp02aa1n06x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nona22aa1n03x5               g008(.a(new_n102), .b(new_n103), .c(new_n101), .out0(new_n104));
  nor042aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n10x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano22aa1n03x7               g011(.a(new_n105), .b(new_n102), .c(new_n106), .out0(new_n107));
  nanp03aa1d12x5               g012(.a(new_n104), .b(new_n107), .c(new_n100), .o1(new_n108));
  xnrc02aa1n12x5               g013(.a(\b[5] ), .b(\a[6] ), .out0(new_n109));
  xorc02aa1n12x5               g014(.a(\a[5] ), .b(\b[4] ), .out0(new_n110));
  xorc02aa1n12x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  nor022aa1n08x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  tech160nm_finand02aa1n05x5   g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanb02aa1n02x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  nona23aa1n09x5               g019(.a(new_n110), .b(new_n111), .c(new_n109), .d(new_n114), .out0(new_n115));
  nand42aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nano22aa1n02x5               g021(.a(new_n112), .b(new_n116), .c(new_n113), .out0(new_n117));
  oai022aa1n02x5               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  orn002aa1n02x5               g023(.a(\a[7] ), .b(\b[6] ), .o(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  aoi013aa1n06x4               g025(.a(new_n120), .b(new_n117), .c(new_n111), .d(new_n118), .o1(new_n121));
  aoai13aa1n12x5               g026(.a(new_n121), .b(new_n115), .c(new_n99), .d(new_n108), .o1(new_n122));
  tech160nm_fixorc02aa1n03p5x5 g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  tech160nm_fixorc02aa1n03p5x5 g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n125));
  aoi112aa1n02x5               g030(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n125), .b(new_n126), .out0(\s[10] ));
  norp02aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  tech160nm_fiaoi012aa1n04x5   g034(.a(new_n128), .b(new_n97), .c(new_n129), .o1(new_n130));
  xnrc02aa1n12x5               g035(.a(\b[10] ), .b(\a[11] ), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n125), .c(new_n130), .out0(\s[11] ));
  aob012aa1n03x5               g038(.a(new_n132), .b(new_n125), .c(new_n130), .out0(new_n134));
  xnrc02aa1n12x5               g039(.a(\b[11] ), .b(\a[12] ), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nor042aa1n06x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n135), .b(new_n137), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n137), .o1(new_n139));
  aoai13aa1n02x7               g044(.a(new_n139), .b(new_n131), .c(new_n125), .d(new_n130), .o1(new_n140));
  aoi022aa1n03x5               g045(.a(new_n140), .b(new_n136), .c(new_n134), .d(new_n138), .o1(\s[12] ));
  nano23aa1n06x5               g046(.a(new_n135), .b(new_n131), .c(new_n124), .d(new_n123), .out0(new_n142));
  nanp02aa1n02x5               g047(.a(new_n122), .b(new_n142), .o1(new_n143));
  oao003aa1n02x5               g048(.a(\a[12] ), .b(\b[11] ), .c(new_n139), .carry(new_n144));
  oai013aa1n02x4               g049(.a(new_n144), .b(new_n131), .c(new_n135), .d(new_n130), .o1(new_n145));
  nanb02aa1n02x5               g050(.a(new_n145), .b(new_n143), .out0(new_n146));
  xorb03aa1n02x5               g051(.a(new_n146), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g052(.a(\a[13] ), .o1(new_n148));
  nanb02aa1n12x5               g053(.a(\b[12] ), .b(new_n148), .out0(new_n149));
  xorc02aa1n02x5               g054(.a(\a[13] ), .b(\b[12] ), .out0(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n145), .c(new_n122), .d(new_n142), .o1(new_n151));
  xorc02aa1n02x5               g056(.a(\a[14] ), .b(\b[13] ), .out0(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n151), .c(new_n149), .out0(\s[14] ));
  inv000aa1d42x5               g058(.a(\a[14] ), .o1(new_n154));
  xroi22aa1d06x4               g059(.a(new_n148), .b(\b[12] ), .c(new_n154), .d(\b[13] ), .out0(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n145), .c(new_n122), .d(new_n142), .o1(new_n156));
  oaoi03aa1n12x5               g061(.a(\a[14] ), .b(\b[13] ), .c(new_n149), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  xorc02aa1n12x5               g063(.a(\a[15] ), .b(\b[14] ), .out0(new_n159));
  xnbna2aa1n03x5               g064(.a(new_n159), .b(new_n156), .c(new_n158), .out0(\s[15] ));
  aob012aa1n03x5               g065(.a(new_n159), .b(new_n156), .c(new_n158), .out0(new_n161));
  xorc02aa1n02x5               g066(.a(\a[16] ), .b(\b[15] ), .out0(new_n162));
  nor002aa1n06x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  norp02aa1n02x5               g068(.a(new_n162), .b(new_n163), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n163), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n159), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n165), .b(new_n166), .c(new_n156), .d(new_n158), .o1(new_n167));
  aoi022aa1n03x5               g072(.a(new_n167), .b(new_n162), .c(new_n161), .d(new_n164), .o1(\s[16] ));
  nor042aa1n02x5               g073(.a(new_n135), .b(new_n131), .o1(new_n169));
  and002aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .o(new_n170));
  xnrc02aa1n02x5               g075(.a(\b[15] ), .b(\a[16] ), .out0(new_n171));
  nona32aa1n02x4               g076(.a(new_n155), .b(new_n171), .c(new_n170), .d(new_n163), .out0(new_n172));
  nano32aa1n03x7               g077(.a(new_n172), .b(new_n169), .c(new_n124), .d(new_n123), .out0(new_n173));
  nand42aa1n04x5               g078(.a(new_n122), .b(new_n173), .o1(new_n174));
  nona22aa1n09x5               g079(.a(new_n136), .b(new_n131), .c(new_n130), .out0(new_n175));
  oaoi03aa1n02x5               g080(.a(\a[16] ), .b(\b[15] ), .c(new_n165), .o1(new_n176));
  aoi013aa1n06x4               g081(.a(new_n176), .b(new_n157), .c(new_n159), .d(new_n162), .o1(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n172), .c(new_n175), .d(new_n144), .o1(new_n178));
  nanb02aa1n06x5               g083(.a(new_n178), .b(new_n174), .out0(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g085(.a(\a[17] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\b[16] ), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(new_n182), .b(new_n181), .o1(new_n183));
  tech160nm_fixorc02aa1n02p5x5 g088(.a(\a[17] ), .b(\b[16] ), .out0(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n185));
  nor042aa1n02x5               g090(.a(\b[17] ), .b(\a[18] ), .o1(new_n186));
  nand22aa1n03x5               g091(.a(\b[17] ), .b(\a[18] ), .o1(new_n187));
  norb02aa1n06x5               g092(.a(new_n187), .b(new_n186), .out0(new_n188));
  xnbna2aa1n03x5               g093(.a(new_n188), .b(new_n185), .c(new_n183), .out0(\s[18] ));
  and002aa1n02x5               g094(.a(new_n184), .b(new_n188), .o(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n191));
  aoi013aa1n06x4               g096(.a(new_n186), .b(new_n187), .c(new_n181), .d(new_n182), .o1(new_n192));
  nor002aa1d32x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nand02aa1d04x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n191), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g102(.a(new_n195), .b(new_n191), .c(new_n192), .out0(new_n198));
  norp02aa1n12x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanp02aa1n06x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  norb02aa1n02x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  aoib12aa1n02x5               g106(.a(new_n193), .b(new_n200), .c(new_n199), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n193), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n195), .o1(new_n204));
  aoai13aa1n02x5               g109(.a(new_n203), .b(new_n204), .c(new_n191), .d(new_n192), .o1(new_n205));
  aoi022aa1n03x5               g110(.a(new_n205), .b(new_n201), .c(new_n198), .d(new_n202), .o1(\s[20] ));
  nano23aa1n06x5               g111(.a(new_n193), .b(new_n199), .c(new_n200), .d(new_n194), .out0(new_n207));
  nand23aa1n04x5               g112(.a(new_n207), .b(new_n184), .c(new_n188), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n210));
  nona23aa1n06x5               g115(.a(new_n200), .b(new_n194), .c(new_n193), .d(new_n199), .out0(new_n211));
  oaoi03aa1n09x5               g116(.a(\a[20] ), .b(\b[19] ), .c(new_n203), .o1(new_n212));
  oabi12aa1n12x5               g117(.a(new_n212), .b(new_n211), .c(new_n192), .out0(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  xnrc02aa1n12x5               g119(.a(\b[20] ), .b(\a[21] ), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n210), .c(new_n214), .out0(\s[21] ));
  aob012aa1n03x5               g122(.a(new_n216), .b(new_n210), .c(new_n214), .out0(new_n218));
  tech160nm_fixnrc02aa1n04x5   g123(.a(\b[21] ), .b(\a[22] ), .out0(new_n219));
  nor042aa1n03x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  norb02aa1n02x5               g125(.a(new_n219), .b(new_n220), .out0(new_n221));
  inv000aa1n03x5               g126(.a(new_n220), .o1(new_n222));
  aoai13aa1n02x5               g127(.a(new_n222), .b(new_n215), .c(new_n210), .d(new_n214), .o1(new_n223));
  aboi22aa1n03x5               g128(.a(new_n219), .b(new_n223), .c(new_n218), .d(new_n221), .out0(\s[22] ));
  nor042aa1n06x5               g129(.a(new_n219), .b(new_n215), .o1(new_n225));
  norb02aa1n03x5               g130(.a(new_n225), .b(new_n208), .out0(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n227));
  oaoi03aa1n02x5               g132(.a(\a[22] ), .b(\b[21] ), .c(new_n222), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n213), .c(new_n225), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[22] ), .b(\a[23] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  xnbna2aa1n03x5               g136(.a(new_n231), .b(new_n227), .c(new_n229), .out0(\s[23] ));
  aob012aa1n03x5               g137(.a(new_n231), .b(new_n227), .c(new_n229), .out0(new_n233));
  xorc02aa1n12x5               g138(.a(\a[24] ), .b(\b[23] ), .out0(new_n234));
  nor042aa1n06x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  norp02aa1n02x5               g140(.a(new_n234), .b(new_n235), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n235), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n230), .c(new_n227), .d(new_n229), .o1(new_n238));
  aoi022aa1n02x5               g143(.a(new_n238), .b(new_n234), .c(new_n233), .d(new_n236), .o1(\s[24] ));
  nano32aa1n02x5               g144(.a(new_n208), .b(new_n234), .c(new_n225), .d(new_n231), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[18] ), .b(\b[17] ), .c(new_n183), .o1(new_n242));
  aoai13aa1n06x5               g147(.a(new_n225), .b(new_n212), .c(new_n207), .d(new_n242), .o1(new_n243));
  inv000aa1n02x5               g148(.a(new_n228), .o1(new_n244));
  norb02aa1n06x4               g149(.a(new_n234), .b(new_n230), .out0(new_n245));
  inv000aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  oao003aa1n02x5               g151(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .carry(new_n247));
  aoai13aa1n12x5               g152(.a(new_n247), .b(new_n246), .c(new_n243), .d(new_n244), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[25] ), .b(\b[24] ), .out0(new_n250));
  xnbna2aa1n03x5               g155(.a(new_n250), .b(new_n241), .c(new_n249), .out0(\s[25] ));
  aob012aa1n03x5               g156(.a(new_n250), .b(new_n241), .c(new_n249), .out0(new_n252));
  tech160nm_fixorc02aa1n02p5x5 g157(.a(\a[26] ), .b(\b[25] ), .out0(new_n253));
  norp02aa1n02x5               g158(.a(\b[24] ), .b(\a[25] ), .o1(new_n254));
  norp02aa1n02x5               g159(.a(new_n253), .b(new_n254), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n254), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n250), .o1(new_n257));
  aoai13aa1n02x5               g162(.a(new_n256), .b(new_n257), .c(new_n241), .d(new_n249), .o1(new_n258));
  aoi022aa1n02x7               g163(.a(new_n258), .b(new_n253), .c(new_n252), .d(new_n255), .o1(\s[26] ));
  and002aa1n12x5               g164(.a(new_n253), .b(new_n250), .o(new_n260));
  nano32aa1n03x7               g165(.a(new_n208), .b(new_n260), .c(new_n225), .d(new_n245), .out0(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n178), .c(new_n122), .d(new_n173), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(\b[25] ), .b(\a[26] ), .o1(new_n263));
  oai022aa1n02x5               g168(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n264));
  aoi022aa1n12x5               g169(.a(new_n248), .b(new_n260), .c(new_n263), .d(new_n264), .o1(new_n265));
  xorc02aa1n12x5               g170(.a(\a[27] ), .b(\b[26] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n265), .c(new_n262), .out0(\s[27] ));
  aoai13aa1n03x5               g172(.a(new_n245), .b(new_n228), .c(new_n213), .d(new_n225), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n260), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(new_n264), .b(new_n263), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n269), .c(new_n268), .d(new_n247), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n266), .b(new_n271), .c(new_n179), .d(new_n261), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[28] ), .b(\b[27] ), .out0(new_n273));
  norp02aa1n02x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  norp02aa1n02x5               g179(.a(new_n273), .b(new_n274), .o1(new_n275));
  inv000aa1n03x5               g180(.a(new_n274), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n266), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n276), .b(new_n277), .c(new_n265), .d(new_n262), .o1(new_n278));
  aoi022aa1n03x5               g183(.a(new_n278), .b(new_n273), .c(new_n272), .d(new_n275), .o1(\s[28] ));
  and002aa1n02x5               g184(.a(new_n273), .b(new_n266), .o(new_n280));
  aoai13aa1n02x5               g185(.a(new_n280), .b(new_n271), .c(new_n179), .d(new_n261), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n280), .o1(new_n282));
  oao003aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n276), .carry(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n282), .c(new_n265), .d(new_n262), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[29] ), .b(\b[28] ), .out0(new_n285));
  norb02aa1n02x5               g190(.a(new_n283), .b(new_n285), .out0(new_n286));
  aoi022aa1n03x5               g191(.a(new_n284), .b(new_n285), .c(new_n281), .d(new_n286), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g193(.a(new_n277), .b(new_n273), .c(new_n285), .out0(new_n289));
  aoai13aa1n02x5               g194(.a(new_n289), .b(new_n271), .c(new_n179), .d(new_n261), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n289), .o1(new_n291));
  oaoi03aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .c(new_n283), .o1(new_n292));
  inv000aa1n03x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n291), .c(new_n265), .d(new_n262), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[30] ), .b(\b[29] ), .out0(new_n295));
  and002aa1n02x5               g200(.a(\b[28] ), .b(\a[29] ), .o(new_n296));
  oabi12aa1n02x5               g201(.a(new_n295), .b(\a[29] ), .c(\b[28] ), .out0(new_n297));
  oab012aa1n02x4               g202(.a(new_n297), .b(new_n283), .c(new_n296), .out0(new_n298));
  aoi022aa1n03x5               g203(.a(new_n294), .b(new_n295), .c(new_n290), .d(new_n298), .o1(\s[30] ));
  nano32aa1n06x5               g204(.a(new_n277), .b(new_n295), .c(new_n273), .d(new_n285), .out0(new_n300));
  aoai13aa1n02x5               g205(.a(new_n300), .b(new_n271), .c(new_n179), .d(new_n261), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[31] ), .b(\b[30] ), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n303));
  norb02aa1n02x5               g208(.a(new_n303), .b(new_n302), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n300), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n303), .b(new_n305), .c(new_n265), .d(new_n262), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[31] ));
  norb02aa1n02x5               g212(.a(new_n106), .b(new_n105), .out0(new_n308));
  xobna2aa1n03x5               g213(.a(new_n308), .b(new_n104), .c(new_n102), .out0(\s[3] ));
  nanp02aa1n02x5               g214(.a(new_n108), .b(new_n99), .o1(new_n310));
  aoi112aa1n02x5               g215(.a(new_n105), .b(new_n100), .c(new_n107), .d(new_n104), .o1(new_n311));
  oaoi13aa1n02x5               g216(.a(new_n311), .b(new_n310), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g217(.a(new_n110), .b(new_n108), .c(new_n99), .out0(\s[5] ));
  nanp02aa1n02x5               g218(.a(new_n310), .b(new_n110), .o1(new_n314));
  oai012aa1n02x5               g219(.a(new_n314), .b(\b[4] ), .c(\a[5] ), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oai012aa1n02x5               g221(.a(new_n117), .b(new_n315), .c(new_n109), .o1(new_n317));
  oai012aa1n02x5               g222(.a(new_n116), .b(new_n315), .c(new_n109), .o1(new_n318));
  aobi12aa1n02x5               g223(.a(new_n317), .b(new_n318), .c(new_n114), .out0(\s[7] ));
  xnbna2aa1n03x5               g224(.a(new_n111), .b(new_n317), .c(new_n119), .out0(\s[8] ));
  xorb03aa1n02x5               g225(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


