// Benchmark "adder" written by ABC on Thu Jul 18 07:19:07 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n326, new_n328, new_n329, new_n331, new_n333,
    new_n334, new_n335, new_n337, new_n338, new_n340, new_n341, new_n342,
    new_n344, new_n345, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1n03x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nona22aa1n03x5               g005(.a(new_n99), .b(new_n98), .c(new_n100), .out0(new_n101));
  aoi022aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .c(\a[2] ), .d(\b[1] ), .o1(new_n102));
  nor002aa1n06x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n08x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb03aa1n12x5               g010(.a(new_n105), .b(new_n103), .c(new_n104), .out0(new_n106));
  nanp03aa1n06x5               g011(.a(new_n101), .b(new_n106), .c(new_n102), .o1(new_n107));
  tech160nm_fioai012aa1n03p5x5 g012(.a(new_n105), .b(new_n104), .c(new_n103), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1n06x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor002aa1n03x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nanp02aa1n09x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nano23aa1n03x5               g017(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n113));
  tech160nm_fixorc02aa1n02p5x5 g018(.a(\a[8] ), .b(\b[7] ), .out0(new_n114));
  xorc02aa1n02x5               g019(.a(\a[6] ), .b(\b[5] ), .out0(new_n115));
  nand23aa1n03x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  norp02aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  aoi112aa1n03x5               g022(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n118));
  oai022aa1n04x5               g023(.a(\a[6] ), .b(\b[5] ), .c(\b[6] ), .d(\a[7] ), .o1(new_n119));
  aoi022aa1n02x5               g024(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n120));
  oaoi13aa1n09x5               g025(.a(new_n117), .b(new_n120), .c(new_n118), .d(new_n119), .o1(new_n121));
  aoai13aa1n12x5               g026(.a(new_n121), .b(new_n116), .c(new_n107), .d(new_n108), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  xorc02aa1n12x5               g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  aoai13aa1n09x5               g029(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n125));
  aoi112aa1n02x5               g030(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n125), .b(new_n126), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(\a[10] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(\b[9] ), .o1(new_n129));
  oao003aa1n09x5               g034(.a(new_n128), .b(new_n129), .c(new_n97), .carry(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  nor042aa1n09x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n125), .c(new_n131), .out0(\s[11] ));
  aob012aa1n03x5               g040(.a(new_n134), .b(new_n125), .c(new_n131), .out0(new_n136));
  inv000aa1d42x5               g041(.a(new_n132), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n134), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n137), .b(new_n138), .c(new_n125), .d(new_n131), .o1(new_n139));
  nor042aa1n02x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  aoib12aa1n02x5               g047(.a(new_n132), .b(new_n141), .c(new_n140), .out0(new_n143));
  aoi022aa1n03x5               g048(.a(new_n139), .b(new_n142), .c(new_n136), .d(new_n143), .o1(\s[12] ));
  nano23aa1n06x5               g049(.a(new_n132), .b(new_n140), .c(new_n141), .d(new_n133), .out0(new_n145));
  nand23aa1n06x5               g050(.a(new_n145), .b(new_n123), .c(new_n124), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  tech160nm_finand02aa1n03p5x5 g052(.a(new_n145), .b(new_n130), .o1(new_n148));
  aoi012aa1n09x5               g053(.a(new_n140), .b(new_n132), .c(new_n141), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n148), .b(new_n149), .o1(new_n150));
  xnrc02aa1n12x5               g055(.a(\b[12] ), .b(\a[13] ), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n06x5               g057(.a(new_n152), .b(new_n150), .c(new_n122), .d(new_n147), .o1(new_n153));
  and003aa1n02x5               g058(.a(new_n148), .b(new_n151), .c(new_n149), .o(new_n154));
  aobi12aa1n02x5               g059(.a(new_n154), .b(new_n147), .c(new_n122), .out0(new_n155));
  norb02aa1n02x5               g060(.a(new_n153), .b(new_n155), .out0(\s[13] ));
  orn002aa1n24x5               g061(.a(\a[13] ), .b(\b[12] ), .o(new_n157));
  tech160nm_fixnrc02aa1n04x5   g062(.a(\b[13] ), .b(\a[14] ), .out0(new_n158));
  xobna2aa1n03x5               g063(.a(new_n158), .b(new_n153), .c(new_n157), .out0(\s[14] ));
  nor022aa1n04x5               g064(.a(new_n158), .b(new_n151), .o1(new_n160));
  aoai13aa1n06x5               g065(.a(new_n160), .b(new_n150), .c(new_n122), .d(new_n147), .o1(new_n161));
  oaoi03aa1n12x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  tech160nm_fixorc02aa1n02p5x5 g068(.a(\a[15] ), .b(\b[14] ), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n161), .c(new_n163), .out0(\s[15] ));
  aob012aa1n03x5               g070(.a(new_n164), .b(new_n161), .c(new_n163), .out0(new_n166));
  nor042aa1n06x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  xnrc02aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n168), .b(new_n169), .c(new_n161), .d(new_n163), .o1(new_n170));
  xorc02aa1n02x5               g075(.a(\a[16] ), .b(\b[15] ), .out0(new_n171));
  norp02aa1n02x5               g076(.a(new_n171), .b(new_n167), .o1(new_n172));
  aoi022aa1n02x5               g077(.a(new_n170), .b(new_n171), .c(new_n166), .d(new_n172), .o1(\s[16] ));
  xnrc02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .out0(new_n174));
  norp02aa1n02x5               g079(.a(new_n174), .b(new_n169), .o1(new_n175));
  nano22aa1n12x5               g080(.a(new_n146), .b(new_n160), .c(new_n175), .out0(new_n176));
  nanp02aa1n09x5               g081(.a(new_n122), .b(new_n176), .o1(new_n177));
  nand22aa1n03x5               g082(.a(new_n175), .b(new_n160), .o1(new_n178));
  oaoi03aa1n02x5               g083(.a(\a[16] ), .b(\b[15] ), .c(new_n168), .o1(new_n179));
  aoi013aa1n06x5               g084(.a(new_n179), .b(new_n162), .c(new_n164), .d(new_n171), .o1(new_n180));
  aoai13aa1n12x5               g085(.a(new_n180), .b(new_n178), .c(new_n148), .d(new_n149), .o1(new_n181));
  nanb02aa1n12x5               g086(.a(new_n181), .b(new_n177), .out0(new_n182));
  xorc02aa1n02x5               g087(.a(\a[17] ), .b(\b[16] ), .out0(new_n183));
  aoi113aa1n02x5               g088(.a(new_n179), .b(new_n183), .c(new_n162), .d(new_n164), .e(new_n171), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n178), .c(new_n148), .d(new_n149), .o1(new_n185));
  aboi22aa1n03x5               g090(.a(new_n185), .b(new_n177), .c(new_n182), .d(new_n183), .out0(\s[17] ));
  nor042aa1n09x5               g091(.a(\b[16] ), .b(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n183), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n189));
  nor042aa1n02x5               g094(.a(\b[17] ), .b(\a[18] ), .o1(new_n190));
  nand02aa1n03x5               g095(.a(\b[17] ), .b(\a[18] ), .o1(new_n191));
  norb02aa1n03x5               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n192), .b(new_n189), .c(new_n188), .out0(\s[18] ));
  and002aa1n02x5               g098(.a(new_n183), .b(new_n192), .o(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n195));
  oaoi03aa1n02x5               g100(.a(\a[18] ), .b(\b[17] ), .c(new_n188), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  tech160nm_fixorc02aa1n05x5   g102(.a(\a[19] ), .b(\b[18] ), .out0(new_n198));
  xnbna2aa1n03x5               g103(.a(new_n198), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g105(.a(new_n198), .b(new_n195), .c(new_n197), .out0(new_n201));
  inv000aa1d42x5               g106(.a(\a[19] ), .o1(new_n202));
  inv000aa1d42x5               g107(.a(\b[18] ), .o1(new_n203));
  nand02aa1d12x5               g108(.a(new_n203), .b(new_n202), .o1(new_n204));
  inv030aa1n02x5               g109(.a(new_n198), .o1(new_n205));
  aoai13aa1n02x5               g110(.a(new_n204), .b(new_n205), .c(new_n195), .d(new_n197), .o1(new_n206));
  nor002aa1n02x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nanp02aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  aboi22aa1n03x5               g114(.a(new_n207), .b(new_n208), .c(new_n202), .d(new_n203), .out0(new_n210));
  aoi022aa1n02x5               g115(.a(new_n206), .b(new_n209), .c(new_n201), .d(new_n210), .o1(\s[20] ));
  nano32aa1n03x7               g116(.a(new_n205), .b(new_n183), .c(new_n209), .d(new_n192), .out0(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n213));
  oaoi03aa1n03x5               g118(.a(\a[20] ), .b(\b[19] ), .c(new_n204), .o1(new_n214));
  inv030aa1n02x5               g119(.a(new_n214), .o1(new_n215));
  nanp02aa1n02x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  nanb03aa1n06x5               g121(.a(new_n207), .b(new_n208), .c(new_n216), .out0(new_n217));
  oai112aa1n06x5               g122(.a(new_n191), .b(new_n204), .c(new_n190), .d(new_n187), .o1(new_n218));
  oai012aa1n18x5               g123(.a(new_n215), .b(new_n218), .c(new_n217), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  nor042aa1n12x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  nanp02aa1n03x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1d27x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  aob012aa1n03x5               g128(.a(new_n223), .b(new_n213), .c(new_n220), .out0(new_n224));
  nano22aa1n03x5               g129(.a(new_n207), .b(new_n216), .c(new_n208), .out0(new_n225));
  oai012aa1n02x5               g130(.a(new_n191), .b(\b[18] ), .c(\a[19] ), .o1(new_n226));
  oab012aa1n02x5               g131(.a(new_n226), .b(new_n187), .c(new_n190), .out0(new_n227));
  aoi112aa1n02x5               g132(.a(new_n223), .b(new_n214), .c(new_n227), .d(new_n225), .o1(new_n228));
  aobi12aa1n02x7               g133(.a(new_n224), .b(new_n228), .c(new_n213), .out0(\s[21] ));
  inv000aa1d42x5               g134(.a(new_n221), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n223), .o1(new_n231));
  aoai13aa1n02x5               g136(.a(new_n230), .b(new_n231), .c(new_n213), .d(new_n220), .o1(new_n232));
  nor042aa1n03x5               g137(.a(\b[21] ), .b(\a[22] ), .o1(new_n233));
  nand22aa1n04x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  aoib12aa1n02x5               g140(.a(new_n221), .b(new_n234), .c(new_n233), .out0(new_n236));
  aoi022aa1n02x5               g141(.a(new_n232), .b(new_n235), .c(new_n224), .d(new_n236), .o1(\s[22] ));
  inv000aa1n02x5               g142(.a(new_n212), .o1(new_n238));
  nano22aa1n03x7               g143(.a(new_n238), .b(new_n223), .c(new_n235), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n240));
  nano23aa1n06x5               g145(.a(new_n221), .b(new_n233), .c(new_n234), .d(new_n222), .out0(new_n241));
  aoi012aa1d18x5               g146(.a(new_n233), .b(new_n221), .c(new_n234), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n243), .b(new_n219), .c(new_n241), .o1(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  aob012aa1n03x5               g150(.a(new_n245), .b(new_n240), .c(new_n244), .out0(new_n246));
  aoi112aa1n02x5               g151(.a(new_n245), .b(new_n243), .c(new_n219), .d(new_n241), .o1(new_n247));
  aobi12aa1n02x7               g152(.a(new_n246), .b(new_n247), .c(new_n240), .out0(\s[23] ));
  nor042aa1n06x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n245), .o1(new_n251));
  aoai13aa1n02x5               g156(.a(new_n250), .b(new_n251), .c(new_n240), .d(new_n244), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .out0(new_n253));
  norp02aa1n02x5               g158(.a(new_n253), .b(new_n249), .o1(new_n254));
  aoi022aa1n03x5               g159(.a(new_n252), .b(new_n253), .c(new_n246), .d(new_n254), .o1(\s[24] ));
  and002aa1n02x7               g160(.a(new_n253), .b(new_n245), .o(new_n256));
  nano22aa1n02x4               g161(.a(new_n238), .b(new_n256), .c(new_n241), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n258));
  aoai13aa1n06x5               g163(.a(new_n241), .b(new_n214), .c(new_n227), .d(new_n225), .o1(new_n259));
  inv000aa1n03x5               g164(.a(new_n256), .o1(new_n260));
  oao003aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .c(new_n250), .carry(new_n261));
  aoai13aa1n12x5               g166(.a(new_n261), .b(new_n260), .c(new_n259), .d(new_n242), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  aob012aa1n03x5               g169(.a(new_n264), .b(new_n258), .c(new_n263), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n256), .b(new_n243), .c(new_n219), .d(new_n241), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n264), .o1(new_n267));
  and003aa1n02x5               g172(.a(new_n266), .b(new_n267), .c(new_n261), .o(new_n268));
  aobi12aa1n02x7               g173(.a(new_n265), .b(new_n268), .c(new_n258), .out0(\s[25] ));
  nor042aa1n03x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n271), .b(new_n267), .c(new_n258), .d(new_n263), .o1(new_n272));
  tech160nm_fixorc02aa1n03p5x5 g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  norp02aa1n02x5               g178(.a(new_n273), .b(new_n270), .o1(new_n274));
  aoi022aa1n03x5               g179(.a(new_n272), .b(new_n273), .c(new_n265), .d(new_n274), .o1(\s[26] ));
  and002aa1n18x5               g180(.a(new_n273), .b(new_n264), .o(new_n276));
  nano32aa1n03x7               g181(.a(new_n238), .b(new_n276), .c(new_n241), .d(new_n256), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n181), .c(new_n122), .d(new_n176), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n276), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n279), .c(new_n266), .d(new_n261), .o1(new_n281));
  xorc02aa1n02x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n281), .c(new_n182), .d(new_n277), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n280), .o1(new_n284));
  aoi112aa1n02x5               g189(.a(new_n282), .b(new_n284), .c(new_n262), .d(new_n276), .o1(new_n285));
  aobi12aa1n02x7               g190(.a(new_n283), .b(new_n285), .c(new_n278), .out0(\s[27] ));
  tech160nm_fiaoi012aa1n05x5   g191(.a(new_n284), .b(new_n262), .c(new_n276), .o1(new_n287));
  nor042aa1d18x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv000aa1n06x5               g193(.a(new_n288), .o1(new_n289));
  inv000aa1n02x5               g194(.a(new_n282), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n289), .b(new_n290), .c(new_n287), .d(new_n278), .o1(new_n291));
  xorc02aa1n12x5               g196(.a(\a[28] ), .b(\b[27] ), .out0(new_n292));
  norp02aa1n02x5               g197(.a(new_n292), .b(new_n288), .o1(new_n293));
  aoi022aa1n03x5               g198(.a(new_n291), .b(new_n292), .c(new_n283), .d(new_n293), .o1(\s[28] ));
  and002aa1n02x5               g199(.a(new_n292), .b(new_n282), .o(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n281), .c(new_n182), .d(new_n277), .o1(new_n296));
  inv000aa1n02x5               g201(.a(new_n295), .o1(new_n297));
  oao003aa1n03x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n297), .c(new_n287), .d(new_n278), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n298), .b(new_n300), .out0(new_n301));
  aoi022aa1n03x5               g206(.a(new_n299), .b(new_n300), .c(new_n296), .d(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d33x5               g208(.a(new_n290), .b(new_n292), .c(new_n300), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n281), .c(new_n182), .d(new_n277), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n304), .o1(new_n306));
  tech160nm_fioaoi03aa1n02p5x5 g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n306), .c(new_n287), .d(new_n278), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .out0(new_n310));
  and002aa1n02x5               g215(.a(\b[28] ), .b(\a[29] ), .o(new_n311));
  oabi12aa1n02x5               g216(.a(new_n310), .b(\a[29] ), .c(\b[28] ), .out0(new_n312));
  oab012aa1n02x4               g217(.a(new_n312), .b(new_n298), .c(new_n311), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n309), .b(new_n310), .c(new_n305), .d(new_n313), .o1(\s[30] ));
  nano32aa1d15x5               g219(.a(new_n290), .b(new_n310), .c(new_n292), .d(new_n300), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n281), .c(new_n182), .d(new_n277), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[31] ), .b(\b[30] ), .out0(new_n317));
  inv000aa1d42x5               g222(.a(\a[30] ), .o1(new_n318));
  inv000aa1d42x5               g223(.a(\b[29] ), .o1(new_n319));
  oabi12aa1n02x5               g224(.a(new_n317), .b(\a[30] ), .c(\b[29] ), .out0(new_n320));
  oaoi13aa1n02x5               g225(.a(new_n320), .b(new_n307), .c(new_n318), .d(new_n319), .o1(new_n321));
  inv000aa1d42x5               g226(.a(new_n315), .o1(new_n322));
  oaoi03aa1n02x5               g227(.a(new_n318), .b(new_n319), .c(new_n307), .o1(new_n323));
  aoai13aa1n03x5               g228(.a(new_n323), .b(new_n322), .c(new_n287), .d(new_n278), .o1(new_n324));
  aoi022aa1n03x5               g229(.a(new_n324), .b(new_n317), .c(new_n316), .d(new_n321), .o1(\s[31] ));
  xorc02aa1n02x5               g230(.a(\a[3] ), .b(\b[2] ), .out0(new_n326));
  xobna2aa1n03x5               g231(.a(new_n326), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  aob012aa1n02x5               g232(.a(new_n326), .b(new_n101), .c(new_n99), .out0(new_n328));
  aboi22aa1n03x5               g233(.a(new_n103), .b(new_n105), .c(\a[3] ), .d(\b[2] ), .out0(new_n329));
  ao0022aa1n03x5               g234(.a(new_n328), .b(new_n329), .c(new_n107), .d(new_n106), .o(\s[4] ));
  norb02aa1n02x5               g235(.a(new_n112), .b(new_n111), .out0(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n331), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  nanp02aa1n02x5               g237(.a(new_n107), .b(new_n108), .o1(new_n333));
  aoai13aa1n02x5               g238(.a(new_n115), .b(new_n111), .c(new_n333), .d(new_n112), .o1(new_n334));
  aoi112aa1n02x5               g239(.a(new_n111), .b(new_n115), .c(new_n333), .d(new_n331), .o1(new_n335));
  norb02aa1n02x5               g240(.a(new_n334), .b(new_n335), .out0(\s[6] ));
  norb02aa1n02x5               g241(.a(new_n110), .b(new_n109), .out0(new_n337));
  oab012aa1n02x4               g242(.a(new_n118), .b(\a[6] ), .c(\b[5] ), .out0(new_n338));
  xnbna2aa1n03x5               g243(.a(new_n337), .b(new_n334), .c(new_n338), .out0(\s[7] ));
  aob012aa1n02x5               g244(.a(new_n337), .b(new_n334), .c(new_n338), .out0(new_n340));
  oai012aa1n02x5               g245(.a(new_n340), .b(\b[6] ), .c(\a[7] ), .o1(new_n341));
  norp02aa1n02x5               g246(.a(new_n114), .b(new_n109), .o1(new_n342));
  aoi022aa1n02x5               g247(.a(new_n341), .b(new_n114), .c(new_n340), .d(new_n342), .o1(\s[8] ));
  nanb02aa1n02x5               g248(.a(new_n116), .b(new_n333), .out0(new_n344));
  oai012aa1n02x5               g249(.a(new_n120), .b(new_n118), .c(new_n119), .o1(new_n345));
  norb03aa1n02x5               g250(.a(new_n345), .b(new_n117), .c(new_n123), .out0(new_n346));
  aoi022aa1n02x5               g251(.a(new_n122), .b(new_n123), .c(new_n344), .d(new_n346), .o1(\s[9] ));
endmodule


