// Benchmark "adder" written by ABC on Thu Jul 18 03:08:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n332, new_n334, new_n335, new_n337, new_n339, new_n341,
    new_n342, new_n343, new_n346, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oao003aa1n02x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n101));
  nand42aa1n06x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor042aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  tech160nm_finand02aa1n03p5x5 g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano23aa1n02x4               g010(.a(new_n104), .b(new_n103), .c(new_n105), .d(new_n102), .out0(new_n106));
  tech160nm_fiaoi012aa1n03p5x5 g011(.a(new_n103), .b(new_n104), .c(new_n102), .o1(new_n107));
  aobi12aa1n02x7               g012(.a(new_n107), .b(new_n106), .c(new_n101), .out0(new_n108));
  xnrc02aa1n12x5               g013(.a(\b[5] ), .b(\a[6] ), .out0(new_n109));
  xnrc02aa1n12x5               g014(.a(\b[4] ), .b(\a[5] ), .out0(new_n110));
  inv000aa1d42x5               g015(.a(new_n110), .o1(new_n111));
  nor022aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanb02aa1n03x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  nanp02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nor002aa1d32x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  inv030aa1n02x5               g022(.a(new_n117), .o1(new_n118));
  nona23aa1n09x5               g023(.a(new_n111), .b(new_n118), .c(new_n109), .d(new_n114), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\a[6] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[5] ), .o1(new_n121));
  nor002aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(new_n120), .b(new_n121), .c(new_n122), .o1(new_n123));
  nona23aa1n02x4               g028(.a(new_n115), .b(new_n113), .c(new_n116), .d(new_n112), .out0(new_n124));
  inv000aa1d42x5               g029(.a(new_n116), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[8] ), .b(\b[7] ), .c(new_n125), .o1(new_n126));
  oabi12aa1n06x5               g031(.a(new_n126), .b(new_n124), .c(new_n123), .out0(new_n127));
  oabi12aa1n09x5               g032(.a(new_n127), .b(new_n108), .c(new_n119), .out0(new_n128));
  nand42aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  aoi012aa1n02x5               g034(.a(new_n97), .b(new_n128), .c(new_n129), .o1(new_n130));
  xnrb03aa1n02x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  oaoi03aa1n09x5               g036(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n132));
  nona23aa1n09x5               g037(.a(new_n102), .b(new_n105), .c(new_n104), .d(new_n103), .out0(new_n133));
  oai012aa1n06x5               g038(.a(new_n107), .b(new_n133), .c(new_n132), .o1(new_n134));
  nona23aa1n02x4               g039(.a(new_n115), .b(new_n113), .c(new_n116), .d(new_n112), .out0(new_n135));
  nor043aa1n03x5               g040(.a(new_n135), .b(new_n110), .c(new_n109), .o1(new_n136));
  nor042aa1n06x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nand22aa1n12x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  nano23aa1n06x5               g043(.a(new_n137), .b(new_n97), .c(new_n129), .d(new_n138), .out0(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n127), .c(new_n134), .d(new_n136), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n137), .b(new_n97), .c(new_n138), .o1(new_n141));
  nor022aa1n08x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand02aa1n06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n144), .b(new_n140), .c(new_n141), .out0(\s[11] ));
  inv030aa1n02x5               g050(.a(new_n142), .o1(new_n146));
  aob012aa1n02x5               g051(.a(new_n144), .b(new_n140), .c(new_n141), .out0(new_n147));
  norp02aa1n12x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nand42aa1n03x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nanb02aa1n02x5               g054(.a(new_n148), .b(new_n149), .out0(new_n150));
  xobna2aa1n03x5               g055(.a(new_n150), .b(new_n147), .c(new_n146), .out0(\s[12] ));
  nano23aa1n03x7               g056(.a(new_n142), .b(new_n148), .c(new_n149), .d(new_n143), .out0(new_n152));
  and002aa1n02x5               g057(.a(new_n152), .b(new_n139), .o(new_n153));
  aoai13aa1n03x5               g058(.a(new_n153), .b(new_n127), .c(new_n134), .d(new_n136), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n148), .o1(new_n155));
  inv020aa1n04x5               g060(.a(new_n149), .o1(new_n156));
  aoai13aa1n12x5               g061(.a(new_n143), .b(new_n137), .c(new_n97), .d(new_n138), .o1(new_n157));
  aoai13aa1n12x5               g062(.a(new_n155), .b(new_n156), .c(new_n157), .d(new_n146), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  nor042aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand42aa1n06x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n154), .c(new_n159), .out0(\s[13] ));
  aoi012aa1n03x5               g068(.a(new_n158), .b(new_n128), .c(new_n153), .o1(new_n164));
  oaoi03aa1n03x5               g069(.a(\a[13] ), .b(\b[12] ), .c(new_n164), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n03x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand02aa1d08x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nano23aa1n03x7               g073(.a(new_n160), .b(new_n167), .c(new_n168), .d(new_n161), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n158), .c(new_n128), .d(new_n153), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n167), .b(new_n160), .c(new_n168), .o1(new_n171));
  norp02aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nanp02aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x7               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n171), .out0(\s[15] ));
  nona23aa1n03x5               g080(.a(new_n168), .b(new_n161), .c(new_n160), .d(new_n167), .out0(new_n176));
  aoai13aa1n03x5               g081(.a(new_n171), .b(new_n176), .c(new_n154), .d(new_n159), .o1(new_n177));
  nor042aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand22aa1n09x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n172), .c(new_n177), .d(new_n173), .o1(new_n181));
  aoi112aa1n03x5               g086(.a(new_n172), .b(new_n180), .c(new_n177), .d(new_n173), .o1(new_n182));
  nanb02aa1n02x5               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano23aa1n06x5               g088(.a(new_n172), .b(new_n178), .c(new_n179), .d(new_n173), .out0(new_n184));
  nand22aa1n03x5               g089(.a(new_n184), .b(new_n169), .o1(new_n185));
  nano22aa1n12x5               g090(.a(new_n185), .b(new_n139), .c(new_n152), .out0(new_n186));
  aoai13aa1n09x5               g091(.a(new_n186), .b(new_n127), .c(new_n134), .d(new_n136), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n178), .o1(new_n188));
  nano32aa1n03x7               g093(.a(new_n176), .b(new_n179), .c(new_n174), .d(new_n188), .out0(new_n189));
  inv000aa1n02x5               g094(.a(new_n172), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n179), .o1(new_n191));
  aoai13aa1n02x5               g096(.a(new_n173), .b(new_n167), .c(new_n160), .d(new_n168), .o1(new_n192));
  aoai13aa1n06x5               g097(.a(new_n188), .b(new_n191), .c(new_n192), .d(new_n190), .o1(new_n193));
  aoi012aa1d18x5               g098(.a(new_n193), .b(new_n158), .c(new_n189), .o1(new_n194));
  nor022aa1n06x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  nand42aa1n03x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  norb02aa1n02x5               g101(.a(new_n196), .b(new_n195), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n187), .c(new_n194), .out0(\s[17] ));
  nand02aa1d04x5               g103(.a(new_n187), .b(new_n194), .o1(new_n199));
  tech160nm_fiaoi012aa1n05x5   g104(.a(new_n195), .b(new_n199), .c(new_n197), .o1(new_n200));
  xnrb03aa1n03x5               g105(.a(new_n200), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n06x5               g106(.a(new_n158), .b(new_n189), .o1(new_n202));
  inv000aa1n02x5               g107(.a(new_n193), .o1(new_n203));
  nanp02aa1n06x5               g108(.a(new_n202), .b(new_n203), .o1(new_n204));
  nor002aa1n02x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nand42aa1n06x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nano23aa1n06x5               g111(.a(new_n195), .b(new_n205), .c(new_n206), .d(new_n196), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n204), .c(new_n128), .d(new_n186), .o1(new_n208));
  oa0012aa1n06x5               g113(.a(new_n206), .b(new_n205), .c(new_n195), .o(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor042aa1n03x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand42aa1n03x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n03x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n208), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand22aa1n02x5               g120(.a(new_n208), .b(new_n210), .o1(new_n216));
  nor042aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanp02aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n211), .c(new_n216), .d(new_n212), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n213), .b(new_n209), .c(new_n199), .d(new_n207), .o1(new_n221));
  nona22aa1n02x5               g126(.a(new_n221), .b(new_n219), .c(new_n211), .out0(new_n222));
  nanp02aa1n02x5               g127(.a(new_n220), .b(new_n222), .o1(\s[20] ));
  nanb03aa1n12x5               g128(.a(new_n219), .b(new_n207), .c(new_n213), .out0(new_n224));
  nanb03aa1n06x5               g129(.a(new_n217), .b(new_n218), .c(new_n212), .out0(new_n225));
  oaih22aa1n04x5               g130(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[18] ), .o1(new_n227));
  nanb02aa1n02x5               g132(.a(\a[19] ), .b(new_n227), .out0(new_n228));
  nanp03aa1n03x5               g133(.a(new_n226), .b(new_n228), .c(new_n206), .o1(new_n229));
  aoi012aa1n09x5               g134(.a(new_n217), .b(new_n211), .c(new_n218), .o1(new_n230));
  oai012aa1n18x5               g135(.a(new_n230), .b(new_n229), .c(new_n225), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n224), .c(new_n187), .d(new_n194), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[20] ), .b(\a[21] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  inv030aa1n02x5               g140(.a(new_n224), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(new_n235), .b(new_n231), .c(new_n199), .d(new_n236), .o1(new_n237));
  aoi012aa1n02x5               g142(.a(new_n237), .b(new_n233), .c(new_n235), .o1(\s[21] ));
  norp02aa1n02x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  tech160nm_fixnrc02aa1n04x5   g144(.a(\b[21] ), .b(\a[22] ), .out0(new_n240));
  aoai13aa1n04x5               g145(.a(new_n240), .b(new_n239), .c(new_n233), .d(new_n235), .o1(new_n241));
  aoi112aa1n03x5               g146(.a(new_n239), .b(new_n240), .c(new_n233), .d(new_n235), .o1(new_n242));
  nanb02aa1n03x5               g147(.a(new_n242), .b(new_n241), .out0(\s[22] ));
  nor042aa1n04x5               g148(.a(new_n240), .b(new_n234), .o1(new_n244));
  nanb02aa1n02x5               g149(.a(new_n224), .b(new_n244), .out0(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oao003aa1n02x5               g152(.a(new_n246), .b(new_n247), .c(new_n239), .carry(new_n248));
  aoi012aa1n02x5               g153(.a(new_n248), .b(new_n231), .c(new_n244), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n245), .c(new_n187), .d(new_n194), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  xnrc02aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .out0(new_n254));
  aoai13aa1n02x7               g159(.a(new_n254), .b(new_n252), .c(new_n250), .d(new_n253), .o1(new_n255));
  aoi112aa1n03x5               g160(.a(new_n252), .b(new_n254), .c(new_n250), .d(new_n253), .o1(new_n256));
  nanb02aa1n03x5               g161(.a(new_n256), .b(new_n255), .out0(\s[24] ));
  inv000aa1n02x5               g162(.a(new_n244), .o1(new_n258));
  nanb02aa1d24x5               g163(.a(new_n254), .b(new_n253), .out0(new_n259));
  nor043aa1n02x5               g164(.a(new_n224), .b(new_n258), .c(new_n259), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n204), .c(new_n128), .d(new_n186), .o1(new_n261));
  nano22aa1n02x4               g166(.a(new_n217), .b(new_n212), .c(new_n218), .out0(new_n262));
  oai012aa1n02x5               g167(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .o1(new_n263));
  oab012aa1n06x5               g168(.a(new_n263), .b(new_n195), .c(new_n205), .out0(new_n264));
  inv000aa1n02x5               g169(.a(new_n230), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n244), .b(new_n265), .c(new_n264), .d(new_n262), .o1(new_n266));
  inv000aa1n02x5               g171(.a(new_n248), .o1(new_n267));
  orn002aa1n02x5               g172(.a(\a[23] ), .b(\b[22] ), .o(new_n268));
  oao003aa1n02x5               g173(.a(\a[24] ), .b(\b[23] ), .c(new_n268), .carry(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n259), .c(new_n266), .d(new_n267), .o1(new_n270));
  nanb02aa1n06x5               g175(.a(new_n270), .b(new_n261), .out0(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  norp02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .o1(new_n275));
  nanp02aa1n02x5               g180(.a(\b[25] ), .b(\a[26] ), .o1(new_n276));
  nanb02aa1n02x5               g181(.a(new_n275), .b(new_n276), .out0(new_n277));
  aoai13aa1n02x5               g182(.a(new_n277), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n274), .b(new_n270), .c(new_n199), .d(new_n260), .o1(new_n279));
  nona22aa1n02x5               g184(.a(new_n279), .b(new_n277), .c(new_n273), .out0(new_n280));
  nanp02aa1n02x5               g185(.a(new_n278), .b(new_n280), .o1(\s[26] ));
  norb02aa1n06x5               g186(.a(new_n274), .b(new_n277), .out0(new_n282));
  nano23aa1n06x5               g187(.a(new_n224), .b(new_n259), .c(new_n282), .d(new_n244), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n204), .c(new_n128), .d(new_n186), .o1(new_n284));
  oai012aa1n02x5               g189(.a(new_n276), .b(new_n275), .c(new_n273), .o1(new_n285));
  aobi12aa1n06x5               g190(.a(new_n285), .b(new_n270), .c(new_n282), .out0(new_n286));
  xorc02aa1n02x5               g191(.a(\a[27] ), .b(\b[26] ), .out0(new_n287));
  xnbna2aa1n03x5               g192(.a(new_n287), .b(new_n286), .c(new_n284), .out0(\s[27] ));
  nand42aa1n04x5               g193(.a(new_n286), .b(new_n284), .o1(new_n289));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[28] ), .b(\b[27] ), .out0(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n290), .c(new_n289), .d(new_n287), .o1(new_n293));
  nona23aa1n06x5               g198(.a(new_n236), .b(new_n282), .c(new_n259), .d(new_n258), .out0(new_n294));
  aoi012aa1n06x5               g199(.a(new_n294), .b(new_n187), .c(new_n194), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n259), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n248), .c(new_n231), .d(new_n244), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n282), .o1(new_n298));
  aoai13aa1n06x5               g203(.a(new_n285), .b(new_n298), .c(new_n297), .d(new_n269), .o1(new_n299));
  oaih12aa1n02x5               g204(.a(new_n287), .b(new_n299), .c(new_n295), .o1(new_n300));
  nona22aa1n03x5               g205(.a(new_n300), .b(new_n292), .c(new_n290), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n293), .b(new_n301), .o1(\s[28] ));
  xnrc02aa1n02x5               g207(.a(\b[28] ), .b(\a[29] ), .out0(new_n303));
  and002aa1n06x5               g208(.a(new_n291), .b(new_n287), .o(new_n304));
  oaih12aa1n02x5               g209(.a(new_n304), .b(new_n299), .c(new_n295), .o1(new_n305));
  aoi112aa1n09x5               g210(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n306));
  oab012aa1n06x5               g211(.a(new_n306), .b(\a[28] ), .c(\b[27] ), .out0(new_n307));
  aoi012aa1n03x5               g212(.a(new_n303), .b(new_n305), .c(new_n307), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n304), .o1(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n309), .b(new_n286), .c(new_n284), .o1(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n303), .c(new_n307), .out0(new_n311));
  nor002aa1n02x5               g216(.a(new_n308), .b(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g217(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g218(.a(new_n303), .b(new_n287), .c(new_n291), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n314), .b(new_n299), .c(new_n295), .o1(new_n315));
  tech160nm_fioaoi03aa1n03p5x5 g220(.a(\a[29] ), .b(\b[28] ), .c(new_n307), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n316), .o1(new_n317));
  nanp02aa1n03x5               g222(.a(new_n315), .b(new_n317), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  norp02aa1n02x5               g224(.a(new_n316), .b(new_n319), .o1(new_n320));
  aoi022aa1n02x7               g225(.a(new_n318), .b(new_n319), .c(new_n315), .d(new_n320), .o1(\s[30] ));
  nano32aa1n02x4               g226(.a(new_n303), .b(new_n319), .c(new_n287), .d(new_n291), .out0(new_n322));
  oaih12aa1n02x5               g227(.a(new_n322), .b(new_n299), .c(new_n295), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[31] ), .b(\b[30] ), .out0(new_n324));
  inv000aa1d42x5               g229(.a(\a[30] ), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[29] ), .o1(new_n326));
  oabi12aa1n02x5               g231(.a(new_n324), .b(\a[30] ), .c(\b[29] ), .out0(new_n327));
  oaoi13aa1n02x5               g232(.a(new_n327), .b(new_n316), .c(new_n325), .d(new_n326), .o1(new_n328));
  oaoi03aa1n02x5               g233(.a(new_n325), .b(new_n326), .c(new_n316), .o1(new_n329));
  nanp02aa1n03x5               g234(.a(new_n323), .b(new_n329), .o1(new_n330));
  aoi022aa1n02x7               g235(.a(new_n330), .b(new_n324), .c(new_n323), .d(new_n328), .o1(\s[31] ));
  norb02aa1n02x5               g236(.a(new_n105), .b(new_n104), .out0(new_n332));
  xnrc02aa1n02x5               g237(.a(new_n132), .b(new_n332), .out0(\s[3] ));
  obai22aa1n02x7               g238(.a(new_n102), .b(new_n103), .c(\a[3] ), .d(\b[2] ), .out0(new_n334));
  aoi012aa1n02x5               g239(.a(new_n334), .b(new_n101), .c(new_n332), .o1(new_n335));
  oaoi13aa1n02x5               g240(.a(new_n335), .b(new_n134), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  oai112aa1n02x5               g241(.a(new_n107), .b(new_n110), .c(new_n133), .d(new_n132), .o1(new_n337));
  aobi12aa1n02x5               g242(.a(new_n337), .b(new_n111), .c(new_n134), .out0(\s[5] ));
  tech160nm_fiaoi012aa1n05x5   g243(.a(new_n122), .b(new_n134), .c(new_n111), .o1(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(new_n120), .out0(\s[6] ));
  nanb02aa1n02x5               g245(.a(new_n109), .b(new_n339), .out0(new_n341));
  oai112aa1n03x5               g246(.a(new_n341), .b(new_n118), .c(new_n121), .d(new_n120), .o1(new_n342));
  oaoi13aa1n02x5               g247(.a(new_n118), .b(new_n341), .c(new_n120), .d(new_n121), .o1(new_n343));
  norb02aa1n02x5               g248(.a(new_n342), .b(new_n343), .out0(\s[7] ));
  xobna2aa1n03x5               g249(.a(new_n114), .b(new_n342), .c(new_n125), .out0(\s[8] ));
  norb02aa1n02x5               g250(.a(new_n129), .b(new_n97), .out0(new_n346));
  aoi112aa1n02x5               g251(.a(new_n346), .b(new_n127), .c(new_n134), .d(new_n136), .o1(new_n347));
  aoi012aa1n02x5               g252(.a(new_n347), .b(new_n128), .c(new_n346), .o1(\s[9] ));
endmodule


