// Benchmark "adder" written by ABC on Thu Jul 11 11:55:28 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n174,
    new_n175, new_n176, new_n177, new_n179, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n292, new_n295, new_n297, new_n298, new_n300;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  and002aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o(new_n98));
  nanp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  norp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai012aa1n02x5               g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  norp02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n02x4               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  aoi012aa1n02x5               g012(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n108));
  oai012aa1n02x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  norp02aa1n02x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n02x4               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  norp03aa1n02x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n109), .b(new_n117), .o1(new_n118));
  orn002aa1n02x5               g023(.a(\a[5] ), .b(\b[4] ), .o(new_n119));
  oao003aa1n02x5               g024(.a(\a[6] ), .b(\b[5] ), .c(new_n119), .carry(new_n120));
  160nm_fiao0012aa1n02p5x5     g025(.a(new_n110), .b(new_n112), .c(new_n111), .o(new_n121));
  oab012aa1n02x4               g026(.a(new_n121), .b(new_n120), .c(new_n114), .out0(new_n122));
  aoai13aa1n02x5               g027(.a(new_n97), .b(new_n98), .c(new_n122), .d(new_n118), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xorc02aa1n02x5               g029(.a(\a[10] ), .b(\b[9] ), .out0(new_n125));
  norp02aa1n02x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  oaoi03aa1n02x5               g033(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n129));
  aoai13aa1n02x5               g034(.a(new_n128), .b(new_n129), .c(new_n123), .d(new_n125), .o1(new_n130));
  aoi112aa1n02x5               g035(.a(new_n128), .b(new_n129), .c(new_n123), .d(new_n125), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(\s[11] ));
  norp02aa1n02x5               g037(.a(\b[11] ), .b(\a[12] ), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  nona22aa1n02x4               g040(.a(new_n130), .b(new_n135), .c(new_n126), .out0(new_n136));
  160nm_ficinv00aa1n08x5       g041(.clk(new_n126), .clkout(new_n137));
  aobi12aa1n02x5               g042(.a(new_n135), .b(new_n130), .c(new_n137), .out0(new_n138));
  norb02aa1n02x5               g043(.a(new_n136), .b(new_n138), .out0(\s[12] ));
  oabi12aa1n02x5               g044(.a(new_n121), .b(new_n120), .c(new_n114), .out0(new_n140));
  nano23aa1n02x4               g045(.a(new_n126), .b(new_n133), .c(new_n134), .d(new_n127), .out0(new_n141));
  xorc02aa1n02x5               g046(.a(\a[9] ), .b(\b[8] ), .out0(new_n142));
  and003aa1n02x5               g047(.a(new_n141), .b(new_n125), .c(new_n142), .o(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n140), .c(new_n109), .d(new_n117), .o1(new_n144));
  oaoi03aa1n02x5               g049(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .o1(new_n145));
  aoi012aa1n02x5               g050(.a(new_n145), .b(new_n141), .c(new_n129), .o1(new_n146));
  xorc02aa1n02x5               g051(.a(\a[13] ), .b(\b[12] ), .out0(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n146), .out0(\s[13] ));
  orn002aa1n02x5               g053(.a(\a[13] ), .b(\b[12] ), .o(new_n149));
  aob012aa1n02x5               g054(.a(new_n147), .b(new_n144), .c(new_n146), .out0(new_n150));
  xorc02aa1n02x5               g055(.a(\a[14] ), .b(\b[13] ), .out0(new_n151));
  xnbna2aa1n03x5               g056(.a(new_n151), .b(new_n150), .c(new_n149), .out0(\s[14] ));
  nanp02aa1n02x5               g057(.a(new_n151), .b(new_n147), .o1(new_n153));
  oao003aa1n02x5               g058(.a(\a[14] ), .b(\b[13] ), .c(new_n149), .carry(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n153), .c(new_n144), .d(new_n146), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g061(.a(\b[14] ), .b(\a[15] ), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(\b[14] ), .b(\a[15] ), .o1(new_n158));
  norp02aa1n02x5               g063(.a(\b[15] ), .b(\a[16] ), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(\b[15] ), .b(\a[16] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  aoi112aa1n02x5               g066(.a(new_n161), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n162));
  aoai13aa1n02x5               g067(.a(new_n161), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(\s[16] ));
  nano23aa1n02x4               g069(.a(new_n157), .b(new_n159), .c(new_n160), .d(new_n158), .out0(new_n165));
  nanp03aa1n02x5               g070(.a(new_n165), .b(new_n147), .c(new_n151), .o1(new_n166));
  nano32aa1n02x4               g071(.a(new_n166), .b(new_n142), .c(new_n141), .d(new_n125), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n140), .c(new_n109), .d(new_n117), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n169));
  oaib12aa1n02x5               g074(.a(new_n169), .b(new_n154), .c(new_n165), .out0(new_n170));
  oab012aa1n02x4               g075(.a(new_n170), .b(new_n146), .c(new_n166), .out0(new_n171));
  nanp02aa1n02x5               g076(.a(new_n168), .b(new_n171), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g078(.clk(\a[18] ), .clkout(new_n174));
  160nm_ficinv00aa1n08x5       g079(.clk(\a[17] ), .clkout(new_n175));
  160nm_ficinv00aa1n08x5       g080(.clk(\b[16] ), .clkout(new_n176));
  oaoi03aa1n02x5               g081(.a(new_n175), .b(new_n176), .c(new_n172), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[17] ), .c(new_n174), .out0(\s[18] ));
  xroi22aa1d04x5               g083(.a(new_n175), .b(\b[16] ), .c(new_n174), .d(\b[17] ), .out0(new_n179));
  nanp02aa1n02x5               g084(.a(new_n176), .b(new_n175), .o1(new_n180));
  oaoi03aa1n02x5               g085(.a(\a[18] ), .b(\b[17] ), .c(new_n180), .o1(new_n181));
  norp02aa1n02x5               g086(.a(\b[18] ), .b(\a[19] ), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(\b[18] ), .b(\a[19] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n181), .c(new_n172), .d(new_n179), .o1(new_n185));
  aoi112aa1n02x5               g090(.a(new_n184), .b(new_n181), .c(new_n172), .d(new_n179), .o1(new_n186));
  norb02aa1n02x5               g091(.a(new_n185), .b(new_n186), .out0(\s[19] ));
  xnrc02aa1n02x5               g092(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g093(.a(\b[19] ), .b(\a[20] ), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(\b[19] ), .b(\a[20] ), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n190), .b(new_n189), .out0(new_n191));
  nona22aa1n02x4               g096(.a(new_n185), .b(new_n191), .c(new_n182), .out0(new_n192));
  160nm_ficinv00aa1n08x5       g097(.clk(new_n191), .clkout(new_n193));
  oaoi13aa1n02x5               g098(.a(new_n193), .b(new_n185), .c(\a[19] ), .d(\b[18] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n192), .b(new_n194), .out0(\s[20] ));
  nano23aa1n02x4               g100(.a(new_n182), .b(new_n189), .c(new_n190), .d(new_n183), .out0(new_n196));
  nanp02aa1n02x5               g101(.a(new_n179), .b(new_n196), .o1(new_n197));
  oai022aa1n02x5               g102(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n198));
  oaib12aa1n02x5               g103(.a(new_n198), .b(new_n174), .c(\b[17] ), .out0(new_n199));
  nona23aa1n02x4               g104(.a(new_n190), .b(new_n183), .c(new_n182), .d(new_n189), .out0(new_n200));
  aoi012aa1n02x5               g105(.a(new_n189), .b(new_n182), .c(new_n190), .o1(new_n201));
  oai012aa1n02x5               g106(.a(new_n201), .b(new_n200), .c(new_n199), .o1(new_n202));
  160nm_ficinv00aa1n08x5       g107(.clk(new_n202), .clkout(new_n203));
  aoai13aa1n02x5               g108(.a(new_n203), .b(new_n197), .c(new_n168), .d(new_n171), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g110(.a(\b[20] ), .b(\a[21] ), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[21] ), .b(\b[20] ), .out0(new_n207));
  xorc02aa1n02x5               g112(.a(\a[22] ), .b(\b[21] ), .out0(new_n208));
  aoi112aa1n02x5               g113(.a(new_n206), .b(new_n208), .c(new_n204), .d(new_n207), .o1(new_n209));
  aoai13aa1n02x5               g114(.a(new_n208), .b(new_n206), .c(new_n204), .d(new_n207), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(\s[22] ));
  160nm_ficinv00aa1n08x5       g116(.clk(\a[21] ), .clkout(new_n212));
  160nm_ficinv00aa1n08x5       g117(.clk(\a[22] ), .clkout(new_n213));
  xroi22aa1d04x5               g118(.a(new_n212), .b(\b[20] ), .c(new_n213), .d(\b[21] ), .out0(new_n214));
  nanp03aa1n02x5               g119(.a(new_n214), .b(new_n179), .c(new_n196), .o1(new_n215));
  160nm_ficinv00aa1n08x5       g120(.clk(\b[21] ), .clkout(new_n216));
  oaoi03aa1n02x5               g121(.a(new_n213), .b(new_n216), .c(new_n206), .o1(new_n217));
  160nm_ficinv00aa1n08x5       g122(.clk(new_n217), .clkout(new_n218));
  aoi012aa1n02x5               g123(.a(new_n218), .b(new_n202), .c(new_n214), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n215), .c(new_n168), .d(new_n171), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g126(.a(\b[22] ), .b(\a[23] ), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[23] ), .b(\b[22] ), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[24] ), .b(\b[23] ), .out0(new_n224));
  aoi112aa1n02x5               g129(.a(new_n222), .b(new_n224), .c(new_n220), .d(new_n223), .o1(new_n225));
  aoai13aa1n02x5               g130(.a(new_n224), .b(new_n222), .c(new_n220), .d(new_n223), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(\s[24] ));
  and002aa1n02x5               g132(.a(new_n224), .b(new_n223), .o(new_n228));
  160nm_ficinv00aa1n08x5       g133(.clk(new_n228), .clkout(new_n229));
  nano32aa1n02x4               g134(.a(new_n229), .b(new_n214), .c(new_n179), .d(new_n196), .out0(new_n230));
  160nm_ficinv00aa1n08x5       g135(.clk(new_n201), .clkout(new_n231));
  aoai13aa1n02x5               g136(.a(new_n214), .b(new_n231), .c(new_n196), .d(new_n181), .o1(new_n232));
  aoi112aa1n02x5               g137(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n233));
  oab012aa1n02x4               g138(.a(new_n233), .b(\a[24] ), .c(\b[23] ), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n229), .c(new_n232), .d(new_n217), .o1(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(new_n172), .c(new_n230), .o1(new_n236));
  xnrc02aa1n02x5               g141(.a(\b[24] ), .b(\a[25] ), .out0(new_n237));
  160nm_ficinv00aa1n08x5       g142(.clk(new_n237), .clkout(new_n238));
  xnrc02aa1n02x5               g143(.a(new_n236), .b(new_n238), .out0(\s[25] ));
  norp02aa1n02x5               g144(.a(\b[24] ), .b(\a[25] ), .o1(new_n240));
  160nm_ficinv00aa1n08x5       g145(.clk(new_n240), .clkout(new_n241));
  aoai13aa1n02x5               g146(.a(new_n238), .b(new_n235), .c(new_n172), .d(new_n230), .o1(new_n242));
  xnrc02aa1n02x5               g147(.a(\b[25] ), .b(\a[26] ), .out0(new_n243));
  nanp03aa1n02x5               g148(.a(new_n242), .b(new_n241), .c(new_n243), .o1(new_n244));
  aoi012aa1n02x5               g149(.a(new_n243), .b(new_n242), .c(new_n241), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n244), .b(new_n245), .out0(\s[26] ));
  norp02aa1n02x5               g151(.a(new_n243), .b(new_n237), .o1(new_n247));
  nano22aa1n02x4               g152(.a(new_n215), .b(new_n228), .c(new_n247), .out0(new_n248));
  nanp02aa1n02x5               g153(.a(new_n172), .b(new_n248), .o1(new_n249));
  oao003aa1n02x5               g154(.a(\a[26] ), .b(\b[25] ), .c(new_n241), .carry(new_n250));
  aobi12aa1n02x5               g155(.a(new_n250), .b(new_n235), .c(new_n247), .out0(new_n251));
  xorc02aa1n02x5               g156(.a(\a[27] ), .b(\b[26] ), .out0(new_n252));
  xnbna2aa1n03x5               g157(.a(new_n252), .b(new_n251), .c(new_n249), .out0(\s[27] ));
  norp02aa1n02x5               g158(.a(\b[26] ), .b(\a[27] ), .o1(new_n254));
  160nm_ficinv00aa1n08x5       g159(.clk(new_n254), .clkout(new_n255));
  aobi12aa1n02x5               g160(.a(new_n252), .b(new_n251), .c(new_n249), .out0(new_n256));
  xnrc02aa1n02x5               g161(.a(\b[27] ), .b(\a[28] ), .out0(new_n257));
  nano22aa1n02x4               g162(.a(new_n256), .b(new_n255), .c(new_n257), .out0(new_n258));
  aobi12aa1n02x5               g163(.a(new_n248), .b(new_n168), .c(new_n171), .out0(new_n259));
  aoai13aa1n02x5               g164(.a(new_n228), .b(new_n218), .c(new_n202), .d(new_n214), .o1(new_n260));
  160nm_ficinv00aa1n08x5       g165(.clk(new_n247), .clkout(new_n261));
  aoai13aa1n02x5               g166(.a(new_n250), .b(new_n261), .c(new_n260), .d(new_n234), .o1(new_n262));
  oai012aa1n02x5               g167(.a(new_n252), .b(new_n262), .c(new_n259), .o1(new_n263));
  aoi012aa1n02x5               g168(.a(new_n257), .b(new_n263), .c(new_n255), .o1(new_n264));
  norp02aa1n02x5               g169(.a(new_n264), .b(new_n258), .o1(\s[28] ));
  norb02aa1n02x5               g170(.a(new_n252), .b(new_n257), .out0(new_n266));
  oai012aa1n02x5               g171(.a(new_n266), .b(new_n262), .c(new_n259), .o1(new_n267));
  oao003aa1n02x5               g172(.a(\a[28] ), .b(\b[27] ), .c(new_n255), .carry(new_n268));
  xnrc02aa1n02x5               g173(.a(\b[28] ), .b(\a[29] ), .out0(new_n269));
  aoi012aa1n02x5               g174(.a(new_n269), .b(new_n267), .c(new_n268), .o1(new_n270));
  aobi12aa1n02x5               g175(.a(new_n266), .b(new_n251), .c(new_n249), .out0(new_n271));
  nano22aa1n02x4               g176(.a(new_n271), .b(new_n268), .c(new_n269), .out0(new_n272));
  norp02aa1n02x5               g177(.a(new_n270), .b(new_n272), .o1(\s[29] ));
  xorb03aa1n02x5               g178(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g179(.a(new_n252), .b(new_n269), .c(new_n257), .out0(new_n275));
  oai012aa1n02x5               g180(.a(new_n275), .b(new_n262), .c(new_n259), .o1(new_n276));
  oao003aa1n02x5               g181(.a(\a[29] ), .b(\b[28] ), .c(new_n268), .carry(new_n277));
  xnrc02aa1n02x5               g182(.a(\b[29] ), .b(\a[30] ), .out0(new_n278));
  aoi012aa1n02x5               g183(.a(new_n278), .b(new_n276), .c(new_n277), .o1(new_n279));
  aobi12aa1n02x5               g184(.a(new_n275), .b(new_n251), .c(new_n249), .out0(new_n280));
  nano22aa1n02x4               g185(.a(new_n280), .b(new_n277), .c(new_n278), .out0(new_n281));
  norp02aa1n02x5               g186(.a(new_n279), .b(new_n281), .o1(\s[30] ));
  xnrc02aa1n02x5               g187(.a(\b[30] ), .b(\a[31] ), .out0(new_n283));
  norb02aa1n02x5               g188(.a(new_n275), .b(new_n278), .out0(new_n284));
  aobi12aa1n02x5               g189(.a(new_n284), .b(new_n251), .c(new_n249), .out0(new_n285));
  oao003aa1n02x5               g190(.a(\a[30] ), .b(\b[29] ), .c(new_n277), .carry(new_n286));
  nano22aa1n02x4               g191(.a(new_n285), .b(new_n283), .c(new_n286), .out0(new_n287));
  oai012aa1n02x5               g192(.a(new_n284), .b(new_n262), .c(new_n259), .o1(new_n288));
  aoi012aa1n02x5               g193(.a(new_n283), .b(new_n288), .c(new_n286), .o1(new_n289));
  norp02aa1n02x5               g194(.a(new_n289), .b(new_n287), .o1(\s[31] ));
  xnrb03aa1n02x5               g195(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g196(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n292));
  xorb03aa1n02x5               g197(.a(new_n292), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g198(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g199(.a(new_n116), .b(new_n109), .out0(new_n295));
  xobna2aa1n03x5               g200(.a(new_n115), .b(new_n295), .c(new_n119), .out0(\s[6] ));
  norp02aa1n02x5               g201(.a(new_n116), .b(new_n115), .o1(new_n297));
  aob012aa1n02x5               g202(.a(new_n120), .b(new_n109), .c(new_n297), .out0(new_n298));
  xorb03aa1n02x5               g203(.a(new_n298), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g204(.a(new_n112), .b(new_n298), .c(new_n113), .o1(new_n300));
  xnrb03aa1n02x5               g205(.a(new_n300), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g206(.a(new_n142), .b(new_n122), .c(new_n118), .out0(\s[9] ));
endmodule


