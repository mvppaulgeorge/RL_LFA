// Benchmark "adder" written by ABC on Wed Jul 17 13:49:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n156, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n327, new_n330, new_n332, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv030aa1d32x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1n16x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  and002aa1n06x5               g004(.a(\b[3] ), .b(\a[4] ), .o(new_n100));
  inv000aa1d42x5               g005(.a(\a[3] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[2] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(new_n103), .b(new_n104), .o1(new_n105));
  norp02aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  aoi022aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n107));
  nor042aa1n02x5               g012(.a(new_n107), .b(new_n106), .o1(new_n108));
  oa0022aa1n09x5               g013(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n109));
  oaoi13aa1n12x5               g014(.a(new_n100), .b(new_n109), .c(new_n108), .d(new_n105), .o1(new_n110));
  xorc02aa1n02x5               g015(.a(\a[6] ), .b(\b[5] ), .out0(new_n111));
  nor042aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  norb02aa1n06x4               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  xorc02aa1n12x5               g019(.a(\a[7] ), .b(\b[6] ), .out0(new_n115));
  nanp02aa1n02x5               g020(.a(new_n115), .b(new_n114), .o1(new_n116));
  xorc02aa1n02x5               g021(.a(\a[5] ), .b(\b[4] ), .out0(new_n117));
  nano22aa1n02x4               g022(.a(new_n116), .b(new_n111), .c(new_n117), .out0(new_n118));
  nanp02aa1n02x5               g023(.a(new_n110), .b(new_n118), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n112), .o1(new_n120));
  aoi112aa1n02x5               g025(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n121), .o1(new_n122));
  and002aa1n18x5               g027(.a(\b[5] ), .b(\a[6] ), .o(new_n123));
  inv000aa1d42x5               g028(.a(new_n123), .o1(new_n124));
  nanb02aa1n02x5               g029(.a(new_n112), .b(new_n113), .out0(new_n125));
  xnrc02aa1n02x5               g030(.a(\b[6] ), .b(\a[7] ), .out0(new_n126));
  oai022aa1n02x5               g031(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n127));
  nano23aa1n02x4               g032(.a(new_n126), .b(new_n125), .c(new_n124), .d(new_n127), .out0(new_n128));
  nano22aa1n02x4               g033(.a(new_n128), .b(new_n120), .c(new_n122), .out0(new_n129));
  nanp02aa1n02x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(new_n99), .b(new_n130), .o1(new_n131));
  aoai13aa1n06x5               g036(.a(new_n99), .b(new_n131), .c(new_n119), .d(new_n129), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1d32x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nand42aa1d28x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanb02aa1d24x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  inv000aa1d42x5               g041(.a(new_n100), .o1(new_n137));
  xorc02aa1n02x5               g042(.a(\a[3] ), .b(\b[2] ), .out0(new_n138));
  and002aa1n02x5               g043(.a(\b[0] ), .b(\a[1] ), .o(new_n139));
  oaoi03aa1n02x5               g044(.a(\a[2] ), .b(\b[1] ), .c(new_n139), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n109), .o1(new_n141));
  aoai13aa1n02x5               g046(.a(new_n137), .b(new_n141), .c(new_n140), .d(new_n138), .o1(new_n142));
  nona23aa1n02x4               g047(.a(new_n111), .b(new_n117), .c(new_n126), .d(new_n125), .out0(new_n143));
  oai012aa1n02x5               g048(.a(new_n129), .b(new_n142), .c(new_n143), .o1(new_n144));
  oaoi03aa1n02x5               g049(.a(new_n97), .b(new_n98), .c(new_n144), .o1(new_n145));
  nor002aa1n03x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  nand22aa1n03x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n12x5               g054(.a(new_n135), .b(new_n134), .c(new_n97), .d(new_n98), .o1(new_n150));
  oaoi13aa1n02x5               g055(.a(new_n149), .b(new_n150), .c(new_n145), .d(new_n136), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n136), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n150), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n148), .b(new_n153), .c(new_n132), .d(new_n152), .o1(new_n154));
  norp02aa1n02x5               g059(.a(new_n151), .b(new_n154), .o1(\s[11] ));
  aoai13aa1n02x5               g060(.a(new_n148), .b(new_n153), .c(new_n132), .d(new_n152), .o1(new_n156));
  nor042aa1n12x5               g061(.a(\b[11] ), .b(\a[12] ), .o1(new_n157));
  nand02aa1n04x5               g062(.a(\b[11] ), .b(\a[12] ), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n157), .b(new_n158), .out0(new_n159));
  oai112aa1n02x5               g064(.a(new_n156), .b(new_n159), .c(\b[10] ), .d(\a[11] ), .o1(new_n160));
  oaoi13aa1n02x5               g065(.a(new_n159), .b(new_n156), .c(\a[11] ), .d(\b[10] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(\s[12] ));
  nano23aa1n06x5               g067(.a(new_n146), .b(new_n157), .c(new_n158), .d(new_n147), .out0(new_n163));
  nona22aa1d18x5               g068(.a(new_n163), .b(new_n136), .c(new_n131), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n157), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n158), .b(new_n147), .c(new_n146), .d(new_n157), .out0(new_n166));
  nanp02aa1n02x5               g071(.a(new_n146), .b(new_n158), .o1(new_n167));
  oai112aa1n06x5               g072(.a(new_n167), .b(new_n165), .c(new_n166), .d(new_n150), .o1(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n164), .c(new_n119), .d(new_n129), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[12] ), .b(\a[13] ), .o1(new_n173));
  aoi012aa1n02x5               g078(.a(new_n172), .b(new_n170), .c(new_n173), .o1(new_n174));
  xnrb03aa1n02x5               g079(.a(new_n174), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g080(.a(\a[6] ), .o1(new_n176));
  inv000aa1d42x5               g081(.a(\b[5] ), .o1(new_n177));
  norp02aa1n02x5               g082(.a(\b[4] ), .b(\a[5] ), .o1(new_n178));
  aoi012aa1n02x5               g083(.a(new_n178), .b(new_n176), .c(new_n177), .o1(new_n179));
  nona23aa1n02x4               g084(.a(new_n115), .b(new_n114), .c(new_n179), .d(new_n123), .out0(new_n180));
  nona22aa1n02x4               g085(.a(new_n180), .b(new_n121), .c(new_n112), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n164), .o1(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n181), .c(new_n110), .d(new_n118), .o1(new_n183));
  norp02aa1n02x5               g088(.a(\b[13] ), .b(\a[14] ), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(\b[13] ), .b(\a[14] ), .o1(new_n185));
  nona23aa1n02x4               g090(.a(new_n185), .b(new_n173), .c(new_n172), .d(new_n184), .out0(new_n186));
  oai012aa1n02x5               g091(.a(new_n185), .b(new_n184), .c(new_n172), .o1(new_n187));
  aoai13aa1n02x5               g092(.a(new_n187), .b(new_n186), .c(new_n183), .d(new_n169), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g094(.a(\b[14] ), .b(\a[15] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(\b[14] ), .b(\a[15] ), .o1(new_n191));
  nanb02aa1n09x5               g096(.a(new_n190), .b(new_n191), .out0(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  norp02aa1n02x5               g098(.a(\b[15] ), .b(\a[16] ), .o1(new_n194));
  nanp02aa1n02x5               g099(.a(\b[15] ), .b(\a[16] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aoi112aa1n02x5               g101(.a(new_n196), .b(new_n190), .c(new_n188), .d(new_n193), .o1(new_n197));
  aoai13aa1n02x5               g102(.a(new_n196), .b(new_n190), .c(new_n188), .d(new_n191), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(\s[16] ));
  nano23aa1n02x4               g104(.a(new_n172), .b(new_n184), .c(new_n185), .d(new_n173), .out0(new_n200));
  nano32aa1n03x7               g105(.a(new_n164), .b(new_n196), .c(new_n193), .d(new_n200), .out0(new_n201));
  aoai13aa1n09x5               g106(.a(new_n201), .b(new_n181), .c(new_n110), .d(new_n118), .o1(new_n202));
  nona23aa1n02x4               g107(.a(new_n195), .b(new_n191), .c(new_n190), .d(new_n194), .out0(new_n203));
  norp02aa1n02x5               g108(.a(new_n203), .b(new_n186), .o1(new_n204));
  aoi112aa1n02x5               g109(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n205));
  oai022aa1n02x5               g110(.a(new_n203), .b(new_n187), .c(\b[15] ), .d(\a[16] ), .o1(new_n206));
  aoi112aa1n09x5               g111(.a(new_n206), .b(new_n205), .c(new_n168), .d(new_n204), .o1(new_n207));
  nand02aa1d10x5               g112(.a(new_n207), .b(new_n202), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g114(.a(\a[18] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(\a[17] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(\b[16] ), .o1(new_n212));
  oaoi03aa1n03x5               g117(.a(new_n211), .b(new_n212), .c(new_n208), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[17] ), .c(new_n210), .out0(\s[18] ));
  xroi22aa1d04x5               g119(.a(new_n211), .b(\b[16] ), .c(new_n210), .d(\b[17] ), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n212), .b(new_n211), .o1(new_n216));
  oaoi03aa1n02x5               g121(.a(\a[18] ), .b(\b[17] ), .c(new_n216), .o1(new_n217));
  nor002aa1n02x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nand42aa1n03x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n217), .c(new_n208), .d(new_n215), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(new_n220), .b(new_n217), .c(new_n208), .d(new_n215), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n221), .b(new_n222), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n03x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand42aa1n03x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  nona22aa1n03x5               g132(.a(new_n221), .b(new_n227), .c(new_n218), .out0(new_n228));
  orn002aa1n02x5               g133(.a(\a[19] ), .b(\b[18] ), .o(new_n229));
  aobi12aa1n02x7               g134(.a(new_n227), .b(new_n221), .c(new_n229), .out0(new_n230));
  norb02aa1n03x4               g135(.a(new_n228), .b(new_n230), .out0(\s[20] ));
  nano23aa1n02x4               g136(.a(new_n218), .b(new_n225), .c(new_n226), .d(new_n219), .out0(new_n232));
  nanp02aa1n02x5               g137(.a(new_n215), .b(new_n232), .o1(new_n233));
  oai022aa1n02x5               g138(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n234));
  oaib12aa1n02x5               g139(.a(new_n234), .b(new_n210), .c(\b[17] ), .out0(new_n235));
  nona23aa1n02x4               g140(.a(new_n226), .b(new_n219), .c(new_n218), .d(new_n225), .out0(new_n236));
  oaoi03aa1n02x5               g141(.a(\a[20] ), .b(\b[19] ), .c(new_n229), .o1(new_n237));
  oabi12aa1n12x5               g142(.a(new_n237), .b(new_n236), .c(new_n235), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n233), .c(new_n207), .d(new_n202), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  xorc02aa1n02x5               g147(.a(\a[21] ), .b(\b[20] ), .out0(new_n243));
  xorc02aa1n02x5               g148(.a(\a[22] ), .b(\b[21] ), .out0(new_n244));
  aoi112aa1n03x5               g149(.a(new_n242), .b(new_n244), .c(new_n240), .d(new_n243), .o1(new_n245));
  aoai13aa1n03x5               g150(.a(new_n244), .b(new_n242), .c(new_n240), .d(new_n243), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n246), .b(new_n245), .out0(\s[22] ));
  inv000aa1d42x5               g152(.a(\a[21] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(\a[22] ), .o1(new_n249));
  xroi22aa1d04x5               g154(.a(new_n248), .b(\b[20] ), .c(new_n249), .d(\b[21] ), .out0(new_n250));
  nanp03aa1n02x5               g155(.a(new_n250), .b(new_n215), .c(new_n232), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\b[21] ), .o1(new_n252));
  oaoi03aa1n12x5               g157(.a(new_n249), .b(new_n252), .c(new_n242), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  aoi012aa1n02x5               g159(.a(new_n254), .b(new_n238), .c(new_n250), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n251), .c(new_n207), .d(new_n202), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  xorc02aa1n02x5               g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  xorc02aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .out0(new_n260));
  aoi112aa1n02x7               g165(.a(new_n258), .b(new_n260), .c(new_n256), .d(new_n259), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n260), .b(new_n258), .c(new_n256), .d(new_n259), .o1(new_n262));
  norb02aa1n03x4               g167(.a(new_n262), .b(new_n261), .out0(\s[24] ));
  and002aa1n06x5               g168(.a(new_n260), .b(new_n259), .o(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  nano32aa1n02x4               g170(.a(new_n265), .b(new_n250), .c(new_n215), .d(new_n232), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n250), .b(new_n237), .c(new_n232), .d(new_n217), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n268));
  oab012aa1n02x4               g173(.a(new_n268), .b(\a[24] ), .c(\b[23] ), .out0(new_n269));
  aoai13aa1n04x5               g174(.a(new_n269), .b(new_n265), .c(new_n267), .d(new_n253), .o1(new_n270));
  tech160nm_fixorc02aa1n05x5   g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n270), .c(new_n208), .d(new_n266), .o1(new_n272));
  aoi112aa1n02x5               g177(.a(new_n271), .b(new_n270), .c(new_n208), .d(new_n266), .o1(new_n273));
  norb02aa1n02x5               g178(.a(new_n272), .b(new_n273), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .out0(new_n276));
  nona22aa1n03x5               g181(.a(new_n272), .b(new_n276), .c(new_n275), .out0(new_n277));
  inv000aa1n02x5               g182(.a(new_n275), .o1(new_n278));
  aobi12aa1n02x7               g183(.a(new_n276), .b(new_n272), .c(new_n278), .out0(new_n279));
  norb02aa1n03x4               g184(.a(new_n277), .b(new_n279), .out0(\s[26] ));
  and002aa1n06x5               g185(.a(new_n276), .b(new_n271), .o(new_n281));
  nano22aa1n03x7               g186(.a(new_n251), .b(new_n264), .c(new_n281), .out0(new_n282));
  nand22aa1n12x5               g187(.a(new_n208), .b(new_n282), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .c(new_n278), .carry(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n270), .c(new_n281), .out0(new_n285));
  xorc02aa1n02x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n285), .out0(\s[27] ));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv040aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  aobi12aa1n06x5               g194(.a(new_n286), .b(new_n283), .c(new_n285), .out0(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  nano22aa1n03x7               g196(.a(new_n290), .b(new_n289), .c(new_n291), .out0(new_n292));
  inv000aa1n02x5               g197(.a(new_n282), .o1(new_n293));
  tech160nm_fiaoi012aa1n05x5   g198(.a(new_n293), .b(new_n207), .c(new_n202), .o1(new_n294));
  aoai13aa1n02x5               g199(.a(new_n264), .b(new_n254), .c(new_n238), .d(new_n250), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n281), .o1(new_n296));
  aoai13aa1n06x5               g201(.a(new_n284), .b(new_n296), .c(new_n295), .d(new_n269), .o1(new_n297));
  oaih12aa1n02x5               g202(.a(new_n286), .b(new_n297), .c(new_n294), .o1(new_n298));
  aoi012aa1n03x5               g203(.a(new_n291), .b(new_n298), .c(new_n289), .o1(new_n299));
  nor002aa1n02x5               g204(.a(new_n299), .b(new_n292), .o1(\s[28] ));
  norb02aa1n02x5               g205(.a(new_n286), .b(new_n291), .out0(new_n301));
  aobi12aa1n06x5               g206(.a(new_n301), .b(new_n283), .c(new_n285), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  nano22aa1n03x7               g209(.a(new_n302), .b(new_n303), .c(new_n304), .out0(new_n305));
  oaih12aa1n02x5               g210(.a(new_n301), .b(new_n297), .c(new_n294), .o1(new_n306));
  aoi012aa1n03x5               g211(.a(new_n304), .b(new_n306), .c(new_n303), .o1(new_n307));
  nor002aa1n02x5               g212(.a(new_n307), .b(new_n305), .o1(\s[29] ));
  xnrb03aa1n02x5               g213(.a(new_n139), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g214(.a(new_n286), .b(new_n304), .c(new_n291), .out0(new_n310));
  aobi12aa1n06x5               g215(.a(new_n310), .b(new_n283), .c(new_n285), .out0(new_n311));
  oao003aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[29] ), .b(\a[30] ), .out0(new_n313));
  nano22aa1n03x7               g218(.a(new_n311), .b(new_n312), .c(new_n313), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n310), .b(new_n297), .c(new_n294), .o1(new_n315));
  aoi012aa1n03x5               g220(.a(new_n313), .b(new_n315), .c(new_n312), .o1(new_n316));
  nor002aa1n02x5               g221(.a(new_n316), .b(new_n314), .o1(\s[30] ));
  norb02aa1n02x5               g222(.a(new_n310), .b(new_n313), .out0(new_n318));
  aobi12aa1n06x5               g223(.a(new_n318), .b(new_n283), .c(new_n285), .out0(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n320));
  xnrc02aa1n02x5               g225(.a(\b[30] ), .b(\a[31] ), .out0(new_n321));
  nano22aa1n03x7               g226(.a(new_n319), .b(new_n320), .c(new_n321), .out0(new_n322));
  oaih12aa1n02x5               g227(.a(new_n318), .b(new_n297), .c(new_n294), .o1(new_n323));
  aoi012aa1n03x5               g228(.a(new_n321), .b(new_n323), .c(new_n320), .o1(new_n324));
  nor002aa1n02x5               g229(.a(new_n324), .b(new_n322), .o1(\s[31] ));
  xnbna2aa1n03x5               g230(.a(new_n108), .b(new_n103), .c(new_n104), .out0(\s[3] ));
  oaoi03aa1n02x5               g231(.a(\a[3] ), .b(\b[2] ), .c(new_n108), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g233(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g234(.a(\a[5] ), .b(\b[4] ), .c(new_n142), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g236(.a(new_n176), .b(new_n177), .c(new_n330), .o1(new_n332));
  xnrc02aa1n02x5               g237(.a(new_n332), .b(new_n115), .out0(\s[7] ));
  oaoi03aa1n02x5               g238(.a(\a[7] ), .b(\b[6] ), .c(new_n332), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g240(.a(new_n144), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


