// Benchmark "adder" written by ABC on Wed Jul 17 19:35:38 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n296, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n316, new_n318,
    new_n319, new_n321, new_n322, new_n324, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  aoi022aa1d24x5               g003(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n99));
  oab012aa1n09x5               g004(.a(new_n99), .b(\a[2] ), .c(\b[1] ), .out0(new_n100));
  xnrc02aa1n02x5               g005(.a(\b[2] ), .b(\a[3] ), .out0(new_n101));
  inv000aa1d42x5               g006(.a(\a[3] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[2] ), .o1(new_n103));
  and002aa1n24x5               g008(.a(\b[3] ), .b(\a[4] ), .o(new_n104));
  nor042aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  aoi112aa1n06x5               g010(.a(new_n104), .b(new_n105), .c(new_n102), .d(new_n103), .o1(new_n106));
  oai012aa1n06x5               g011(.a(new_n106), .b(new_n100), .c(new_n101), .o1(new_n107));
  orn002aa1n24x5               g012(.a(\a[5] ), .b(\b[4] ), .o(new_n108));
  norp02aa1n04x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nand22aa1n09x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nanb03aa1d18x5               g015(.a(new_n109), .b(new_n108), .c(new_n110), .out0(new_n111));
  oai022aa1n02x5               g016(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n112));
  aoi022aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  aoi022aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(new_n114), .b(new_n113), .o1(new_n115));
  nor043aa1n02x5               g020(.a(new_n111), .b(new_n115), .c(new_n112), .o1(new_n116));
  nanp02aa1n09x5               g021(.a(new_n116), .b(new_n107), .o1(new_n117));
  nor042aa1d18x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(new_n118), .o1(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  and002aa1n12x5               g025(.a(\b[6] ), .b(\a[7] ), .o(new_n121));
  aoi112aa1n06x5               g026(.a(new_n121), .b(new_n118), .c(\a[6] ), .d(\b[5] ), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .out0(new_n123));
  aoi013aa1n09x5               g028(.a(new_n120), .b(new_n111), .c(new_n122), .d(new_n123), .o1(new_n124));
  xnrc02aa1n12x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n98), .b(new_n125), .c(new_n117), .d(new_n124), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xorc02aa1n03x5               g032(.a(\a[10] ), .b(\b[9] ), .out0(new_n128));
  nor042aa1n06x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  oai012aa1d24x5               g035(.a(new_n130), .b(new_n129), .c(new_n97), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nor042aa1d18x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  aoai13aa1n03x5               g040(.a(new_n135), .b(new_n132), .c(new_n126), .d(new_n128), .o1(new_n136));
  aoi112aa1n02x5               g041(.a(new_n135), .b(new_n132), .c(new_n126), .d(new_n128), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n136), .b(new_n137), .out0(\s[11] ));
  inv040aa1n06x5               g043(.a(new_n133), .o1(new_n139));
  nor022aa1n16x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  tech160nm_fiaoi012aa1n03p5x5 g048(.a(new_n143), .b(new_n136), .c(new_n139), .o1(new_n144));
  nona22aa1n02x4               g049(.a(new_n136), .b(new_n142), .c(new_n133), .out0(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(\s[12] ));
  nona23aa1d18x5               g051(.a(new_n141), .b(new_n134), .c(new_n133), .d(new_n140), .out0(new_n147));
  nona22aa1n02x4               g052(.a(new_n128), .b(new_n147), .c(new_n125), .out0(new_n148));
  oaoi03aa1n02x5               g053(.a(\a[12] ), .b(\b[11] ), .c(new_n139), .o1(new_n149));
  oab012aa1n02x4               g054(.a(new_n149), .b(new_n147), .c(new_n131), .out0(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n148), .c(new_n117), .d(new_n124), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand02aa1n04x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n16x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand02aa1n08x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nona23aa1d18x5               g063(.a(new_n158), .b(new_n154), .c(new_n153), .d(new_n157), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  oa0012aa1n02x5               g065(.a(new_n158), .b(new_n157), .c(new_n153), .o(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[14] ), .b(\a[15] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n161), .c(new_n151), .d(new_n160), .o1(new_n164));
  aoi112aa1n02x5               g069(.a(new_n163), .b(new_n161), .c(new_n151), .d(new_n160), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(\s[15] ));
  inv000aa1d42x5               g071(.a(\a[15] ), .o1(new_n167));
  inv000aa1d42x5               g072(.a(\b[14] ), .o1(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n167), .o1(new_n169));
  xnrc02aa1n12x5               g074(.a(\b[15] ), .b(\a[16] ), .out0(new_n170));
  aoi012aa1n02x5               g075(.a(new_n170), .b(new_n164), .c(new_n169), .o1(new_n171));
  nanp03aa1n02x5               g076(.a(new_n164), .b(new_n169), .c(new_n170), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(\s[16] ));
  norb03aa1n03x5               g078(.a(new_n128), .b(new_n147), .c(new_n125), .out0(new_n174));
  nor043aa1d12x5               g079(.a(new_n159), .b(new_n162), .c(new_n170), .o1(new_n175));
  nand22aa1n09x5               g080(.a(new_n174), .b(new_n175), .o1(new_n176));
  oabi12aa1n03x5               g081(.a(new_n149), .b(new_n147), .c(new_n131), .out0(new_n177));
  inv000aa1d42x5               g082(.a(\a[16] ), .o1(new_n178));
  inv000aa1d42x5               g083(.a(\b[15] ), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(new_n179), .b(new_n178), .o1(new_n180));
  and002aa1n02x5               g085(.a(\b[15] ), .b(\a[16] ), .o(new_n181));
  oai122aa1n02x7               g086(.a(new_n158), .b(new_n157), .c(new_n153), .d(new_n168), .e(new_n167), .o1(new_n182));
  aoai13aa1n06x5               g087(.a(new_n180), .b(new_n181), .c(new_n182), .d(new_n169), .o1(new_n183));
  aoi012aa1n12x5               g088(.a(new_n183), .b(new_n177), .c(new_n175), .o1(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n176), .c(new_n117), .d(new_n124), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g091(.a(\a[18] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[16] ), .o1(new_n189));
  tech160nm_fioaoi03aa1n03p5x5 g094(.a(new_n188), .b(new_n189), .c(new_n185), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(new_n187), .out0(\s[18] ));
  xroi22aa1d06x4               g096(.a(new_n188), .b(\b[16] ), .c(new_n187), .d(\b[17] ), .out0(new_n192));
  oaih22aa1n04x5               g097(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n193));
  oaib12aa1n18x5               g098(.a(new_n193), .b(new_n187), .c(\b[17] ), .out0(new_n194));
  inv000aa1d42x5               g099(.a(new_n194), .o1(new_n195));
  tech160nm_fiaoi012aa1n05x5   g100(.a(new_n195), .b(new_n185), .c(new_n192), .o1(new_n196));
  nor022aa1n16x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  nand02aa1n04x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n196), .b(new_n199), .c(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norb02aa1n02x5               g106(.a(new_n199), .b(new_n197), .out0(new_n202));
  aoai13aa1n03x5               g107(.a(new_n202), .b(new_n195), .c(new_n185), .d(new_n192), .o1(new_n203));
  norp02aa1n04x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nanp02aa1n04x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  tech160nm_fiaoi012aa1n02p5x5 g111(.a(new_n206), .b(new_n203), .c(new_n198), .o1(new_n207));
  nanp03aa1n03x5               g112(.a(new_n203), .b(new_n198), .c(new_n206), .o1(new_n208));
  norb02aa1n02x7               g113(.a(new_n208), .b(new_n207), .out0(\s[20] ));
  nona23aa1n12x5               g114(.a(new_n205), .b(new_n199), .c(new_n197), .d(new_n204), .out0(new_n210));
  inv040aa1n08x5               g115(.a(new_n210), .o1(new_n211));
  nand02aa1d06x5               g116(.a(new_n192), .b(new_n211), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  aoi012aa1n02x5               g118(.a(new_n204), .b(new_n197), .c(new_n205), .o1(new_n214));
  oai012aa1n12x5               g119(.a(new_n214), .b(new_n210), .c(new_n194), .o1(new_n215));
  tech160nm_fiaoi012aa1n05x5   g120(.a(new_n215), .b(new_n185), .c(new_n213), .o1(new_n216));
  nor002aa1n20x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  nanp02aa1n02x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n216), .b(new_n219), .c(new_n218), .out0(\s[21] ));
  norb02aa1n02x5               g125(.a(new_n219), .b(new_n217), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n215), .c(new_n185), .d(new_n213), .o1(new_n222));
  norp02aa1n04x5               g127(.a(\b[21] ), .b(\a[22] ), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(\b[21] ), .b(\a[22] ), .o1(new_n224));
  nanb02aa1n02x5               g129(.a(new_n223), .b(new_n224), .out0(new_n225));
  tech160nm_fiaoi012aa1n02p5x5 g130(.a(new_n225), .b(new_n222), .c(new_n218), .o1(new_n226));
  nanp03aa1n03x5               g131(.a(new_n222), .b(new_n218), .c(new_n225), .o1(new_n227));
  norb02aa1n02x7               g132(.a(new_n227), .b(new_n226), .out0(\s[22] ));
  nona23aa1n06x5               g133(.a(new_n224), .b(new_n219), .c(new_n217), .d(new_n223), .out0(new_n229));
  nano22aa1n02x4               g134(.a(new_n229), .b(new_n192), .c(new_n211), .out0(new_n230));
  inv000aa1n02x5               g135(.a(new_n229), .o1(new_n231));
  aoi012aa1n02x5               g136(.a(new_n223), .b(new_n217), .c(new_n224), .o1(new_n232));
  aobi12aa1n02x5               g137(.a(new_n232), .b(new_n215), .c(new_n231), .out0(new_n233));
  inv040aa1n03x5               g138(.a(new_n233), .o1(new_n234));
  tech160nm_fiaoi012aa1n05x5   g139(.a(new_n234), .b(new_n185), .c(new_n230), .o1(new_n235));
  nor002aa1n06x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nanp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  xnbna2aa1n03x5               g143(.a(new_n235), .b(new_n238), .c(new_n237), .out0(\s[23] ));
  norb02aa1n02x5               g144(.a(new_n238), .b(new_n236), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n185), .d(new_n230), .o1(new_n241));
  nor002aa1n02x5               g146(.a(\b[23] ), .b(\a[24] ), .o1(new_n242));
  nanp02aa1n02x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  tech160nm_fiaoi012aa1n02p5x5 g149(.a(new_n244), .b(new_n241), .c(new_n237), .o1(new_n245));
  nanp03aa1n03x5               g150(.a(new_n241), .b(new_n237), .c(new_n244), .o1(new_n246));
  norb02aa1n02x7               g151(.a(new_n246), .b(new_n245), .out0(\s[24] ));
  nand42aa1n02x5               g152(.a(new_n117), .b(new_n124), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n176), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(new_n177), .b(new_n175), .o1(new_n250));
  nanb02aa1n02x5               g155(.a(new_n183), .b(new_n250), .out0(new_n251));
  nona23aa1n03x5               g156(.a(new_n243), .b(new_n238), .c(new_n236), .d(new_n242), .out0(new_n252));
  norp02aa1n09x5               g157(.a(new_n252), .b(new_n229), .o1(new_n253));
  norb02aa1n06x4               g158(.a(new_n253), .b(new_n212), .out0(new_n254));
  aoai13aa1n02x5               g159(.a(new_n254), .b(new_n251), .c(new_n249), .d(new_n248), .o1(new_n255));
  aoai13aa1n02x5               g160(.a(new_n238), .b(new_n223), .c(new_n217), .d(new_n224), .o1(new_n256));
  aoi022aa1n06x5               g161(.a(new_n256), .b(new_n237), .c(\a[24] ), .d(\b[23] ), .o1(new_n257));
  aoi112aa1n03x5               g162(.a(new_n242), .b(new_n257), .c(new_n215), .d(new_n253), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[24] ), .b(\a[25] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n255), .c(new_n258), .out0(\s[25] ));
  nor042aa1n03x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  nanp02aa1n03x5               g168(.a(new_n215), .b(new_n253), .o1(new_n264));
  nona22aa1n03x5               g169(.a(new_n264), .b(new_n257), .c(new_n242), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n260), .b(new_n265), .c(new_n185), .d(new_n254), .o1(new_n266));
  xnrc02aa1n02x5               g171(.a(\b[25] ), .b(\a[26] ), .out0(new_n267));
  tech160nm_fiaoi012aa1n02p5x5 g172(.a(new_n267), .b(new_n266), .c(new_n263), .o1(new_n268));
  nanp03aa1n03x5               g173(.a(new_n266), .b(new_n263), .c(new_n267), .o1(new_n269));
  norb02aa1n02x7               g174(.a(new_n269), .b(new_n268), .out0(\s[26] ));
  nor042aa1n04x5               g175(.a(new_n267), .b(new_n259), .o1(new_n271));
  nano22aa1d15x5               g176(.a(new_n212), .b(new_n253), .c(new_n271), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n251), .c(new_n249), .d(new_n248), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n274));
  aobi12aa1n09x5               g179(.a(new_n274), .b(new_n265), .c(new_n271), .out0(new_n275));
  xorc02aa1n12x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n273), .c(new_n275), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  inv040aa1n03x5               g183(.a(new_n278), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n271), .o1(new_n280));
  tech160nm_fioai012aa1n05x5   g185(.a(new_n274), .b(new_n258), .c(new_n280), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n276), .b(new_n281), .c(new_n185), .d(new_n272), .o1(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  aoi012aa1n03x5               g188(.a(new_n283), .b(new_n282), .c(new_n279), .o1(new_n284));
  aobi12aa1n06x5               g189(.a(new_n276), .b(new_n273), .c(new_n275), .out0(new_n285));
  nano22aa1n03x7               g190(.a(new_n285), .b(new_n279), .c(new_n283), .out0(new_n286));
  norp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n276), .b(new_n283), .out0(new_n288));
  aoai13aa1n02x7               g193(.a(new_n288), .b(new_n281), .c(new_n185), .d(new_n272), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n279), .carry(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  aobi12aa1n03x5               g197(.a(new_n288), .b(new_n273), .c(new_n275), .out0(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n291), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[29] ));
  nanp02aa1n02x5               g200(.a(\b[0] ), .b(\a[1] ), .o1(new_n296));
  xorb03aa1n02x5               g201(.a(new_n296), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g202(.a(new_n276), .b(new_n291), .c(new_n283), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n281), .c(new_n185), .d(new_n272), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[29] ), .b(\a[30] ), .out0(new_n301));
  tech160nm_fiaoi012aa1n02p5x5 g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  aobi12aa1n03x5               g207(.a(new_n298), .b(new_n273), .c(new_n275), .out0(new_n303));
  nano22aa1n03x5               g208(.a(new_n303), .b(new_n300), .c(new_n301), .out0(new_n304));
  nor002aa1n02x5               g209(.a(new_n302), .b(new_n304), .o1(\s[30] ));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  norb02aa1n03x4               g211(.a(new_n298), .b(new_n301), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n281), .c(new_n185), .d(new_n272), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  aobi12aa1n06x5               g215(.a(new_n307), .b(new_n273), .c(new_n275), .out0(new_n311));
  nano22aa1n03x7               g216(.a(new_n311), .b(new_n306), .c(new_n309), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n310), .b(new_n312), .o1(\s[31] ));
  xorb03aa1n02x5               g218(.a(new_n100), .b(\b[2] ), .c(new_n102), .out0(\s[3] ));
  xnrc02aa1n02x5               g219(.a(\b[3] ), .b(\a[4] ), .out0(new_n315));
  oaoi03aa1n02x5               g220(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n316));
  aob012aa1n02x5               g221(.a(new_n107), .b(new_n316), .c(new_n315), .out0(\s[4] ));
  inv000aa1d42x5               g222(.a(new_n104), .o1(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[4] ), .b(\a[5] ), .out0(new_n319));
  xnbna2aa1n03x5               g224(.a(new_n319), .b(new_n107), .c(new_n318), .out0(\s[5] ));
  norb02aa1n02x5               g225(.a(new_n110), .b(new_n109), .out0(new_n321));
  nona22aa1n02x4               g226(.a(new_n107), .b(new_n319), .c(new_n104), .out0(new_n322));
  xnbna2aa1n03x5               g227(.a(new_n321), .b(new_n322), .c(new_n108), .out0(\s[6] ));
  norp02aa1n02x5               g228(.a(new_n121), .b(new_n118), .o1(new_n324));
  nanb02aa1n02x5               g229(.a(new_n111), .b(new_n322), .out0(new_n325));
  xobna2aa1n03x5               g230(.a(new_n324), .b(new_n325), .c(new_n110), .out0(\s[7] ));
  nanp02aa1n02x5               g231(.a(new_n325), .b(new_n122), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n123), .b(new_n327), .c(new_n119), .out0(\s[8] ));
  xobna2aa1n03x5               g233(.a(new_n125), .b(new_n117), .c(new_n124), .out0(\s[9] ));
endmodule


