// Benchmark "adder" written by ABC on Thu Jul 18 03:10:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n339, new_n340, new_n343, new_n344, new_n346, new_n347, new_n349,
    new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  nor002aa1d32x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[2] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[1] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  oaoi03aa1n02x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n02x4               g012(.a(new_n104), .b(new_n107), .c(new_n106), .d(new_n105), .out0(new_n108));
  norp02aa1n02x5               g013(.a(new_n106), .b(new_n105), .o1(new_n109));
  obai22aa1n06x5               g014(.a(new_n104), .b(new_n109), .c(new_n108), .d(new_n103), .out0(new_n110));
  nor002aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nor002aa1n12x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n03x5               g019(.a(new_n113), .b(new_n112), .c(new_n114), .d(new_n111), .out0(new_n115));
  nor002aa1n03x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanp02aa1n09x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nanb02aa1n12x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  xnrc02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .out0(new_n119));
  nor043aa1n03x5               g024(.a(new_n115), .b(new_n118), .c(new_n119), .o1(new_n120));
  aoi112aa1n02x5               g025(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n121));
  nano23aa1n02x4               g026(.a(new_n114), .b(new_n111), .c(new_n112), .d(new_n113), .out0(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  nanp03aa1n02x5               g028(.a(new_n122), .b(new_n117), .c(new_n123), .o1(new_n124));
  nona22aa1n06x5               g029(.a(new_n124), .b(new_n121), .c(new_n111), .out0(new_n125));
  tech160nm_fixorc02aa1n04x5   g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n125), .c(new_n110), .d(new_n120), .o1(new_n127));
  xobna2aa1n03x5               g032(.a(new_n97), .b(new_n127), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g033(.a(\a[10] ), .o1(new_n129));
  inv040aa1d32x5               g034(.a(\b[9] ), .o1(new_n130));
  aoi012aa1n02x5               g035(.a(new_n98), .b(new_n129), .c(new_n130), .o1(new_n131));
  aoi022aa1n06x5               g036(.a(new_n127), .b(new_n131), .c(\b[9] ), .d(\a[10] ), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv040aa1d32x5               g038(.a(\a[11] ), .o1(new_n134));
  inv000aa1d42x5               g039(.a(\b[10] ), .o1(new_n135));
  nand42aa1n03x5               g040(.a(new_n135), .b(new_n134), .o1(new_n136));
  xnrc02aa1n02x5               g041(.a(\b[10] ), .b(\a[11] ), .out0(new_n137));
  nanb02aa1n06x5               g042(.a(new_n137), .b(new_n132), .out0(new_n138));
  xorc02aa1n12x5               g043(.a(\a[12] ), .b(\b[11] ), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nanp03aa1n02x5               g045(.a(new_n138), .b(new_n136), .c(new_n140), .o1(new_n141));
  tech160nm_fiaoi012aa1n04x5   g046(.a(new_n140), .b(new_n138), .c(new_n136), .o1(new_n142));
  norb02aa1n03x4               g047(.a(new_n141), .b(new_n142), .out0(\s[12] ));
  oao003aa1n02x5               g048(.a(new_n100), .b(new_n101), .c(new_n102), .carry(new_n144));
  nano23aa1n06x5               g049(.a(new_n106), .b(new_n105), .c(new_n107), .d(new_n104), .out0(new_n145));
  inv020aa1n02x5               g050(.a(new_n106), .o1(new_n146));
  oaoi03aa1n02x5               g051(.a(\a[4] ), .b(\b[3] ), .c(new_n146), .o1(new_n147));
  aoai13aa1n06x5               g052(.a(new_n120), .b(new_n147), .c(new_n144), .d(new_n145), .o1(new_n148));
  nano22aa1n03x5               g053(.a(new_n115), .b(new_n117), .c(new_n123), .out0(new_n149));
  nor003aa1n03x5               g054(.a(new_n149), .b(new_n121), .c(new_n111), .o1(new_n150));
  nona23aa1n02x4               g055(.a(new_n139), .b(new_n126), .c(new_n97), .d(new_n137), .out0(new_n151));
  inv040aa1d32x5               g056(.a(\a[12] ), .o1(new_n152));
  inv040aa1n18x5               g057(.a(\b[11] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(new_n153), .b(new_n152), .o1(new_n154));
  tech160nm_fioaoi03aa1n03p5x5 g059(.a(new_n129), .b(new_n130), .c(new_n98), .o1(new_n155));
  oaih22aa1n04x5               g060(.a(new_n134), .b(new_n135), .c(new_n153), .d(new_n152), .o1(new_n156));
  aoai13aa1n12x5               g061(.a(new_n154), .b(new_n156), .c(new_n155), .d(new_n136), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n151), .c(new_n148), .d(new_n150), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d28x5               g065(.a(\a[14] ), .o1(new_n161));
  nor042aa1d18x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  xorc02aa1n02x5               g067(.a(\a[13] ), .b(\b[12] ), .out0(new_n163));
  aoi012aa1n02x5               g068(.a(new_n162), .b(new_n159), .c(new_n163), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(new_n161), .out0(\s[14] ));
  nano23aa1n02x4               g070(.a(new_n97), .b(new_n137), .c(new_n139), .d(new_n126), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n125), .c(new_n110), .d(new_n120), .o1(new_n167));
  xorc02aa1n02x5               g072(.a(\a[14] ), .b(\b[13] ), .out0(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n163), .o1(new_n169));
  inv040aa1d32x5               g074(.a(\b[13] ), .o1(new_n170));
  oaoi03aa1n12x5               g075(.a(new_n161), .b(new_n170), .c(new_n162), .o1(new_n171));
  aoai13aa1n03x5               g076(.a(new_n171), .b(new_n169), .c(new_n167), .d(new_n158), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n12x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nand42aa1n16x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  xorc02aa1n02x5               g080(.a(\a[16] ), .b(\b[15] ), .out0(new_n176));
  aoi112aa1n02x5               g081(.a(new_n174), .b(new_n176), .c(new_n172), .d(new_n175), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n174), .o1(new_n178));
  inv000aa1d42x5               g083(.a(\a[13] ), .o1(new_n179));
  xroi22aa1d04x5               g084(.a(new_n179), .b(\b[12] ), .c(new_n161), .d(\b[13] ), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n171), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n175), .b(new_n174), .out0(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n181), .c(new_n159), .d(new_n180), .o1(new_n183));
  aobi12aa1n02x5               g088(.a(new_n176), .b(new_n183), .c(new_n178), .out0(new_n184));
  norp02aa1n02x5               g089(.a(new_n184), .b(new_n177), .o1(\s[16] ));
  nor002aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nand42aa1n04x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nano23aa1n06x5               g092(.a(new_n174), .b(new_n186), .c(new_n187), .d(new_n175), .out0(new_n188));
  norb02aa1n06x4               g093(.a(new_n188), .b(new_n169), .out0(new_n189));
  nand02aa1n02x5               g094(.a(new_n166), .b(new_n189), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n175), .o1(new_n191));
  oai022aa1n02x5               g096(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n192));
  oabi12aa1n09x5               g097(.a(new_n192), .b(new_n171), .c(new_n191), .out0(new_n193));
  aoi022aa1d18x5               g098(.a(new_n157), .b(new_n189), .c(new_n187), .d(new_n193), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n190), .c(new_n148), .d(new_n150), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g101(.a(\a[18] ), .o1(new_n197));
  norp02aa1n02x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  tech160nm_fiaoi012aa1n05x5   g104(.a(new_n198), .b(new_n195), .c(new_n199), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n197), .out0(\s[18] ));
  nano22aa1n03x7               g106(.a(new_n151), .b(new_n180), .c(new_n188), .out0(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n125), .c(new_n110), .d(new_n120), .o1(new_n203));
  inv000aa1d42x5               g108(.a(\a[17] ), .o1(new_n204));
  xroi22aa1d06x4               g109(.a(new_n204), .b(\b[16] ), .c(new_n197), .d(\b[17] ), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[17] ), .o1(new_n207));
  oao003aa1n02x5               g112(.a(new_n197), .b(new_n207), .c(new_n198), .carry(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n206), .c(new_n203), .d(new_n194), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n02x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand02aa1n03x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nor042aa1n02x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nand02aa1n03x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  aoi112aa1n02x5               g122(.a(new_n213), .b(new_n217), .c(new_n210), .d(new_n214), .o1(new_n218));
  inv000aa1d42x5               g123(.a(\b[18] ), .o1(new_n219));
  nanb02aa1n02x5               g124(.a(\a[19] ), .b(new_n219), .out0(new_n220));
  norb02aa1n02x5               g125(.a(new_n214), .b(new_n213), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n208), .c(new_n195), .d(new_n205), .o1(new_n222));
  aobi12aa1n03x5               g127(.a(new_n217), .b(new_n222), .c(new_n220), .out0(new_n223));
  nor002aa1n02x5               g128(.a(new_n223), .b(new_n218), .o1(\s[20] ));
  nanb03aa1n12x5               g129(.a(new_n215), .b(new_n216), .c(new_n214), .out0(new_n225));
  nona22aa1n03x5               g130(.a(new_n205), .b(new_n213), .c(new_n225), .out0(new_n226));
  nanp02aa1n02x5               g131(.a(\b[17] ), .b(\a[18] ), .o1(new_n227));
  oai022aa1n02x5               g132(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n228));
  nand03aa1n02x5               g133(.a(new_n228), .b(new_n220), .c(new_n227), .o1(new_n229));
  aoi012aa1n06x5               g134(.a(new_n215), .b(new_n213), .c(new_n216), .o1(new_n230));
  oai012aa1n18x5               g135(.a(new_n230), .b(new_n229), .c(new_n225), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n226), .c(new_n203), .d(new_n194), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[21] ), .b(\a[22] ), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoi112aa1n03x4               g144(.a(new_n235), .b(new_n239), .c(new_n233), .d(new_n237), .o1(new_n240));
  inv000aa1n03x5               g145(.a(new_n235), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n226), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n237), .b(new_n231), .c(new_n195), .d(new_n242), .o1(new_n243));
  aoi012aa1n03x5               g148(.a(new_n238), .b(new_n243), .c(new_n241), .o1(new_n244));
  norp02aa1n03x5               g149(.a(new_n244), .b(new_n240), .o1(\s[22] ));
  nor042aa1n06x5               g150(.a(new_n238), .b(new_n236), .o1(new_n246));
  nona23aa1d18x5               g151(.a(new_n205), .b(new_n246), .c(new_n225), .d(new_n213), .out0(new_n247));
  oao003aa1n02x5               g152(.a(\a[22] ), .b(\b[21] ), .c(new_n241), .carry(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoi012aa1n09x5               g154(.a(new_n249), .b(new_n231), .c(new_n246), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n247), .c(new_n203), .d(new_n194), .o1(new_n251));
  xorb03aa1n02x5               g156(.a(new_n251), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  tech160nm_fixorc02aa1n02p5x5 g158(.a(\a[23] ), .b(\b[22] ), .out0(new_n254));
  xorc02aa1n02x5               g159(.a(\a[24] ), .b(\b[23] ), .out0(new_n255));
  aoi112aa1n03x4               g160(.a(new_n253), .b(new_n255), .c(new_n251), .d(new_n254), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n253), .o1(new_n257));
  inv030aa1n02x5               g162(.a(new_n247), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n250), .o1(new_n259));
  aoai13aa1n04x5               g164(.a(new_n254), .b(new_n259), .c(new_n195), .d(new_n258), .o1(new_n260));
  aobi12aa1n03x5               g165(.a(new_n255), .b(new_n260), .c(new_n257), .out0(new_n261));
  norp02aa1n02x5               g166(.a(new_n261), .b(new_n256), .o1(\s[24] ));
  nano32aa1n03x7               g167(.a(new_n226), .b(new_n255), .c(new_n246), .d(new_n254), .out0(new_n263));
  inv000aa1n02x5               g168(.a(new_n263), .o1(new_n264));
  nano22aa1n02x4               g169(.a(new_n215), .b(new_n214), .c(new_n216), .out0(new_n265));
  oai012aa1n02x5               g170(.a(new_n227), .b(\b[18] ), .c(\a[19] ), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n228), .b(new_n266), .out0(new_n267));
  inv040aa1n02x5               g172(.a(new_n230), .o1(new_n268));
  aoai13aa1n06x5               g173(.a(new_n246), .b(new_n268), .c(new_n267), .d(new_n265), .o1(new_n269));
  and002aa1n02x5               g174(.a(new_n255), .b(new_n254), .o(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  oao003aa1n03x5               g176(.a(\a[24] ), .b(\b[23] ), .c(new_n257), .carry(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n271), .c(new_n269), .d(new_n248), .o1(new_n273));
  inv000aa1n02x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n264), .c(new_n203), .d(new_n194), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  xorc02aa1n03x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  xorc02aa1n03x5               g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  aoi112aa1n02x5               g184(.a(new_n277), .b(new_n279), .c(new_n275), .d(new_n278), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n277), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n278), .b(new_n273), .c(new_n195), .d(new_n263), .o1(new_n282));
  aobi12aa1n03x5               g187(.a(new_n279), .b(new_n282), .c(new_n281), .out0(new_n283));
  norp02aa1n03x5               g188(.a(new_n283), .b(new_n280), .o1(\s[26] ));
  tech160nm_fiaoi012aa1n03p5x5 g189(.a(new_n147), .b(new_n145), .c(new_n144), .o1(new_n285));
  nona22aa1n02x4               g190(.a(new_n122), .b(new_n119), .c(new_n118), .out0(new_n286));
  oai012aa1n03x5               g191(.a(new_n150), .b(new_n286), .c(new_n285), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(new_n157), .b(new_n189), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(new_n193), .b(new_n187), .o1(new_n289));
  nanp02aa1n02x5               g194(.a(new_n288), .b(new_n289), .o1(new_n290));
  and002aa1n02x5               g195(.a(new_n279), .b(new_n278), .o(new_n291));
  nano22aa1n12x5               g196(.a(new_n247), .b(new_n270), .c(new_n291), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n290), .c(new_n287), .d(new_n202), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[26] ), .b(\b[25] ), .c(new_n281), .carry(new_n294));
  aobi12aa1n12x5               g199(.a(new_n294), .b(new_n273), .c(new_n291), .out0(new_n295));
  xorc02aa1n12x5               g200(.a(\a[27] ), .b(\b[26] ), .out0(new_n296));
  xnbna2aa1n06x5               g201(.a(new_n296), .b(new_n295), .c(new_n293), .out0(\s[27] ));
  norp02aa1n02x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  inv040aa1n03x5               g203(.a(new_n298), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n296), .o1(new_n300));
  tech160nm_fiaoi012aa1n03p5x5 g205(.a(new_n300), .b(new_n295), .c(new_n293), .o1(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[27] ), .b(\a[28] ), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n301), .b(new_n299), .c(new_n302), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n270), .b(new_n249), .c(new_n231), .d(new_n246), .o1(new_n304));
  inv000aa1n02x5               g209(.a(new_n291), .o1(new_n305));
  aoai13aa1n04x5               g210(.a(new_n294), .b(new_n305), .c(new_n304), .d(new_n272), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n296), .b(new_n306), .c(new_n195), .d(new_n292), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n302), .b(new_n307), .c(new_n299), .o1(new_n308));
  norp02aa1n03x5               g213(.a(new_n308), .b(new_n303), .o1(\s[28] ));
  xnrc02aa1n02x5               g214(.a(\b[28] ), .b(\a[29] ), .out0(new_n310));
  norb02aa1n03x4               g215(.a(new_n296), .b(new_n302), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n306), .c(new_n195), .d(new_n292), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[28] ), .b(\b[27] ), .c(new_n299), .carry(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n310), .b(new_n312), .c(new_n313), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n311), .o1(new_n315));
  tech160nm_fiaoi012aa1n03p5x5 g220(.a(new_n315), .b(new_n295), .c(new_n293), .o1(new_n316));
  nano22aa1n03x5               g221(.a(new_n316), .b(new_n310), .c(new_n313), .out0(new_n317));
  norp02aa1n03x5               g222(.a(new_n314), .b(new_n317), .o1(\s[29] ));
  xorb03aa1n02x5               g223(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n03x5               g224(.a(new_n296), .b(new_n310), .c(new_n302), .out0(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n306), .c(new_n195), .d(new_n292), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .carry(new_n322));
  xnrc02aa1n02x5               g227(.a(\b[29] ), .b(\a[30] ), .out0(new_n323));
  tech160nm_fiaoi012aa1n02p5x5 g228(.a(new_n323), .b(new_n321), .c(new_n322), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n320), .o1(new_n325));
  tech160nm_fiaoi012aa1n03p5x5 g230(.a(new_n325), .b(new_n295), .c(new_n293), .o1(new_n326));
  nano22aa1n03x5               g231(.a(new_n326), .b(new_n322), .c(new_n323), .out0(new_n327));
  norp02aa1n03x5               g232(.a(new_n324), .b(new_n327), .o1(\s[30] ));
  norb02aa1n09x5               g233(.a(new_n320), .b(new_n323), .out0(new_n329));
  inv000aa1n02x5               g234(.a(new_n329), .o1(new_n330));
  tech160nm_fiaoi012aa1n03p5x5 g235(.a(new_n330), .b(new_n295), .c(new_n293), .o1(new_n331));
  oao003aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .c(new_n322), .carry(new_n332));
  xnrc02aa1n02x5               g237(.a(\b[30] ), .b(\a[31] ), .out0(new_n333));
  nano22aa1n03x5               g238(.a(new_n331), .b(new_n332), .c(new_n333), .out0(new_n334));
  aoai13aa1n02x5               g239(.a(new_n329), .b(new_n306), .c(new_n195), .d(new_n292), .o1(new_n335));
  tech160nm_fiaoi012aa1n02p5x5 g240(.a(new_n333), .b(new_n335), .c(new_n332), .o1(new_n336));
  norp02aa1n03x5               g241(.a(new_n336), .b(new_n334), .o1(\s[31] ));
  xnbna2aa1n03x5               g242(.a(new_n103), .b(new_n107), .c(new_n146), .out0(\s[3] ));
  norb02aa1n02x5               g243(.a(new_n104), .b(new_n105), .out0(new_n339));
  aoi112aa1n02x5               g244(.a(new_n106), .b(new_n339), .c(new_n144), .d(new_n107), .o1(new_n340));
  aoib12aa1n02x5               g245(.a(new_n340), .b(new_n110), .c(new_n105), .out0(\s[4] ));
  xnrb03aa1n02x5               g246(.a(new_n285), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g247(.a(new_n118), .o1(new_n343));
  oao003aa1n03x5               g248(.a(\a[5] ), .b(\b[4] ), .c(new_n285), .carry(new_n344));
  xnrc02aa1n02x5               g249(.a(new_n344), .b(new_n343), .out0(\s[6] ));
  norb02aa1n02x5               g250(.a(new_n113), .b(new_n114), .out0(new_n346));
  nanp02aa1n02x5               g251(.a(new_n344), .b(new_n343), .o1(new_n347));
  xobna2aa1n03x5               g252(.a(new_n346), .b(new_n347), .c(new_n117), .out0(\s[7] ));
  orn002aa1n02x5               g253(.a(\a[8] ), .b(\b[7] ), .o(new_n349));
  aoi013aa1n03x5               g254(.a(new_n114), .b(new_n347), .c(new_n117), .d(new_n113), .o1(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n350), .b(new_n349), .c(new_n112), .out0(\s[8] ));
  xnbna2aa1n03x5               g256(.a(new_n126), .b(new_n148), .c(new_n150), .out0(\s[9] ));
endmodule


