// Benchmark "adder" written by ABC on Thu Jul 18 15:06:29 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n312, new_n315, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[6] ), .b(\a[7] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  oaoi03aa1n02x5               g003(.a(\a[8] ), .b(\b[7] ), .c(new_n98), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[6] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[5] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[4] ), .b(\a[5] ), .o1(new_n102));
  oaoi03aa1n02x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  norp02aa1n04x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  nand02aa1n03x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nand02aa1d28x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n105), .b(new_n106), .c(new_n97), .d(new_n104), .out0(new_n107));
  oabi12aa1n06x5               g012(.a(new_n99), .b(new_n107), .c(new_n103), .out0(new_n108));
  inv040aa1d32x5               g013(.a(\a[4] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[3] ), .o1(new_n110));
  nand22aa1n03x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(new_n111), .b(new_n112), .o1(new_n113));
  norp02aa1n04x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  oaoi03aa1n02x5               g019(.a(new_n109), .b(new_n110), .c(new_n114), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nanb02aa1n06x5               g021(.a(new_n114), .b(new_n116), .out0(new_n117));
  nand42aa1n03x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  nand02aa1d04x5               g023(.a(\b[0] ), .b(\a[1] ), .o1(new_n119));
  nor042aa1n02x5               g024(.a(\b[1] ), .b(\a[2] ), .o1(new_n120));
  oai012aa1n12x5               g025(.a(new_n118), .b(new_n120), .c(new_n119), .o1(new_n121));
  oai013aa1n09x5               g026(.a(new_n115), .b(new_n121), .c(new_n117), .d(new_n113), .o1(new_n122));
  xnrc02aa1n02x5               g027(.a(\b[5] ), .b(\a[6] ), .out0(new_n123));
  nanp02aa1n02x5               g028(.a(\b[4] ), .b(\a[5] ), .o1(new_n124));
  nanb02aa1n02x5               g029(.a(new_n102), .b(new_n124), .out0(new_n125));
  nor043aa1n04x5               g030(.a(new_n107), .b(new_n125), .c(new_n123), .o1(new_n126));
  aoi012aa1n02x5               g031(.a(new_n108), .b(new_n122), .c(new_n126), .o1(new_n127));
  oaoi03aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .c(new_n127), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n04x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  norp02aa1n02x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nand02aa1n02x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  aoi012aa1n03x5               g037(.a(new_n131), .b(new_n130), .c(new_n132), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[8] ), .b(\a[9] ), .o1(new_n134));
  nano23aa1n06x5               g039(.a(new_n130), .b(new_n131), .c(new_n132), .d(new_n134), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n108), .c(new_n122), .d(new_n126), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(new_n136), .b(new_n133), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g043(.a(\a[12] ), .o1(new_n139));
  nor042aa1n03x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nand42aa1n03x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  aoi012aa1n02x5               g046(.a(new_n140), .b(new_n137), .c(new_n141), .o1(new_n142));
  xorb03aa1n02x5               g047(.a(new_n142), .b(\b[11] ), .c(new_n139), .out0(\s[12] ));
  nor042aa1n02x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanp02aa1n03x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  ao0012aa1n03x7               g050(.a(new_n144), .b(new_n140), .c(new_n145), .o(new_n146));
  nano23aa1n06x5               g051(.a(new_n140), .b(new_n144), .c(new_n145), .d(new_n141), .out0(new_n147));
  aoib12aa1n02x5               g052(.a(new_n146), .b(new_n147), .c(new_n133), .out0(new_n148));
  nona23aa1n09x5               g053(.a(new_n145), .b(new_n141), .c(new_n140), .d(new_n144), .out0(new_n149));
  norb02aa1n02x5               g054(.a(new_n135), .b(new_n149), .out0(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n108), .c(new_n122), .d(new_n126), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n151), .b(new_n148), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g058(.a(\a[14] ), .o1(new_n154));
  nor042aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n06x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n155), .b(new_n152), .c(new_n156), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[13] ), .c(new_n154), .out0(\s[14] ));
  nor042aa1n02x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nand42aa1n03x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nona23aa1n02x4               g065(.a(new_n160), .b(new_n156), .c(new_n155), .d(new_n159), .out0(new_n161));
  oabi12aa1n06x5               g066(.a(new_n146), .b(new_n149), .c(new_n133), .out0(new_n162));
  aoi012aa1n02x5               g067(.a(new_n159), .b(new_n155), .c(new_n160), .o1(new_n163));
  nano23aa1n03x7               g068(.a(new_n155), .b(new_n159), .c(new_n160), .d(new_n156), .out0(new_n164));
  aobi12aa1n02x5               g069(.a(new_n163), .b(new_n162), .c(new_n164), .out0(new_n165));
  oai012aa1n02x5               g070(.a(new_n165), .b(new_n151), .c(new_n161), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n03x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  norp02aa1n04x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand42aa1n03x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n168), .b(new_n172), .c(new_n166), .d(new_n169), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(\s[16] ));
  nanb02aa1n02x5               g080(.a(new_n168), .b(new_n169), .out0(new_n176));
  aoi012aa1n02x5               g081(.a(new_n170), .b(new_n168), .c(new_n171), .o1(new_n177));
  oai013aa1n02x4               g082(.a(new_n177), .b(new_n163), .c(new_n176), .d(new_n172), .o1(new_n178));
  nano23aa1n03x5               g083(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n179));
  nanp02aa1n03x5               g084(.a(new_n179), .b(new_n164), .o1(new_n180));
  aoib12aa1n12x5               g085(.a(new_n178), .b(new_n162), .c(new_n180), .out0(new_n181));
  nano22aa1n03x7               g086(.a(new_n180), .b(new_n135), .c(new_n147), .out0(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n108), .c(new_n122), .d(new_n126), .o1(new_n183));
  xorc02aa1n12x5               g088(.a(\a[17] ), .b(\b[16] ), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n183), .c(new_n181), .out0(\s[17] ));
  nanp02aa1n06x5               g090(.a(new_n183), .b(new_n181), .o1(new_n186));
  nor042aa1n06x5               g091(.a(\b[16] ), .b(\a[17] ), .o1(new_n187));
  tech160nm_fiaoi012aa1n05x5   g092(.a(new_n187), .b(new_n186), .c(new_n184), .o1(new_n188));
  inv030aa1d32x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[17] ), .o1(new_n190));
  nand42aa1n06x5               g095(.a(new_n190), .b(new_n189), .o1(new_n191));
  nand02aa1d28x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n188), .b(new_n192), .c(new_n191), .out0(\s[18] ));
  aob012aa1d18x5               g098(.a(new_n191), .b(new_n187), .c(new_n192), .out0(new_n194));
  inv000aa1d42x5               g099(.a(new_n194), .o1(new_n195));
  inv000aa1n09x5               g100(.a(new_n184), .o1(new_n196));
  nano22aa1d15x5               g101(.a(new_n196), .b(new_n191), .c(new_n192), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n195), .b(new_n198), .c(new_n183), .d(new_n181), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1n03x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nor042aa1n09x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand02aa1d12x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  norb02aa1n12x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n199), .d(new_n203), .o1(new_n208));
  norb02aa1n06x4               g113(.a(new_n203), .b(new_n202), .out0(new_n209));
  nanp02aa1n02x5               g114(.a(new_n199), .b(new_n209), .o1(new_n210));
  nona22aa1n02x4               g115(.a(new_n210), .b(new_n207), .c(new_n202), .out0(new_n211));
  nanp02aa1n02x5               g116(.a(new_n211), .b(new_n208), .o1(\s[20] ));
  aoi012aa1d24x5               g117(.a(new_n204), .b(new_n202), .c(new_n205), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nano23aa1n06x5               g119(.a(new_n202), .b(new_n204), .c(new_n205), .d(new_n203), .out0(new_n215));
  aoi012aa1n02x5               g120(.a(new_n214), .b(new_n215), .c(new_n194), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(new_n197), .b(new_n215), .o1(new_n217));
  aoai13aa1n06x5               g122(.a(new_n216), .b(new_n217), .c(new_n183), .d(new_n181), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  nand42aa1d28x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  nor002aa1n06x5               g127(.a(\b[21] ), .b(\a[22] ), .o1(new_n223));
  nand02aa1d24x5               g128(.a(\b[21] ), .b(\a[22] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoai13aa1n02x5               g131(.a(new_n226), .b(new_n220), .c(new_n218), .d(new_n222), .o1(new_n227));
  nanp02aa1n02x5               g132(.a(new_n218), .b(new_n222), .o1(new_n228));
  nona22aa1n02x4               g133(.a(new_n228), .b(new_n226), .c(new_n220), .out0(new_n229));
  nanp02aa1n02x5               g134(.a(new_n229), .b(new_n227), .o1(\s[22] ));
  nanp03aa1d12x5               g135(.a(new_n194), .b(new_n209), .c(new_n206), .o1(new_n231));
  nanp02aa1n02x5               g136(.a(new_n231), .b(new_n213), .o1(new_n232));
  ao0012aa1n03x7               g137(.a(new_n223), .b(new_n220), .c(new_n224), .o(new_n233));
  nano23aa1d12x5               g138(.a(new_n220), .b(new_n223), .c(new_n224), .d(new_n221), .out0(new_n234));
  aoi012aa1n02x5               g139(.a(new_n233), .b(new_n232), .c(new_n234), .o1(new_n235));
  nanp03aa1n02x5               g140(.a(new_n197), .b(new_n215), .c(new_n234), .o1(new_n236));
  aoai13aa1n06x5               g141(.a(new_n235), .b(new_n236), .c(new_n183), .d(new_n181), .o1(new_n237));
  xorb03aa1n02x5               g142(.a(new_n237), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  nand02aa1n16x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  nor042aa1n06x5               g146(.a(\b[23] ), .b(\a[24] ), .o1(new_n242));
  nand02aa1d16x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  nanb02aa1n02x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n239), .c(new_n237), .d(new_n241), .o1(new_n245));
  nanp02aa1n02x5               g150(.a(new_n237), .b(new_n241), .o1(new_n246));
  nona22aa1n02x4               g151(.a(new_n246), .b(new_n244), .c(new_n239), .out0(new_n247));
  nanp02aa1n02x5               g152(.a(new_n247), .b(new_n245), .o1(\s[24] ));
  ao0012aa1n03x5               g153(.a(new_n242), .b(new_n239), .c(new_n243), .o(new_n249));
  nano23aa1d15x5               g154(.a(new_n239), .b(new_n242), .c(new_n243), .d(new_n240), .out0(new_n250));
  aoi012aa1n06x5               g155(.a(new_n249), .b(new_n250), .c(new_n233), .o1(new_n251));
  nand22aa1n09x5               g156(.a(new_n250), .b(new_n234), .o1(new_n252));
  aoai13aa1n12x5               g157(.a(new_n251), .b(new_n252), .c(new_n231), .d(new_n213), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  nanb03aa1n02x5               g159(.a(new_n252), .b(new_n197), .c(new_n215), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n254), .b(new_n255), .c(new_n183), .d(new_n181), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  tech160nm_fixorc02aa1n03p5x5 g163(.a(\a[25] ), .b(\b[24] ), .out0(new_n259));
  tech160nm_fixnrc02aa1n04x5   g164(.a(\b[25] ), .b(\a[26] ), .out0(new_n260));
  aoai13aa1n02x5               g165(.a(new_n260), .b(new_n258), .c(new_n256), .d(new_n259), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(new_n256), .b(new_n259), .o1(new_n262));
  nona22aa1n02x4               g167(.a(new_n262), .b(new_n260), .c(new_n258), .out0(new_n263));
  nanp02aa1n03x5               g168(.a(new_n263), .b(new_n261), .o1(\s[26] ));
  inv000aa1d42x5               g169(.a(\a[26] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(\b[25] ), .o1(new_n266));
  oaoi03aa1n12x5               g171(.a(new_n265), .b(new_n266), .c(new_n258), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  norb02aa1n02x7               g173(.a(new_n259), .b(new_n260), .out0(new_n269));
  tech160nm_fiaoi012aa1n05x5   g174(.a(new_n268), .b(new_n253), .c(new_n269), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n252), .o1(new_n271));
  nanb03aa1n02x5               g176(.a(new_n217), .b(new_n269), .c(new_n271), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n270), .b(new_n272), .c(new_n183), .d(new_n181), .o1(new_n273));
  xorb03aa1n03x5               g178(.a(new_n273), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g179(.a(\b[26] ), .b(\a[27] ), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  xnrc02aa1n02x5               g181(.a(\b[27] ), .b(\a[28] ), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .d(new_n276), .o1(new_n278));
  nand22aa1n03x5               g183(.a(new_n253), .b(new_n269), .o1(new_n279));
  nanp02aa1n03x5               g184(.a(new_n279), .b(new_n267), .o1(new_n280));
  nano32aa1n03x7               g185(.a(new_n217), .b(new_n269), .c(new_n234), .d(new_n250), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n276), .b(new_n280), .c(new_n186), .d(new_n281), .o1(new_n282));
  nona22aa1n03x5               g187(.a(new_n282), .b(new_n277), .c(new_n275), .out0(new_n283));
  nanp02aa1n03x5               g188(.a(new_n278), .b(new_n283), .o1(\s[28] ));
  inv000aa1d42x5               g189(.a(\a[28] ), .o1(new_n285));
  inv000aa1d42x5               g190(.a(\b[27] ), .o1(new_n286));
  oaoi03aa1n09x5               g191(.a(new_n285), .b(new_n286), .c(new_n275), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  norb02aa1n02x5               g193(.a(new_n276), .b(new_n277), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n280), .c(new_n186), .d(new_n281), .o1(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  nona22aa1n03x5               g196(.a(new_n290), .b(new_n291), .c(new_n288), .out0(new_n292));
  aoai13aa1n03x5               g197(.a(new_n291), .b(new_n288), .c(new_n273), .d(new_n289), .o1(new_n293));
  nanp02aa1n03x5               g198(.a(new_n293), .b(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n119), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  tech160nm_fioaoi03aa1n03p5x5 g200(.a(\a[29] ), .b(\b[28] ), .c(new_n287), .o1(new_n296));
  norb03aa1n02x5               g201(.a(new_n276), .b(new_n291), .c(new_n277), .out0(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[29] ), .b(\a[30] ), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n296), .c(new_n273), .d(new_n297), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n297), .b(new_n280), .c(new_n186), .d(new_n281), .o1(new_n300));
  nona22aa1n03x5               g205(.a(new_n300), .b(new_n298), .c(new_n296), .out0(new_n301));
  nanp02aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[30] ));
  nanb02aa1n02x5               g207(.a(new_n298), .b(new_n296), .out0(new_n303));
  oai012aa1n02x5               g208(.a(new_n303), .b(\b[29] ), .c(\a[30] ), .o1(new_n304));
  norb02aa1n02x5               g209(.a(new_n297), .b(new_n298), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n280), .c(new_n186), .d(new_n281), .o1(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  nona22aa1n03x5               g212(.a(new_n306), .b(new_n307), .c(new_n304), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n307), .b(new_n304), .c(new_n273), .d(new_n305), .o1(new_n309));
  nanp02aa1n03x5               g214(.a(new_n309), .b(new_n308), .o1(\s[31] ));
  xnrb03aa1n02x5               g215(.a(new_n121), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g216(.a(\a[3] ), .b(\b[2] ), .c(new_n121), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g218(.a(new_n122), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioai012aa1n05x5   g219(.a(new_n124), .b(new_n122), .c(new_n102), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[5] ), .c(new_n100), .out0(\s[6] ));
  and002aa1n02x5               g221(.a(\b[5] ), .b(\a[6] ), .o(new_n317));
  inv000aa1d42x5               g222(.a(new_n106), .o1(new_n318));
  nanb02aa1n02x5               g223(.a(new_n123), .b(new_n315), .out0(new_n319));
  nona32aa1n03x5               g224(.a(new_n319), .b(new_n318), .c(new_n317), .d(new_n97), .out0(new_n320));
  aboi22aa1n03x5               g225(.a(new_n317), .b(new_n319), .c(new_n98), .d(new_n106), .out0(new_n321));
  norb02aa1n02x5               g226(.a(new_n320), .b(new_n321), .out0(\s[7] ));
  norb02aa1n02x5               g227(.a(new_n105), .b(new_n104), .out0(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n323), .b(new_n320), .c(new_n98), .out0(\s[8] ));
  xnrb03aa1n02x5               g229(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


