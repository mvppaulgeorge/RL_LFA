// Benchmark "adder" written by ABC on Wed Jul 17 22:21:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n328, new_n330, new_n333,
    new_n334, new_n335, new_n337, new_n338, new_n339, new_n340, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand22aa1n09x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n09x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1n16x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[3] ), .o1(new_n102));
  oai022aa1n02x5               g007(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  oaib12aa1n06x5               g008(.a(new_n103), .b(new_n102), .c(\a[4] ), .out0(new_n104));
  inv000aa1d42x5               g009(.a(\a[4] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(new_n102), .b(new_n105), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nor042aa1n04x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  oai112aa1n06x5               g014(.a(new_n106), .b(new_n107), .c(new_n109), .d(new_n108), .o1(new_n110));
  orn002aa1n24x5               g015(.a(\a[3] ), .b(\b[2] ), .o(new_n111));
  tech160nm_finand02aa1n03p5x5 g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  oai112aa1n06x5               g017(.a(new_n111), .b(new_n112), .c(new_n102), .d(new_n105), .o1(new_n113));
  oai012aa1n18x5               g018(.a(new_n104), .b(new_n110), .c(new_n113), .o1(new_n114));
  nor042aa1n06x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand42aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor042aa1n04x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  tech160nm_finand02aa1n03p5x5 g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nona23aa1n09x5               g023(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n119));
  nor002aa1n02x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nand42aa1n04x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nor042aa1n06x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  nand42aa1n04x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nona23aa1n09x5               g028(.a(new_n123), .b(new_n121), .c(new_n120), .d(new_n122), .out0(new_n124));
  nor042aa1n04x5               g029(.a(new_n124), .b(new_n119), .o1(new_n125));
  nanb03aa1n03x5               g030(.a(new_n122), .b(new_n123), .c(new_n121), .out0(new_n126));
  oai122aa1n06x5               g031(.a(new_n116), .b(new_n115), .c(new_n117), .d(\b[7] ), .e(\a[8] ), .o1(new_n127));
  tech160nm_fiaoi012aa1n03p5x5 g032(.a(new_n120), .b(new_n122), .c(new_n121), .o1(new_n128));
  oai012aa1n04x7               g033(.a(new_n128), .b(new_n127), .c(new_n126), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n129), .c(new_n114), .d(new_n125), .o1(new_n131));
  xobna2aa1n03x5               g036(.a(new_n99), .b(new_n131), .c(new_n101), .out0(\s[10] ));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1n08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  nona22aa1n06x5               g040(.a(new_n131), .b(new_n100), .c(new_n97), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n135), .b(new_n136), .c(new_n98), .out0(\s[11] ));
  nor002aa1d32x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  nand22aa1n09x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  aoi013aa1n06x4               g045(.a(new_n133), .b(new_n136), .c(new_n134), .d(new_n98), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n139), .c(new_n140), .out0(\s[12] ));
  nona23aa1n09x5               g047(.a(new_n140), .b(new_n134), .c(new_n133), .d(new_n138), .out0(new_n143));
  norb03aa1n06x5               g048(.a(new_n130), .b(new_n143), .c(new_n99), .out0(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n129), .c(new_n114), .d(new_n125), .o1(new_n145));
  nanb03aa1n06x5               g050(.a(new_n138), .b(new_n140), .c(new_n134), .out0(new_n146));
  inv000aa1n02x5               g051(.a(new_n133), .o1(new_n147));
  oai112aa1n06x5               g052(.a(new_n147), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n148));
  aoi012aa1n06x5               g053(.a(new_n138), .b(new_n133), .c(new_n140), .o1(new_n149));
  oai012aa1n02x5               g054(.a(new_n149), .b(new_n148), .c(new_n146), .o1(new_n150));
  inv020aa1n02x5               g055(.a(new_n150), .o1(new_n151));
  nor002aa1d32x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nanp02aa1n06x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanb02aa1n02x5               g058(.a(new_n152), .b(new_n153), .out0(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  xnbna2aa1n03x5               g060(.a(new_n155), .b(new_n145), .c(new_n151), .out0(\s[13] ));
  orn002aa1n24x5               g061(.a(\a[13] ), .b(\b[12] ), .o(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n154), .c(new_n145), .d(new_n151), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n16x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nanp02aa1n04x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nona23aa1d24x5               g066(.a(new_n161), .b(new_n153), .c(new_n152), .d(new_n160), .out0(new_n162));
  oaoi03aa1n12x5               g067(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n163));
  inv030aa1n02x5               g068(.a(new_n163), .o1(new_n164));
  aoai13aa1n04x5               g069(.a(new_n164), .b(new_n162), .c(new_n145), .d(new_n151), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  xnrc02aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  xnrc02aa1n02x5               g074(.a(\b[15] ), .b(\a[16] ), .out0(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n167), .c(new_n165), .d(new_n169), .o1(new_n171));
  aoi112aa1n02x7               g076(.a(new_n167), .b(new_n170), .c(new_n165), .d(new_n169), .o1(new_n172));
  nanb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(\s[16] ));
  nand42aa1n08x5               g078(.a(new_n114), .b(new_n125), .o1(new_n174));
  tech160nm_ficinv00aa1n08x5   g079(.clk(new_n129), .clkout(new_n175));
  nand42aa1n04x5               g080(.a(new_n174), .b(new_n175), .o1(new_n176));
  nona32aa1n09x5               g081(.a(new_n144), .b(new_n170), .c(new_n168), .d(new_n162), .out0(new_n177));
  nanb02aa1n06x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  nor022aa1n03x5               g083(.a(new_n170), .b(new_n168), .o1(new_n179));
  oaoi13aa1n09x5               g084(.a(new_n162), .b(new_n149), .c(new_n148), .d(new_n146), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\a[16] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\b[15] ), .o1(new_n182));
  oao003aa1n06x5               g087(.a(new_n181), .b(new_n182), .c(new_n167), .carry(new_n183));
  oaoi13aa1n09x5               g088(.a(new_n183), .b(new_n179), .c(new_n180), .d(new_n163), .o1(new_n184));
  nor002aa1d32x5               g089(.a(\b[16] ), .b(\a[17] ), .o1(new_n185));
  nand42aa1n04x5               g090(.a(\b[16] ), .b(\a[17] ), .o1(new_n186));
  norb02aa1n02x5               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n184), .c(new_n178), .out0(\s[17] ));
  aoi012aa1d18x5               g093(.a(new_n177), .b(new_n174), .c(new_n175), .o1(new_n189));
  inv000aa1n04x5               g094(.a(new_n179), .o1(new_n190));
  nano22aa1n02x4               g095(.a(new_n138), .b(new_n134), .c(new_n140), .out0(new_n191));
  oai012aa1n02x5               g096(.a(new_n98), .b(\b[10] ), .c(\a[11] ), .o1(new_n192));
  oab012aa1n04x5               g097(.a(new_n192), .b(new_n97), .c(new_n100), .out0(new_n193));
  inv040aa1n03x5               g098(.a(new_n149), .o1(new_n194));
  inv000aa1n02x5               g099(.a(new_n162), .o1(new_n195));
  aoai13aa1n04x5               g100(.a(new_n195), .b(new_n194), .c(new_n193), .d(new_n191), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n183), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n190), .c(new_n196), .d(new_n164), .o1(new_n198));
  oaoi13aa1n06x5               g103(.a(new_n185), .b(new_n187), .c(new_n198), .d(new_n189), .o1(new_n199));
  xnrb03aa1n03x5               g104(.a(new_n199), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor002aa1d32x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand02aa1d24x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nano23aa1d15x5               g107(.a(new_n185), .b(new_n201), .c(new_n202), .d(new_n186), .out0(new_n203));
  oai012aa1n06x5               g108(.a(new_n203), .b(new_n198), .c(new_n189), .o1(new_n204));
  oa0012aa1n02x5               g109(.a(new_n202), .b(new_n201), .c(new_n185), .o(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  nor042aa1d18x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nanp02aa1n09x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n03x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n204), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g116(.a(new_n204), .b(new_n206), .o1(new_n212));
  nor002aa1d32x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d28x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n207), .c(new_n212), .d(new_n208), .o1(new_n216));
  aoi012aa1n06x5               g121(.a(new_n129), .b(new_n114), .c(new_n125), .o1(new_n217));
  oai012aa1n06x5               g122(.a(new_n184), .b(new_n177), .c(new_n217), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n209), .b(new_n205), .c(new_n218), .d(new_n203), .o1(new_n219));
  nona22aa1n02x5               g124(.a(new_n219), .b(new_n215), .c(new_n207), .out0(new_n220));
  nanp02aa1n03x5               g125(.a(new_n216), .b(new_n220), .o1(\s[20] ));
  nano22aa1n03x7               g126(.a(new_n215), .b(new_n203), .c(new_n209), .out0(new_n222));
  inv000aa1n02x5               g127(.a(new_n222), .o1(new_n223));
  nanb03aa1n09x5               g128(.a(new_n213), .b(new_n214), .c(new_n208), .out0(new_n224));
  oai122aa1n12x5               g129(.a(new_n202), .b(new_n201), .c(new_n185), .d(\b[18] ), .e(\a[19] ), .o1(new_n225));
  aoi012aa1d18x5               g130(.a(new_n213), .b(new_n207), .c(new_n214), .o1(new_n226));
  oai012aa1d24x5               g131(.a(new_n226), .b(new_n225), .c(new_n224), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n02x7               g133(.a(new_n228), .b(new_n223), .c(new_n178), .d(new_n184), .o1(new_n229));
  nor002aa1d32x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand42aa1n16x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  aoi112aa1n02x5               g137(.a(new_n232), .b(new_n227), .c(new_n218), .d(new_n222), .o1(new_n233));
  aoi012aa1n02x5               g138(.a(new_n233), .b(new_n229), .c(new_n232), .o1(\s[21] ));
  nor002aa1n16x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  nand42aa1n10x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  nanb02aa1n02x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n230), .c(new_n229), .d(new_n232), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n232), .b(new_n227), .c(new_n218), .d(new_n222), .o1(new_n239));
  nona22aa1n02x5               g144(.a(new_n239), .b(new_n237), .c(new_n230), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n238), .b(new_n240), .o1(\s[22] ));
  nano23aa1d15x5               g146(.a(new_n230), .b(new_n235), .c(new_n236), .d(new_n231), .out0(new_n242));
  nano32aa1n03x7               g147(.a(new_n215), .b(new_n242), .c(new_n203), .d(new_n209), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  oa0012aa1n06x5               g149(.a(new_n236), .b(new_n235), .c(new_n230), .o(new_n245));
  aoi012aa1d18x5               g150(.a(new_n245), .b(new_n227), .c(new_n242), .o1(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n244), .c(new_n178), .d(new_n184), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  tech160nm_fixnrc02aa1n05x5   g155(.a(\b[23] ), .b(\a[24] ), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n249), .c(new_n247), .d(new_n250), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n246), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n250), .b(new_n253), .c(new_n218), .d(new_n243), .o1(new_n254));
  nona22aa1n02x5               g159(.a(new_n254), .b(new_n251), .c(new_n249), .out0(new_n255));
  nanp02aa1n03x5               g160(.a(new_n252), .b(new_n255), .o1(\s[24] ));
  norb02aa1n06x4               g161(.a(new_n250), .b(new_n251), .out0(new_n257));
  nano22aa1n03x7               g162(.a(new_n223), .b(new_n257), .c(new_n242), .out0(new_n258));
  oai012aa1n06x5               g163(.a(new_n258), .b(new_n198), .c(new_n189), .o1(new_n259));
  nano22aa1n03x5               g164(.a(new_n213), .b(new_n208), .c(new_n214), .out0(new_n260));
  tech160nm_fioai012aa1n04x5   g165(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .o1(new_n261));
  oab012aa1n03x5               g166(.a(new_n261), .b(new_n185), .c(new_n201), .out0(new_n262));
  inv020aa1n03x5               g167(.a(new_n226), .o1(new_n263));
  aoai13aa1n06x5               g168(.a(new_n242), .b(new_n263), .c(new_n262), .d(new_n260), .o1(new_n264));
  inv040aa1n02x5               g169(.a(new_n245), .o1(new_n265));
  inv020aa1n04x5               g170(.a(new_n257), .o1(new_n266));
  oai022aa1n02x5               g171(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n267));
  aob012aa1n02x5               g172(.a(new_n267), .b(\b[23] ), .c(\a[24] ), .out0(new_n268));
  aoai13aa1n12x5               g173(.a(new_n268), .b(new_n266), .c(new_n264), .d(new_n265), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  xnbna2aa1n03x5               g176(.a(new_n271), .b(new_n259), .c(new_n270), .out0(\s[25] ));
  tech160nm_finand02aa1n03p5x5 g177(.a(new_n259), .b(new_n270), .o1(new_n273));
  norp02aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  tech160nm_fixnrc02aa1n04x5   g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n274), .c(new_n273), .d(new_n271), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n271), .b(new_n269), .c(new_n218), .d(new_n258), .o1(new_n277));
  nona22aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n274), .out0(new_n278));
  nanp02aa1n03x5               g183(.a(new_n276), .b(new_n278), .o1(\s[26] ));
  norb02aa1n12x5               g184(.a(new_n271), .b(new_n275), .out0(new_n280));
  nano32aa1n06x5               g185(.a(new_n223), .b(new_n280), .c(new_n242), .d(new_n257), .out0(new_n281));
  oai012aa1n12x5               g186(.a(new_n281), .b(new_n198), .c(new_n189), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(\b[25] ), .b(\a[26] ), .o1(new_n283));
  oai022aa1n02x5               g188(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n284));
  aoi022aa1n12x5               g189(.a(new_n269), .b(new_n280), .c(new_n283), .d(new_n284), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n282), .c(new_n285), .out0(\s[27] ));
  xorc02aa1n12x5               g192(.a(\a[28] ), .b(\b[27] ), .out0(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  inv000aa1n03x5               g195(.a(new_n290), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n286), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n291), .b(new_n292), .c(new_n282), .d(new_n285), .o1(new_n293));
  nanp02aa1n03x5               g198(.a(new_n293), .b(new_n289), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n257), .b(new_n245), .c(new_n227), .d(new_n242), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n280), .o1(new_n296));
  nanp02aa1n02x5               g201(.a(new_n284), .b(new_n283), .o1(new_n297));
  aoai13aa1n06x5               g202(.a(new_n297), .b(new_n296), .c(new_n295), .d(new_n268), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n286), .b(new_n298), .c(new_n218), .d(new_n281), .o1(new_n299));
  nona22aa1n02x5               g204(.a(new_n299), .b(new_n289), .c(new_n290), .out0(new_n300));
  nanp02aa1n03x5               g205(.a(new_n294), .b(new_n300), .o1(\s[28] ));
  and002aa1n02x5               g206(.a(new_n288), .b(new_n286), .o(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n298), .c(new_n218), .d(new_n281), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n302), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[28] ), .b(\b[27] ), .c(new_n291), .carry(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n304), .c(new_n282), .d(new_n285), .o1(new_n306));
  tech160nm_fixorc02aa1n02p5x5 g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g215(.a(new_n289), .b(new_n286), .c(new_n307), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n298), .c(new_n218), .d(new_n281), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  oaoi03aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .o1(new_n314));
  inv000aa1n03x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n282), .d(new_n285), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .out0(new_n317));
  norp02aa1n02x5               g222(.a(new_n314), .b(new_n317), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n312), .d(new_n318), .o1(\s[30] ));
  nano32aa1n09x5               g224(.a(new_n292), .b(new_n317), .c(new_n288), .d(new_n307), .out0(new_n320));
  aoai13aa1n02x5               g225(.a(new_n320), .b(new_n298), .c(new_n218), .d(new_n281), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  inv000aa1d42x5               g229(.a(new_n320), .o1(new_n325));
  aoai13aa1n03x5               g230(.a(new_n323), .b(new_n325), .c(new_n282), .d(new_n285), .o1(new_n326));
  aoi022aa1n03x5               g231(.a(new_n326), .b(new_n322), .c(new_n321), .d(new_n324), .o1(\s[31] ));
  oai012aa1n02x5               g232(.a(new_n107), .b(new_n109), .c(new_n108), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n111), .c(new_n112), .out0(\s[3] ));
  oaoi03aa1n02x5               g234(.a(\a[3] ), .b(\b[2] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g236(.a(new_n114), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g237(.a(new_n115), .b(new_n116), .out0(new_n333));
  norb02aa1n02x5               g238(.a(new_n118), .b(new_n117), .out0(new_n334));
  oai112aa1n02x5               g239(.a(new_n104), .b(new_n334), .c(new_n110), .d(new_n113), .o1(new_n335));
  xnbna2aa1n03x5               g240(.a(new_n333), .b(new_n335), .c(new_n118), .out0(\s[6] ));
  nanb02aa1n02x5               g241(.a(new_n122), .b(new_n123), .out0(new_n337));
  aoai13aa1n02x5               g242(.a(new_n116), .b(new_n115), .c(new_n335), .d(new_n118), .o1(new_n338));
  aoi012aa1n02x5               g243(.a(new_n333), .b(new_n335), .c(new_n118), .o1(new_n339));
  nano23aa1n02x4               g244(.a(new_n339), .b(new_n122), .c(new_n116), .d(new_n123), .out0(new_n340));
  aoi012aa1n02x5               g245(.a(new_n340), .b(new_n337), .c(new_n338), .o1(\s[7] ));
  norp02aa1n02x5               g246(.a(new_n340), .b(new_n122), .o1(new_n342));
  xnrb03aa1n02x5               g247(.a(new_n342), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g248(.a(new_n130), .b(new_n174), .c(new_n175), .out0(\s[9] ));
endmodule


