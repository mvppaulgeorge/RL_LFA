// Benchmark "adder" written by ABC on Thu Jul 18 03:40:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n348, new_n349, new_n351, new_n352,
    new_n354, new_n355, new_n356, new_n357, new_n359, new_n360, new_n361,
    new_n363, new_n365, new_n366, new_n367, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\a[3] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[4] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[2] ), .o1(new_n100));
  aboi22aa1n03x5               g005(.a(\b[3] ), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n101));
  nanp02aa1n02x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  oab012aa1n06x5               g007(.a(new_n102), .b(\a[2] ), .c(\b[1] ), .out0(new_n103));
  nand42aa1n02x5               g008(.a(new_n100), .b(new_n98), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand23aa1n03x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  tech160nm_fioai012aa1n05x5   g012(.a(new_n101), .b(new_n107), .c(new_n103), .o1(new_n108));
  nor042aa1n04x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(new_n109), .o1(new_n110));
  nor042aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  aoi012aa1n02x5               g016(.a(new_n111), .b(\a[6] ), .c(\b[5] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[7] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[6] ), .o1(new_n114));
  aoi022aa1n02x5               g019(.a(new_n114), .b(new_n113), .c(\a[8] ), .d(\b[7] ), .o1(new_n115));
  aoi022aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nor042aa1n06x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(new_n118), .o1(new_n119));
  nanp03aa1n02x5               g024(.a(new_n116), .b(new_n119), .c(new_n117), .o1(new_n120));
  nano32aa1n03x7               g025(.a(new_n120), .b(new_n115), .c(new_n112), .d(new_n110), .out0(new_n121));
  nand02aa1d04x5               g026(.a(new_n121), .b(new_n108), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  aoai13aa1n02x5               g028(.a(new_n123), .b(new_n111), .c(new_n113), .d(new_n114), .o1(new_n124));
  aoi122aa1n12x5               g029(.a(new_n111), .b(\b[6] ), .c(\a[7] ), .d(\b[5] ), .e(\a[6] ), .o1(new_n125));
  oai012aa1n02x5               g030(.a(new_n123), .b(\b[6] ), .c(\a[7] ), .o1(new_n126));
  oab012aa1n02x4               g031(.a(new_n126), .b(new_n109), .c(new_n118), .out0(new_n127));
  aobi12aa1n06x5               g032(.a(new_n124), .b(new_n127), .c(new_n125), .out0(new_n128));
  nand02aa1d06x5               g033(.a(new_n122), .b(new_n128), .o1(new_n129));
  xnrc02aa1n12x5               g034(.a(\b[8] ), .b(\a[9] ), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  nor042aa1n03x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nand22aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norb02aa1n06x4               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n134), .b(new_n97), .c(new_n129), .d(new_n131), .o1(new_n135));
  aoi112aa1n02x5               g040(.a(new_n134), .b(new_n97), .c(new_n129), .d(new_n131), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(\s[10] ));
  oai012aa1n02x5               g042(.a(new_n133), .b(new_n132), .c(new_n97), .o1(new_n138));
  nor042aa1d18x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n06x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n135), .c(new_n138), .out0(\s[11] ));
  aob012aa1n03x5               g047(.a(new_n141), .b(new_n135), .c(new_n138), .out0(new_n143));
  inv000aa1d42x5               g048(.a(new_n139), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n141), .o1(new_n145));
  aoai13aa1n02x5               g050(.a(new_n144), .b(new_n145), .c(new_n135), .d(new_n138), .o1(new_n146));
  nor022aa1n08x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand22aa1n04x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nanb02aa1n02x5               g053(.a(new_n147), .b(new_n148), .out0(new_n149));
  aoib12aa1n02x5               g054(.a(new_n139), .b(new_n148), .c(new_n147), .out0(new_n150));
  aboi22aa1n03x5               g055(.a(new_n149), .b(new_n146), .c(new_n143), .d(new_n150), .out0(\s[12] ));
  oai112aa1n03x5               g056(.a(new_n125), .b(new_n115), .c(new_n118), .d(new_n109), .o1(new_n152));
  nand22aa1n02x5               g057(.a(new_n152), .b(new_n124), .o1(new_n153));
  inv040aa1n02x5               g058(.a(new_n134), .o1(new_n154));
  nona23aa1n06x5               g059(.a(new_n148), .b(new_n140), .c(new_n139), .d(new_n147), .out0(new_n155));
  nor043aa1n06x5               g060(.a(new_n155), .b(new_n154), .c(new_n130), .o1(new_n156));
  aoai13aa1n02x5               g061(.a(new_n156), .b(new_n153), .c(new_n108), .d(new_n121), .o1(new_n157));
  nano22aa1n09x5               g062(.a(new_n147), .b(new_n140), .c(new_n148), .out0(new_n158));
  oai012aa1n02x5               g063(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .o1(new_n159));
  oab012aa1n06x5               g064(.a(new_n159), .b(new_n97), .c(new_n132), .out0(new_n160));
  aoi012aa1n02x5               g065(.a(new_n147), .b(new_n139), .c(new_n148), .o1(new_n161));
  aob012aa1n02x5               g066(.a(new_n161), .b(new_n160), .c(new_n158), .out0(new_n162));
  nanb02aa1n02x5               g067(.a(new_n162), .b(new_n157), .out0(new_n163));
  nor042aa1n04x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  inv020aa1n03x5               g071(.a(new_n161), .o1(new_n167));
  aoi112aa1n02x5               g072(.a(new_n167), .b(new_n166), .c(new_n160), .d(new_n158), .o1(new_n168));
  aoi022aa1n02x5               g073(.a(new_n163), .b(new_n166), .c(new_n157), .d(new_n168), .o1(\s[13] ));
  nor042aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand02aa1n04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n164), .c(new_n163), .d(new_n165), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n164), .b(new_n172), .c(new_n163), .d(new_n166), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(\s[14] ));
  nano23aa1n06x5               g080(.a(new_n164), .b(new_n170), .c(new_n171), .d(new_n165), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n162), .c(new_n129), .d(new_n156), .o1(new_n177));
  oai012aa1d24x5               g082(.a(new_n171), .b(new_n170), .c(new_n164), .o1(new_n178));
  nor042aa1n06x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nand42aa1n03x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n177), .c(new_n178), .out0(\s[15] ));
  inv000aa1d42x5               g088(.a(new_n178), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n182), .b(new_n184), .c(new_n163), .d(new_n176), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n179), .o1(new_n186));
  aoai13aa1n02x5               g091(.a(new_n186), .b(new_n181), .c(new_n177), .d(new_n178), .o1(new_n187));
  norp02aa1n04x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  nand42aa1n03x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  nanb02aa1n02x5               g094(.a(new_n188), .b(new_n189), .out0(new_n190));
  aoib12aa1n02x5               g095(.a(new_n179), .b(new_n189), .c(new_n188), .out0(new_n191));
  aboi22aa1n03x5               g096(.a(new_n190), .b(new_n187), .c(new_n191), .d(new_n185), .out0(\s[16] ));
  nona23aa1n02x4               g097(.a(new_n171), .b(new_n165), .c(new_n164), .d(new_n170), .out0(new_n193));
  nona23aa1d18x5               g098(.a(new_n189), .b(new_n180), .c(new_n179), .d(new_n188), .out0(new_n194));
  nona22aa1n09x5               g099(.a(new_n156), .b(new_n193), .c(new_n194), .out0(new_n195));
  aoi012aa1n12x5               g100(.a(new_n195), .b(new_n122), .c(new_n128), .o1(new_n196));
  aoai13aa1n09x5               g101(.a(new_n176), .b(new_n167), .c(new_n160), .d(new_n158), .o1(new_n197));
  tech160nm_fiaoi012aa1n03p5x5 g102(.a(new_n188), .b(new_n179), .c(new_n189), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n194), .c(new_n197), .d(new_n178), .o1(new_n199));
  xorc02aa1n02x5               g104(.a(\a[17] ), .b(\b[16] ), .out0(new_n200));
  tech160nm_fioai012aa1n05x5   g105(.a(new_n200), .b(new_n199), .c(new_n196), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n194), .o1(new_n202));
  aob012aa1n06x5               g107(.a(new_n202), .b(new_n197), .c(new_n178), .out0(new_n203));
  nano23aa1n02x4               g108(.a(new_n200), .b(new_n196), .c(new_n203), .d(new_n198), .out0(new_n204));
  norb02aa1n02x5               g109(.a(new_n201), .b(new_n204), .out0(\s[17] ));
  nor042aa1n12x5               g110(.a(\b[16] ), .b(\a[17] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  nor002aa1n06x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand02aa1n03x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  norb02aa1n09x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  xnbna2aa1n03x5               g115(.a(new_n210), .b(new_n201), .c(new_n207), .out0(\s[18] ));
  and002aa1n02x5               g116(.a(new_n200), .b(new_n210), .o(new_n212));
  tech160nm_fioai012aa1n05x5   g117(.a(new_n212), .b(new_n199), .c(new_n196), .o1(new_n213));
  oaoi03aa1n02x5               g118(.a(\a[18] ), .b(\b[17] ), .c(new_n207), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  nor042aa1n12x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  nanp02aa1n04x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  norb02aa1n12x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  xnbna2aa1n03x5               g123(.a(new_n218), .b(new_n213), .c(new_n215), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fiaoi012aa1n04x5   g125(.a(new_n153), .b(new_n108), .c(new_n121), .o1(new_n221));
  oai112aa1n06x5               g126(.a(new_n203), .b(new_n198), .c(new_n195), .d(new_n221), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n218), .b(new_n214), .c(new_n222), .d(new_n212), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n216), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n218), .o1(new_n225));
  aoai13aa1n02x5               g130(.a(new_n224), .b(new_n225), .c(new_n213), .d(new_n215), .o1(new_n226));
  nor042aa1n04x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nand02aa1d06x5               g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  inv000aa1d42x5               g134(.a(\a[19] ), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\b[18] ), .o1(new_n231));
  aboi22aa1n03x5               g136(.a(new_n227), .b(new_n228), .c(new_n230), .d(new_n231), .out0(new_n232));
  aoi022aa1n03x5               g137(.a(new_n226), .b(new_n229), .c(new_n223), .d(new_n232), .o1(\s[20] ));
  nano32aa1n03x7               g138(.a(new_n225), .b(new_n200), .c(new_n229), .d(new_n210), .out0(new_n234));
  oai012aa1n02x5               g139(.a(new_n234), .b(new_n199), .c(new_n196), .o1(new_n235));
  nanb03aa1n09x5               g140(.a(new_n227), .b(new_n228), .c(new_n217), .out0(new_n236));
  oai112aa1n06x5               g141(.a(new_n224), .b(new_n209), .c(new_n208), .d(new_n206), .o1(new_n237));
  aoi012aa1n12x5               g142(.a(new_n227), .b(new_n216), .c(new_n228), .o1(new_n238));
  oai012aa1d24x5               g143(.a(new_n238), .b(new_n237), .c(new_n236), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[20] ), .b(\a[21] ), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n241), .b(new_n239), .c(new_n222), .d(new_n234), .o1(new_n242));
  nano22aa1n03x7               g147(.a(new_n227), .b(new_n217), .c(new_n228), .out0(new_n243));
  oai012aa1n02x5               g148(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .o1(new_n244));
  oab012aa1n04x5               g149(.a(new_n244), .b(new_n206), .c(new_n208), .out0(new_n245));
  inv020aa1n04x5               g150(.a(new_n238), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n241), .b(new_n246), .c(new_n245), .d(new_n243), .o1(new_n247));
  aobi12aa1n03x7               g152(.a(new_n242), .b(new_n247), .c(new_n235), .out0(\s[21] ));
  inv000aa1d42x5               g153(.a(new_n239), .o1(new_n249));
  nor042aa1n09x5               g154(.a(\b[20] ), .b(\a[21] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n02x7               g156(.a(new_n251), .b(new_n240), .c(new_n235), .d(new_n249), .o1(new_n252));
  xnrc02aa1n12x5               g157(.a(\b[21] ), .b(\a[22] ), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n253), .b(new_n250), .out0(new_n255));
  aoi022aa1n02x5               g160(.a(new_n252), .b(new_n254), .c(new_n242), .d(new_n255), .o1(\s[22] ));
  nor042aa1n06x5               g161(.a(new_n253), .b(new_n240), .o1(new_n257));
  and002aa1n02x5               g162(.a(new_n234), .b(new_n257), .o(new_n258));
  oai012aa1n02x5               g163(.a(new_n258), .b(new_n199), .c(new_n196), .o1(new_n259));
  oao003aa1n12x5               g164(.a(\a[22] ), .b(\b[21] ), .c(new_n251), .carry(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  aoi012aa1n02x5               g166(.a(new_n261), .b(new_n239), .c(new_n257), .o1(new_n262));
  inv040aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n263), .c(new_n222), .d(new_n258), .o1(new_n265));
  aoi112aa1n02x5               g170(.a(new_n264), .b(new_n261), .c(new_n239), .d(new_n257), .o1(new_n266));
  aobi12aa1n03x7               g171(.a(new_n265), .b(new_n266), .c(new_n259), .out0(\s[23] ));
  nor042aa1n06x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n264), .o1(new_n270));
  aoai13aa1n02x7               g175(.a(new_n269), .b(new_n270), .c(new_n259), .d(new_n262), .o1(new_n271));
  xorc02aa1n02x5               g176(.a(\a[24] ), .b(\b[23] ), .out0(new_n272));
  norp02aa1n02x5               g177(.a(new_n272), .b(new_n268), .o1(new_n273));
  aoi022aa1n02x5               g178(.a(new_n271), .b(new_n272), .c(new_n265), .d(new_n273), .o1(\s[24] ));
  inv020aa1n02x5               g179(.a(new_n234), .o1(new_n275));
  and002aa1n06x5               g180(.a(new_n272), .b(new_n264), .o(new_n276));
  nano22aa1n02x4               g181(.a(new_n275), .b(new_n276), .c(new_n257), .out0(new_n277));
  oai012aa1n02x5               g182(.a(new_n277), .b(new_n199), .c(new_n196), .o1(new_n278));
  aoai13aa1n09x5               g183(.a(new_n257), .b(new_n246), .c(new_n245), .d(new_n243), .o1(new_n279));
  inv030aa1n02x5               g184(.a(new_n276), .o1(new_n280));
  oao003aa1n02x5               g185(.a(\a[24] ), .b(\b[23] ), .c(new_n269), .carry(new_n281));
  aoai13aa1n12x5               g186(.a(new_n281), .b(new_n280), .c(new_n279), .d(new_n260), .o1(new_n282));
  xorc02aa1n12x5               g187(.a(\a[25] ), .b(\b[24] ), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n282), .c(new_n222), .d(new_n277), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n276), .b(new_n261), .c(new_n239), .d(new_n257), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n283), .o1(new_n286));
  and003aa1n02x5               g191(.a(new_n285), .b(new_n286), .c(new_n281), .o(new_n287));
  aobi12aa1n03x7               g192(.a(new_n284), .b(new_n287), .c(new_n278), .out0(\s[25] ));
  inv000aa1d42x5               g193(.a(new_n282), .o1(new_n289));
  nor042aa1n03x5               g194(.a(\b[24] ), .b(\a[25] ), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n286), .c(new_n278), .d(new_n289), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .out0(new_n293));
  norp02aa1n02x5               g198(.a(new_n293), .b(new_n290), .o1(new_n294));
  aoi022aa1n02x7               g199(.a(new_n292), .b(new_n293), .c(new_n284), .d(new_n294), .o1(\s[26] ));
  and002aa1n18x5               g200(.a(new_n293), .b(new_n283), .o(new_n296));
  nano32aa1n03x7               g201(.a(new_n275), .b(new_n296), .c(new_n257), .d(new_n276), .out0(new_n297));
  tech160nm_fioai012aa1n05x5   g202(.a(new_n297), .b(new_n199), .c(new_n196), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n296), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[26] ), .b(\b[25] ), .c(new_n291), .carry(new_n300));
  aoai13aa1n04x5               g205(.a(new_n300), .b(new_n299), .c(new_n285), .d(new_n281), .o1(new_n301));
  xorc02aa1n12x5               g206(.a(\a[27] ), .b(\b[26] ), .out0(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n301), .c(new_n222), .d(new_n297), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n300), .o1(new_n304));
  aoi112aa1n02x5               g209(.a(new_n302), .b(new_n304), .c(new_n282), .d(new_n296), .o1(new_n305));
  aobi12aa1n02x7               g210(.a(new_n303), .b(new_n305), .c(new_n298), .out0(\s[27] ));
  aoi012aa1n09x5               g211(.a(new_n304), .b(new_n282), .c(new_n296), .o1(new_n307));
  nor042aa1n03x5               g212(.a(\b[26] ), .b(\a[27] ), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n308), .o1(new_n309));
  inv000aa1n02x5               g214(.a(new_n302), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n309), .b(new_n310), .c(new_n307), .d(new_n298), .o1(new_n311));
  tech160nm_fixorc02aa1n02p5x5 g216(.a(\a[28] ), .b(\b[27] ), .out0(new_n312));
  norp02aa1n02x5               g217(.a(new_n312), .b(new_n308), .o1(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n303), .d(new_n313), .o1(\s[28] ));
  and002aa1n02x5               g219(.a(new_n312), .b(new_n302), .o(new_n315));
  aoai13aa1n02x5               g220(.a(new_n315), .b(new_n301), .c(new_n222), .d(new_n297), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n315), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[28] ), .b(\b[27] ), .c(new_n309), .carry(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n307), .d(new_n298), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .out0(new_n320));
  norb02aa1n02x5               g225(.a(new_n318), .b(new_n320), .out0(new_n321));
  aoi022aa1n03x5               g226(.a(new_n319), .b(new_n320), .c(new_n316), .d(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g228(.a(new_n310), .b(new_n312), .c(new_n320), .out0(new_n324));
  aoai13aa1n02x5               g229(.a(new_n324), .b(new_n301), .c(new_n222), .d(new_n297), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n324), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\b[28] ), .o1(new_n327));
  inv000aa1d42x5               g232(.a(\a[29] ), .o1(new_n328));
  oaib12aa1n02x5               g233(.a(new_n318), .b(\b[28] ), .c(new_n328), .out0(new_n329));
  oaib12aa1n02x5               g234(.a(new_n329), .b(new_n327), .c(\a[29] ), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n326), .c(new_n307), .d(new_n298), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .out0(new_n332));
  oaoi13aa1n02x5               g237(.a(new_n332), .b(new_n329), .c(new_n328), .d(new_n327), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n331), .b(new_n332), .c(new_n325), .d(new_n333), .o1(\s[30] ));
  nanb02aa1n02x5               g239(.a(\b[30] ), .b(\a[31] ), .out0(new_n335));
  nanb02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  nanp02aa1n02x5               g241(.a(new_n336), .b(new_n335), .o1(new_n337));
  nano32aa1n06x5               g242(.a(new_n310), .b(new_n332), .c(new_n312), .d(new_n320), .out0(new_n338));
  aoai13aa1n02x5               g243(.a(new_n338), .b(new_n301), .c(new_n222), .d(new_n297), .o1(new_n339));
  inv000aa1d42x5               g244(.a(new_n338), .o1(new_n340));
  norp02aa1n02x5               g245(.a(\b[29] ), .b(\a[30] ), .o1(new_n341));
  aoi022aa1n02x5               g246(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n342));
  aoi012aa1n02x5               g247(.a(new_n341), .b(new_n329), .c(new_n342), .o1(new_n343));
  aoai13aa1n03x5               g248(.a(new_n343), .b(new_n340), .c(new_n307), .d(new_n298), .o1(new_n344));
  oai112aa1n02x5               g249(.a(new_n335), .b(new_n336), .c(\b[29] ), .d(\a[30] ), .o1(new_n345));
  aoi012aa1n02x5               g250(.a(new_n345), .b(new_n329), .c(new_n342), .o1(new_n346));
  aoi022aa1n03x5               g251(.a(new_n344), .b(new_n337), .c(new_n339), .d(new_n346), .o1(\s[31] ));
  norp02aa1n02x5               g252(.a(new_n107), .b(new_n103), .o1(new_n348));
  aboi22aa1n03x5               g253(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n349));
  norp02aa1n02x5               g254(.a(new_n349), .b(new_n348), .o1(\s[3] ));
  xorc02aa1n02x5               g255(.a(\a[4] ), .b(\b[3] ), .out0(new_n351));
  norb02aa1n02x5               g256(.a(new_n104), .b(new_n351), .out0(new_n352));
  aboi22aa1n03x5               g257(.a(new_n348), .b(new_n352), .c(new_n108), .d(new_n351), .out0(\s[4] ));
  nanb02aa1n02x5               g258(.a(new_n118), .b(new_n117), .out0(new_n354));
  aoi022aa1n02x5               g259(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n355));
  norb02aa1n02x5               g260(.a(new_n355), .b(new_n118), .out0(new_n356));
  oaib12aa1n02x5               g261(.a(new_n108), .b(new_n99), .c(\b[3] ), .out0(new_n357));
  aoi022aa1n02x5               g262(.a(new_n357), .b(new_n354), .c(new_n108), .d(new_n356), .o1(\s[5] ));
  xorc02aa1n02x5               g263(.a(\a[6] ), .b(\b[5] ), .out0(new_n359));
  aoai13aa1n02x5               g264(.a(new_n359), .b(new_n118), .c(new_n108), .d(new_n355), .o1(new_n360));
  aoi112aa1n02x5               g265(.a(new_n118), .b(new_n359), .c(new_n108), .d(new_n355), .o1(new_n361));
  norb02aa1n02x5               g266(.a(new_n360), .b(new_n361), .out0(\s[6] ));
  xorc02aa1n02x5               g267(.a(\a[7] ), .b(\b[6] ), .out0(new_n363));
  xnbna2aa1n03x5               g268(.a(new_n363), .b(new_n360), .c(new_n110), .out0(\s[7] ));
  nanp02aa1n02x5               g269(.a(new_n114), .b(new_n113), .o1(new_n365));
  aob012aa1n02x5               g270(.a(new_n363), .b(new_n360), .c(new_n110), .out0(new_n366));
  norb02aa1n02x5               g271(.a(new_n123), .b(new_n111), .out0(new_n367));
  xnbna2aa1n03x5               g272(.a(new_n367), .b(new_n366), .c(new_n365), .out0(\s[8] ));
  and003aa1n02x5               g273(.a(new_n152), .b(new_n124), .c(new_n130), .o(new_n369));
  aoi022aa1n02x5               g274(.a(new_n129), .b(new_n131), .c(new_n122), .d(new_n369), .o1(\s[9] ));
endmodule


