// Benchmark "adder" written by ABC on Thu Jul 18 05:03:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n328, new_n330, new_n332, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d32x5               g001(.a(\a[3] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[2] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nanp02aa1n03x5               g005(.a(new_n99), .b(new_n100), .o1(new_n101));
  orn002aa1n02x7               g006(.a(\a[2] ), .b(\b[1] ), .o(new_n102));
  nand42aa1n04x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  aob012aa1n03x5               g008(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(new_n104));
  inv000aa1d42x5               g009(.a(\a[4] ), .o1(new_n105));
  aboi22aa1n03x5               g010(.a(\b[3] ), .b(new_n105), .c(new_n97), .d(new_n98), .out0(new_n106));
  aoai13aa1n06x5               g011(.a(new_n106), .b(new_n101), .c(new_n104), .d(new_n102), .o1(new_n107));
  xnrc02aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .out0(new_n108));
  nand02aa1n08x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  nor042aa1d18x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nanb03aa1n06x5               g016(.a(new_n110), .b(new_n111), .c(new_n109), .out0(new_n112));
  nor042aa1n02x5               g017(.a(new_n112), .b(new_n108), .o1(new_n113));
  nand42aa1n20x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nor002aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n08x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nano23aa1n03x5               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nona23aa1n02x4               g023(.a(new_n114), .b(new_n117), .c(new_n116), .d(new_n115), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\a[6] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[5] ), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(new_n120), .b(new_n121), .c(new_n110), .o1(new_n122));
  aoi012aa1n02x5               g027(.a(new_n115), .b(new_n116), .c(new_n114), .o1(new_n123));
  oai012aa1n02x5               g028(.a(new_n123), .b(new_n119), .c(new_n122), .o1(new_n124));
  aoi013aa1n02x4               g029(.a(new_n124), .b(new_n107), .c(new_n113), .d(new_n118), .o1(new_n125));
  tech160nm_fioaoi03aa1n03p5x5 g030(.a(\a[9] ), .b(\b[8] ), .c(new_n125), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand22aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor022aa1n03x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  oaoi13aa1n02x5               g037(.a(new_n132), .b(new_n129), .c(new_n126), .d(new_n128), .o1(new_n133));
  nor042aa1n03x5               g038(.a(new_n126), .b(new_n128), .o1(new_n134));
  nano22aa1n03x7               g039(.a(new_n134), .b(new_n129), .c(new_n132), .out0(new_n135));
  norp02aa1n02x5               g040(.a(new_n133), .b(new_n135), .o1(\s[11] ));
  tech160nm_fixnrc02aa1n02p5x5 g041(.a(\b[11] ), .b(\a[12] ), .out0(new_n137));
  oai012aa1n02x5               g042(.a(new_n137), .b(new_n135), .c(new_n131), .o1(new_n138));
  inv040aa1n03x5               g043(.a(new_n135), .o1(new_n139));
  nona22aa1n02x4               g044(.a(new_n139), .b(new_n137), .c(new_n131), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n140), .b(new_n138), .o1(\s[12] ));
  nanp03aa1n03x5               g046(.a(new_n107), .b(new_n113), .c(new_n118), .o1(new_n142));
  oao003aa1n02x5               g047(.a(new_n120), .b(new_n121), .c(new_n110), .carry(new_n143));
  aobi12aa1n06x5               g048(.a(new_n123), .b(new_n118), .c(new_n143), .out0(new_n144));
  nanp02aa1n02x5               g049(.a(new_n142), .b(new_n144), .o1(new_n145));
  nona23aa1n06x5               g050(.a(new_n130), .b(new_n129), .c(new_n131), .d(new_n128), .out0(new_n146));
  tech160nm_fixnrc02aa1n04x5   g051(.a(\b[8] ), .b(\a[9] ), .out0(new_n147));
  norp03aa1n02x5               g052(.a(new_n146), .b(new_n147), .c(new_n137), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n145), .b(new_n148), .o1(new_n149));
  oai022aa1n02x5               g054(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n150));
  nanp03aa1n02x5               g055(.a(new_n150), .b(new_n129), .c(new_n130), .o1(new_n151));
  oai122aa1n02x7               g056(.a(new_n151), .b(\a[12] ), .c(\b[11] ), .d(\a[11] ), .e(\b[10] ), .o1(new_n152));
  aob012aa1n02x5               g057(.a(new_n152), .b(\b[11] ), .c(\a[12] ), .out0(new_n153));
  nor022aa1n16x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  tech160nm_finand02aa1n05x5   g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n149), .c(new_n153), .out0(\s[13] ));
  inv000aa1n02x5               g062(.a(new_n148), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n153), .b(new_n158), .c(new_n142), .d(new_n144), .o1(new_n159));
  aoi012aa1n02x5               g064(.a(new_n154), .b(new_n159), .c(new_n155), .o1(new_n160));
  xnrb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand02aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nona23aa1d16x5               g068(.a(new_n163), .b(new_n155), .c(new_n154), .d(new_n162), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(new_n159), .b(new_n165), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n162), .b(new_n154), .c(new_n163), .o1(new_n167));
  nor022aa1n16x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nanp02aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nanb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n166), .c(new_n167), .out0(\s[15] ));
  nanp02aa1n02x5               g077(.a(new_n166), .b(new_n167), .o1(new_n173));
  nor002aa1n12x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1n08x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n168), .c(new_n173), .d(new_n169), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(new_n173), .b(new_n171), .o1(new_n178));
  nona22aa1n02x4               g083(.a(new_n178), .b(new_n176), .c(new_n168), .out0(new_n179));
  nanp02aa1n02x5               g084(.a(new_n179), .b(new_n177), .o1(\s[16] ));
  nor042aa1n02x5               g085(.a(new_n147), .b(new_n137), .o1(new_n181));
  nano23aa1n06x5               g086(.a(new_n168), .b(new_n174), .c(new_n175), .d(new_n169), .out0(new_n182));
  nona23aa1d24x5               g087(.a(new_n182), .b(new_n181), .c(new_n146), .d(new_n164), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  nanp02aa1n03x5               g089(.a(new_n145), .b(new_n184), .o1(new_n185));
  tech160nm_fiaoi012aa1n04x5   g090(.a(new_n174), .b(\a[15] ), .c(\b[14] ), .o1(new_n186));
  aoi012aa1n02x5               g091(.a(new_n154), .b(\a[12] ), .c(\b[11] ), .o1(new_n187));
  nona23aa1n02x4               g092(.a(new_n163), .b(new_n155), .c(new_n168), .d(new_n162), .out0(new_n188));
  nano32aa1n02x4               g093(.a(new_n188), .b(new_n187), .c(new_n186), .d(new_n175), .out0(new_n189));
  inv000aa1d42x5               g094(.a(new_n168), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n174), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n175), .o1(new_n192));
  aoai13aa1n04x5               g097(.a(new_n169), .b(new_n162), .c(new_n154), .d(new_n163), .o1(new_n193));
  aoai13aa1n03x5               g098(.a(new_n191), .b(new_n192), .c(new_n193), .d(new_n190), .o1(new_n194));
  aoi012aa1n06x5               g099(.a(new_n194), .b(new_n152), .c(new_n189), .o1(new_n195));
  aoai13aa1n12x5               g100(.a(new_n195), .b(new_n183), .c(new_n142), .d(new_n144), .o1(new_n196));
  xorc02aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  aoi112aa1n02x5               g102(.a(new_n194), .b(new_n197), .c(new_n189), .d(new_n152), .o1(new_n198));
  aoi022aa1n02x5               g103(.a(new_n196), .b(new_n197), .c(new_n185), .d(new_n198), .o1(\s[17] ));
  inv040aa1d32x5               g104(.a(\a[18] ), .o1(new_n200));
  nor002aa1d32x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  aoi012aa1n02x5               g106(.a(new_n201), .b(new_n196), .c(new_n197), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[17] ), .c(new_n200), .out0(\s[18] ));
  inv000aa1d42x5               g108(.a(\a[17] ), .o1(new_n204));
  xroi22aa1d04x5               g109(.a(new_n204), .b(\b[16] ), .c(new_n200), .d(\b[17] ), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n201), .o1(new_n206));
  oaoi03aa1n02x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n206), .o1(new_n207));
  nor002aa1n03x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nanp02aa1n04x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n196), .d(new_n205), .o1(new_n211));
  aoi112aa1n02x5               g116(.a(new_n210), .b(new_n207), .c(new_n196), .d(new_n205), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n211), .b(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  orn002aa1n02x5               g119(.a(\a[19] ), .b(\b[18] ), .o(new_n215));
  nor042aa1n03x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand02aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  xnbna2aa1n03x5               g123(.a(new_n218), .b(new_n211), .c(new_n215), .out0(\s[20] ));
  nano23aa1n03x7               g124(.a(new_n208), .b(new_n216), .c(new_n217), .d(new_n209), .out0(new_n220));
  nand02aa1n02x5               g125(.a(new_n205), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oai022aa1n02x5               g127(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n223));
  oaib12aa1n02x5               g128(.a(new_n223), .b(new_n200), .c(\b[17] ), .out0(new_n224));
  nona23aa1n02x4               g129(.a(new_n217), .b(new_n209), .c(new_n208), .d(new_n216), .out0(new_n225));
  tech160nm_fiaoi012aa1n04x5   g130(.a(new_n216), .b(new_n208), .c(new_n217), .o1(new_n226));
  tech160nm_fioai012aa1n05x5   g131(.a(new_n226), .b(new_n225), .c(new_n224), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[20] ), .b(\a[21] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n227), .c(new_n196), .d(new_n222), .o1(new_n230));
  aoi112aa1n02x5               g135(.a(new_n229), .b(new_n227), .c(new_n196), .d(new_n222), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n230), .b(new_n231), .out0(\s[21] ));
  nor042aa1n03x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[21] ), .b(\a[22] ), .out0(new_n234));
  oaib12aa1n03x5               g139(.a(new_n234), .b(new_n233), .c(new_n230), .out0(new_n235));
  nona22aa1n02x4               g140(.a(new_n230), .b(new_n234), .c(new_n233), .out0(new_n236));
  nanp02aa1n03x5               g141(.a(new_n235), .b(new_n236), .o1(\s[22] ));
  norp02aa1n24x5               g142(.a(new_n234), .b(new_n228), .o1(new_n238));
  nanp03aa1n02x5               g143(.a(new_n205), .b(new_n238), .c(new_n220), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\a[22] ), .o1(new_n240));
  inv000aa1d42x5               g145(.a(\b[21] ), .o1(new_n241));
  oaoi03aa1n09x5               g146(.a(new_n240), .b(new_n241), .c(new_n233), .o1(new_n242));
  inv030aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n243), .b(new_n227), .c(new_n238), .o1(new_n244));
  aoai13aa1n02x5               g149(.a(new_n244), .b(new_n239), .c(new_n185), .d(new_n195), .o1(new_n245));
  xorb03aa1n02x5               g150(.a(new_n245), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[23] ), .b(\b[22] ), .out0(new_n248));
  xnrc02aa1n12x5               g153(.a(\b[23] ), .b(\a[24] ), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n247), .c(new_n245), .d(new_n248), .o1(new_n250));
  oaoi13aa1n04x5               g155(.a(new_n239), .b(new_n195), .c(new_n125), .d(new_n183), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n226), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n238), .b(new_n252), .c(new_n220), .d(new_n207), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n253), .b(new_n242), .o1(new_n254));
  oai012aa1n02x5               g159(.a(new_n248), .b(new_n251), .c(new_n254), .o1(new_n255));
  nona22aa1n02x4               g160(.a(new_n255), .b(new_n249), .c(new_n247), .out0(new_n256));
  nanp02aa1n02x5               g161(.a(new_n250), .b(new_n256), .o1(\s[24] ));
  norb02aa1n02x7               g162(.a(new_n248), .b(new_n249), .out0(new_n258));
  inv000aa1n03x5               g163(.a(new_n258), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n260));
  oab012aa1n02x4               g165(.a(new_n260), .b(\a[24] ), .c(\b[23] ), .out0(new_n261));
  aoai13aa1n12x5               g166(.a(new_n261), .b(new_n259), .c(new_n253), .d(new_n242), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n238), .o1(new_n264));
  nona32aa1n06x5               g169(.a(new_n196), .b(new_n259), .c(new_n264), .d(new_n221), .out0(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n265), .c(new_n263), .out0(\s[25] ));
  nand42aa1n04x5               g172(.a(new_n265), .b(new_n263), .o1(new_n268));
  norp02aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[25] ), .b(\a[26] ), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n268), .d(new_n266), .o1(new_n271));
  nand22aa1n02x5               g176(.a(new_n268), .b(new_n266), .o1(new_n272));
  nona22aa1n02x4               g177(.a(new_n272), .b(new_n270), .c(new_n269), .out0(new_n273));
  nanp02aa1n02x5               g178(.a(new_n273), .b(new_n271), .o1(\s[26] ));
  nona23aa1d18x5               g179(.a(new_n266), .b(new_n248), .c(new_n270), .d(new_n249), .out0(new_n275));
  nona32aa1n09x5               g180(.a(new_n196), .b(new_n275), .c(new_n264), .d(new_n221), .out0(new_n276));
  norb02aa1n02x5               g181(.a(new_n266), .b(new_n270), .out0(new_n277));
  nand42aa1n06x5               g182(.a(new_n262), .b(new_n277), .o1(new_n278));
  aoi112aa1n02x5               g183(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n279));
  oab012aa1n02x4               g184(.a(new_n279), .b(\a[26] ), .c(\b[25] ), .out0(new_n280));
  nanp03aa1n06x5               g185(.a(new_n276), .b(new_n278), .c(new_n280), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  nano22aa1n02x4               g187(.a(new_n282), .b(new_n278), .c(new_n280), .out0(new_n283));
  aoi022aa1n02x5               g188(.a(new_n283), .b(new_n276), .c(new_n281), .d(new_n282), .o1(\s[27] ));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  norp02aa1n02x5               g190(.a(\b[27] ), .b(\a[28] ), .o1(new_n286));
  nand42aa1n03x5               g191(.a(\b[27] ), .b(\a[28] ), .o1(new_n287));
  nanb02aa1n06x5               g192(.a(new_n286), .b(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n285), .c(new_n281), .d(new_n282), .o1(new_n289));
  aoai13aa1n02x5               g194(.a(new_n258), .b(new_n243), .c(new_n227), .d(new_n238), .o1(new_n290));
  inv000aa1n02x5               g195(.a(new_n277), .o1(new_n291));
  aoai13aa1n02x7               g196(.a(new_n280), .b(new_n291), .c(new_n290), .d(new_n261), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n275), .o1(new_n293));
  aoai13aa1n02x5               g198(.a(new_n282), .b(new_n292), .c(new_n251), .d(new_n293), .o1(new_n294));
  nona22aa1n02x4               g199(.a(new_n294), .b(new_n288), .c(new_n285), .out0(new_n295));
  nanp02aa1n03x5               g200(.a(new_n289), .b(new_n295), .o1(\s[28] ));
  norb02aa1n02x5               g201(.a(new_n282), .b(new_n288), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n292), .c(new_n251), .d(new_n293), .o1(new_n298));
  norp02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .o1(new_n299));
  nand42aa1n03x5               g204(.a(\b[28] ), .b(\a[29] ), .o1(new_n300));
  norb02aa1n03x5               g205(.a(new_n300), .b(new_n299), .out0(new_n301));
  oai022aa1n02x5               g206(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n302));
  aboi22aa1n03x5               g207(.a(new_n299), .b(new_n300), .c(new_n302), .d(new_n287), .out0(new_n303));
  aobi12aa1n06x5               g208(.a(new_n280), .b(new_n262), .c(new_n277), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n297), .o1(new_n305));
  oai012aa1n02x5               g210(.a(new_n287), .b(new_n286), .c(new_n285), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n305), .c(new_n304), .d(new_n276), .o1(new_n307));
  aoi022aa1n03x5               g212(.a(new_n307), .b(new_n301), .c(new_n298), .d(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g214(.a(new_n288), .b(new_n282), .c(new_n301), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n292), .c(new_n251), .d(new_n293), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[30] ), .b(\b[29] ), .out0(new_n312));
  aoi113aa1n02x5               g217(.a(new_n312), .b(new_n299), .c(new_n300), .d(new_n302), .e(new_n287), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n310), .o1(new_n314));
  aoi013aa1n02x4               g219(.a(new_n299), .b(new_n302), .c(new_n300), .d(new_n287), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n314), .c(new_n304), .d(new_n276), .o1(new_n316));
  aoi022aa1n02x7               g221(.a(new_n316), .b(new_n312), .c(new_n311), .d(new_n313), .o1(\s[30] ));
  nand23aa1n03x5               g222(.a(new_n297), .b(new_n301), .c(new_n312), .o1(new_n318));
  nanb02aa1n03x5               g223(.a(new_n318), .b(new_n281), .out0(new_n319));
  xorc02aa1n02x5               g224(.a(\a[31] ), .b(\b[30] ), .out0(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(new_n322));
  aoai13aa1n02x7               g227(.a(new_n321), .b(new_n318), .c(new_n304), .d(new_n276), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n323), .b(new_n320), .c(new_n319), .d(new_n322), .o1(\s[31] ));
  xobna2aa1n03x5               g229(.a(new_n101), .b(new_n104), .c(new_n102), .out0(\s[3] ));
  nanb02aa1n02x5               g230(.a(\b[3] ), .b(new_n105), .out0(new_n326));
  aoi012aa1n02x5               g231(.a(new_n101), .b(new_n104), .c(new_n102), .o1(new_n327));
  aoi122aa1n02x5               g232(.a(new_n327), .b(new_n109), .c(new_n326), .d(new_n98), .e(new_n97), .o1(new_n328));
  aoi013aa1n02x4               g233(.a(new_n328), .b(new_n109), .c(new_n107), .d(new_n326), .o1(\s[4] ));
  norb02aa1n02x5               g234(.a(new_n111), .b(new_n110), .out0(new_n330));
  xobna2aa1n03x5               g235(.a(new_n330), .b(new_n107), .c(new_n109), .out0(\s[5] ));
  aoib12aa1n02x5               g236(.a(new_n110), .b(new_n107), .c(new_n112), .out0(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[5] ), .c(new_n120), .out0(\s[6] ));
  aob012aa1n02x5               g238(.a(new_n122), .b(new_n107), .c(new_n113), .out0(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g240(.a(new_n116), .b(new_n334), .c(new_n117), .o1(new_n336));
  xnrb03aa1n02x5               g241(.a(new_n336), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g242(.a(new_n147), .b(new_n142), .c(new_n144), .out0(\s[9] ));
endmodule


