// Benchmark "adder" written by ABC on Wed Jul 17 16:59:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n348, new_n349, new_n350, new_n351,
    new_n353, new_n354, new_n356, new_n358, new_n360, new_n361, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d24x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand02aa1d28x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  tech160nm_fioaoi03aa1n03p5x5 g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor042aa1n06x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n12x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor042aa1n12x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nanp02aa1n04x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1n09x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  aoi012aa1d24x5               g015(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  nand42aa1n16x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor042aa1d18x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand22aa1n12x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n113), .b(new_n116), .c(new_n115), .d(new_n114), .out0(new_n117));
  nor002aa1d24x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1n10x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  norb02aa1n06x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  inv000aa1d42x5               g025(.a(\b[6] ), .o1(new_n121));
  nanb02aa1d36x5               g026(.a(\a[7] ), .b(new_n121), .out0(new_n122));
  nand02aa1n04x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nano32aa1n03x7               g028(.a(new_n117), .b(new_n123), .c(new_n120), .d(new_n122), .out0(new_n124));
  inv000aa1d42x5               g029(.a(new_n118), .o1(new_n125));
  tech160nm_fioai012aa1n03p5x5 g030(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(new_n123), .b(new_n119), .o1(new_n127));
  aoai13aa1n06x5               g032(.a(new_n125), .b(new_n127), .c(new_n126), .d(new_n122), .o1(new_n128));
  nand42aa1n10x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n100), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n128), .c(new_n112), .d(new_n124), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n99), .b(new_n131), .c(new_n101), .out0(\s[10] ));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nona22aa1n02x4               g039(.a(new_n131), .b(new_n100), .c(new_n97), .out0(new_n135));
  nanp02aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  aoi022aa1n02x5               g041(.a(new_n135), .b(new_n98), .c(new_n136), .d(new_n134), .o1(new_n137));
  aoi022aa1n09x5               g042(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n138));
  aoi013aa1n02x4               g043(.a(new_n137), .b(new_n135), .c(new_n134), .d(new_n138), .o1(\s[11] ));
  nanp03aa1n02x5               g044(.a(new_n135), .b(new_n134), .c(new_n138), .o1(new_n140));
  nor002aa1n16x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1d28x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1d36x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n133), .c(new_n135), .d(new_n138), .o1(new_n144));
  norb03aa1n03x5               g049(.a(new_n142), .b(new_n133), .c(new_n141), .out0(new_n145));
  aob012aa1n02x5               g050(.a(new_n144), .b(new_n140), .c(new_n145), .out0(\s[12] ));
  nanb02aa1n12x5               g051(.a(new_n133), .b(new_n136), .out0(new_n147));
  nano23aa1d12x5               g052(.a(new_n97), .b(new_n100), .c(new_n129), .d(new_n98), .out0(new_n148));
  nona22aa1d24x5               g053(.a(new_n148), .b(new_n143), .c(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n128), .c(new_n112), .d(new_n124), .o1(new_n151));
  oai022aa1n02x5               g056(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n152));
  oaoi03aa1n02x5               g057(.a(\a[12] ), .b(\b[11] ), .c(new_n134), .o1(new_n153));
  aoi013aa1n03x5               g058(.a(new_n153), .b(new_n145), .c(new_n138), .d(new_n152), .o1(new_n154));
  nor002aa1d32x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1d28x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n151), .c(new_n154), .out0(\s[13] ));
  inv000aa1d42x5               g063(.a(new_n155), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n104), .o1(new_n160));
  tech160nm_fioaoi03aa1n03p5x5 g065(.a(\a[2] ), .b(\b[1] ), .c(new_n160), .o1(new_n161));
  nano23aa1n09x5               g066(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n162));
  aobi12aa1n06x5               g067(.a(new_n111), .b(new_n162), .c(new_n161), .out0(new_n163));
  nanb02aa1n12x5               g068(.a(new_n114), .b(new_n113), .out0(new_n164));
  nanb02aa1n12x5               g069(.a(new_n115), .b(new_n116), .out0(new_n165));
  inv040aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  nand02aa1d04x5               g071(.a(new_n122), .b(new_n123), .o1(new_n167));
  nona23aa1n02x5               g072(.a(new_n166), .b(new_n120), .c(new_n164), .d(new_n167), .out0(new_n168));
  oabi12aa1n06x5               g073(.a(new_n128), .b(new_n163), .c(new_n168), .out0(new_n169));
  nanp03aa1n03x5               g074(.a(new_n145), .b(new_n152), .c(new_n138), .o1(new_n170));
  oaib12aa1n06x5               g075(.a(new_n170), .b(new_n145), .c(new_n142), .out0(new_n171));
  aoai13aa1n02x5               g076(.a(new_n157), .b(new_n171), .c(new_n169), .d(new_n150), .o1(new_n172));
  nor002aa1d32x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nand42aa1d28x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  nona23aa1n02x4               g080(.a(new_n172), .b(new_n174), .c(new_n173), .d(new_n155), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n175), .c(new_n159), .d(new_n172), .o1(\s[14] ));
  nano23aa1d15x5               g082(.a(new_n155), .b(new_n173), .c(new_n174), .d(new_n156), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n171), .c(new_n169), .d(new_n150), .o1(new_n179));
  tech160nm_fioai012aa1n03p5x5 g084(.a(new_n174), .b(new_n173), .c(new_n155), .o1(new_n180));
  tech160nm_fixorc02aa1n05x5   g085(.a(\a[15] ), .b(\b[14] ), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n179), .c(new_n180), .out0(\s[15] ));
  aobi12aa1n02x5               g087(.a(new_n181), .b(new_n179), .c(new_n180), .out0(new_n183));
  inv000aa1d42x5               g088(.a(\a[15] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\b[14] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n178), .o1(new_n186));
  aoai13aa1n02x5               g091(.a(new_n180), .b(new_n186), .c(new_n151), .d(new_n154), .o1(new_n187));
  oaoi03aa1n02x5               g092(.a(new_n184), .b(new_n185), .c(new_n187), .o1(new_n188));
  tech160nm_fixorc02aa1n04x5   g093(.a(\a[16] ), .b(\b[15] ), .out0(new_n189));
  nanp02aa1n02x5               g094(.a(new_n185), .b(new_n184), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n189), .b(new_n190), .o1(new_n191));
  oai022aa1n02x5               g096(.a(new_n188), .b(new_n189), .c(new_n183), .d(new_n191), .o1(\s[16] ));
  nand23aa1n09x5               g097(.a(new_n178), .b(new_n181), .c(new_n189), .o1(new_n193));
  nor042aa1n09x5               g098(.a(new_n193), .b(new_n149), .o1(new_n194));
  aoai13aa1n12x5               g099(.a(new_n194), .b(new_n128), .c(new_n112), .d(new_n124), .o1(new_n195));
  inv000aa1d42x5               g100(.a(\a[16] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[15] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  oai022aa1n02x5               g103(.a(new_n184), .b(new_n185), .c(new_n197), .d(new_n196), .o1(new_n199));
  aoai13aa1n06x5               g104(.a(new_n198), .b(new_n199), .c(new_n180), .d(new_n190), .o1(new_n200));
  aoib12aa1n12x5               g105(.a(new_n200), .b(new_n171), .c(new_n193), .out0(new_n201));
  nor042aa1n04x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  nand42aa1d28x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n195), .c(new_n201), .out0(\s[17] ));
  nand42aa1n06x5               g110(.a(new_n195), .b(new_n201), .o1(new_n206));
  aoi012aa1n02x5               g111(.a(new_n202), .b(new_n206), .c(new_n203), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand42aa1d28x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  oaih22aa1d12x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  aoi122aa1n06x5               g116(.a(new_n211), .b(\b[17] ), .c(\a[18] ), .d(new_n206), .e(new_n204), .o1(new_n212));
  oabi12aa1n03x5               g117(.a(new_n212), .b(new_n207), .c(new_n210), .out0(\s[18] ));
  oabi12aa1n06x5               g118(.a(new_n200), .b(new_n154), .c(new_n193), .out0(new_n214));
  nano23aa1d15x5               g119(.a(new_n202), .b(new_n208), .c(new_n209), .d(new_n203), .out0(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n214), .c(new_n169), .d(new_n194), .o1(new_n216));
  oai012aa1n02x5               g121(.a(new_n209), .b(new_n208), .c(new_n202), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[19] ), .b(\b[18] ), .out0(new_n218));
  xnbna2aa1n03x5               g123(.a(new_n218), .b(new_n216), .c(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aobi12aa1n02x7               g125(.a(new_n218), .b(new_n216), .c(new_n217), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n215), .o1(new_n222));
  aoai13aa1n02x7               g127(.a(new_n217), .b(new_n222), .c(new_n195), .d(new_n201), .o1(new_n223));
  inv040aa1d32x5               g128(.a(\a[19] ), .o1(new_n224));
  inv040aa1d32x5               g129(.a(\b[18] ), .o1(new_n225));
  nand02aa1n12x5               g130(.a(new_n225), .b(new_n224), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  tech160nm_finand02aa1n03p5x5 g132(.a(\b[18] ), .b(\a[19] ), .o1(new_n228));
  norp02aa1n24x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  nand42aa1d28x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(new_n229), .b(new_n230), .out0(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n227), .c(new_n223), .d(new_n228), .o1(new_n232));
  nano22aa1n02x4               g137(.a(new_n229), .b(new_n226), .c(new_n230), .out0(new_n233));
  oaib12aa1n03x5               g138(.a(new_n232), .b(new_n221), .c(new_n233), .out0(\s[20] ));
  nano22aa1n03x7               g139(.a(new_n231), .b(new_n226), .c(new_n228), .out0(new_n235));
  nand22aa1n12x5               g140(.a(new_n235), .b(new_n215), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n214), .c(new_n169), .d(new_n194), .o1(new_n238));
  nanb03aa1n06x5               g143(.a(new_n229), .b(new_n230), .c(new_n228), .out0(new_n239));
  nand23aa1n04x5               g144(.a(new_n211), .b(new_n226), .c(new_n209), .o1(new_n240));
  aoai13aa1n12x5               g145(.a(new_n230), .b(new_n229), .c(new_n224), .d(new_n225), .o1(new_n241));
  oai012aa1n18x5               g146(.a(new_n241), .b(new_n240), .c(new_n239), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  nor022aa1n08x5               g148(.a(\b[20] ), .b(\a[21] ), .o1(new_n244));
  nand42aa1n16x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  xnbna2aa1n03x5               g151(.a(new_n246), .b(new_n238), .c(new_n243), .out0(\s[21] ));
  aobi12aa1n02x5               g152(.a(new_n246), .b(new_n238), .c(new_n243), .out0(new_n248));
  aoai13aa1n03x5               g153(.a(new_n243), .b(new_n236), .c(new_n195), .d(new_n201), .o1(new_n249));
  aoi012aa1n03x5               g154(.a(new_n244), .b(new_n249), .c(new_n245), .o1(new_n250));
  nor042aa1n04x5               g155(.a(\b[21] ), .b(\a[22] ), .o1(new_n251));
  nand42aa1n08x5               g156(.a(\b[21] ), .b(\a[22] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  nona22aa1n02x4               g158(.a(new_n252), .b(new_n251), .c(new_n244), .out0(new_n254));
  oai022aa1n03x5               g159(.a(new_n250), .b(new_n253), .c(new_n254), .d(new_n248), .o1(\s[22] ));
  nano23aa1d15x5               g160(.a(new_n244), .b(new_n251), .c(new_n252), .d(new_n245), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  nona22aa1n02x4               g162(.a(new_n206), .b(new_n236), .c(new_n257), .out0(new_n258));
  nanp03aa1n02x5               g163(.a(new_n235), .b(new_n215), .c(new_n256), .o1(new_n259));
  nano22aa1n02x4               g164(.a(new_n229), .b(new_n228), .c(new_n230), .out0(new_n260));
  oai012aa1n02x5               g165(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .o1(new_n261));
  oab012aa1n03x5               g166(.a(new_n261), .b(new_n202), .c(new_n208), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n241), .o1(new_n263));
  aoai13aa1n06x5               g168(.a(new_n256), .b(new_n263), .c(new_n262), .d(new_n260), .o1(new_n264));
  oa0012aa1n02x5               g169(.a(new_n252), .b(new_n251), .c(new_n244), .o(new_n265));
  inv020aa1n03x5               g170(.a(new_n265), .o1(new_n266));
  nanp02aa1n02x5               g171(.a(new_n264), .b(new_n266), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n04x5               g173(.a(new_n268), .b(new_n259), .c(new_n195), .d(new_n201), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[23] ), .b(\b[22] ), .out0(new_n270));
  aoi112aa1n02x5               g175(.a(new_n270), .b(new_n265), .c(new_n242), .d(new_n256), .o1(new_n271));
  aoi022aa1n02x5               g176(.a(new_n271), .b(new_n258), .c(new_n269), .d(new_n270), .o1(\s[23] ));
  norp02aa1n02x5               g177(.a(\b[22] ), .b(\a[23] ), .o1(new_n273));
  tech160nm_fixnrc02aa1n04x5   g178(.a(\b[23] ), .b(\a[24] ), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n269), .d(new_n270), .o1(new_n275));
  norp02aa1n02x5               g180(.a(new_n274), .b(new_n273), .o1(new_n276));
  aob012aa1n03x5               g181(.a(new_n276), .b(new_n269), .c(new_n270), .out0(new_n277));
  nanp02aa1n03x5               g182(.a(new_n275), .b(new_n277), .o1(\s[24] ));
  norb02aa1n12x5               g183(.a(new_n270), .b(new_n274), .out0(new_n279));
  nona23aa1n02x4               g184(.a(new_n279), .b(new_n235), .c(new_n222), .d(new_n257), .out0(new_n280));
  inv000aa1d42x5               g185(.a(new_n279), .o1(new_n281));
  orn002aa1n02x5               g186(.a(\a[23] ), .b(\b[22] ), .o(new_n282));
  oao003aa1n02x5               g187(.a(\a[24] ), .b(\b[23] ), .c(new_n282), .carry(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n281), .c(new_n264), .d(new_n266), .o1(new_n284));
  inv040aa1n02x5               g189(.a(new_n284), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n285), .b(new_n280), .c(new_n195), .d(new_n201), .o1(new_n286));
  xorb03aa1n02x5               g191(.a(new_n286), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  xnrc02aa1n12x5               g193(.a(\b[24] ), .b(\a[25] ), .out0(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  tech160nm_fixnrc02aa1n05x5   g195(.a(\b[25] ), .b(\a[26] ), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n288), .c(new_n286), .d(new_n290), .o1(new_n292));
  norp02aa1n02x5               g197(.a(new_n291), .b(new_n288), .o1(new_n293));
  aob012aa1n03x5               g198(.a(new_n293), .b(new_n286), .c(new_n290), .out0(new_n294));
  nanp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[26] ));
  nor002aa1n03x5               g200(.a(new_n291), .b(new_n289), .o1(new_n296));
  inv000aa1n03x5               g201(.a(new_n296), .o1(new_n297));
  nano23aa1d12x5               g202(.a(new_n236), .b(new_n297), .c(new_n279), .d(new_n256), .out0(new_n298));
  aoai13aa1n06x5               g203(.a(new_n298), .b(new_n214), .c(new_n169), .d(new_n194), .o1(new_n299));
  nanp02aa1n02x5               g204(.a(\b[25] ), .b(\a[26] ), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n293), .o1(new_n301));
  aoi022aa1n12x5               g206(.a(new_n284), .b(new_n296), .c(new_n300), .d(new_n301), .o1(new_n302));
  xorc02aa1n12x5               g207(.a(\a[27] ), .b(\b[26] ), .out0(new_n303));
  xnbna2aa1n03x5               g208(.a(new_n303), .b(new_n302), .c(new_n299), .out0(\s[27] ));
  norp02aa1n02x5               g209(.a(\b[26] ), .b(\a[27] ), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n305), .o1(new_n306));
  aoai13aa1n04x5               g211(.a(new_n279), .b(new_n265), .c(new_n242), .d(new_n256), .o1(new_n307));
  oai012aa1n02x5               g212(.a(new_n300), .b(new_n291), .c(new_n288), .o1(new_n308));
  aoai13aa1n04x5               g213(.a(new_n308), .b(new_n297), .c(new_n307), .d(new_n283), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n303), .b(new_n309), .c(new_n206), .d(new_n298), .o1(new_n310));
  tech160nm_fixorc02aa1n02p5x5 g215(.a(\a[28] ), .b(\b[27] ), .out0(new_n311));
  inv000aa1d42x5               g216(.a(new_n303), .o1(new_n312));
  oai022aa1d18x5               g217(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n313));
  aoi012aa1n02x5               g218(.a(new_n313), .b(\a[28] ), .c(\b[27] ), .o1(new_n314));
  aoai13aa1n04x5               g219(.a(new_n314), .b(new_n312), .c(new_n302), .d(new_n299), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n310), .d(new_n306), .o1(\s[28] ));
  and002aa1n02x5               g221(.a(new_n311), .b(new_n303), .o(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n309), .c(new_n206), .d(new_n298), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  aob012aa1n12x5               g224(.a(new_n313), .b(\b[27] ), .c(\a[28] ), .out0(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n319), .c(new_n302), .d(new_n299), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n320), .b(new_n322), .out0(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g230(.a(new_n312), .b(new_n311), .c(new_n322), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n309), .c(new_n206), .d(new_n298), .o1(new_n327));
  inv000aa1d42x5               g232(.a(new_n326), .o1(new_n328));
  tech160nm_fioaoi03aa1n03p5x5 g233(.a(\a[29] ), .b(\b[28] ), .c(new_n320), .o1(new_n329));
  inv000aa1d42x5               g234(.a(new_n329), .o1(new_n330));
  aoai13aa1n06x5               g235(.a(new_n330), .b(new_n328), .c(new_n302), .d(new_n299), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .out0(new_n332));
  norp02aa1n02x5               g237(.a(\b[28] ), .b(\a[29] ), .o1(new_n333));
  aoi012aa1n02x5               g238(.a(new_n320), .b(\a[29] ), .c(\b[28] ), .o1(new_n334));
  norp03aa1n02x5               g239(.a(new_n334), .b(new_n332), .c(new_n333), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n331), .b(new_n332), .c(new_n327), .d(new_n335), .o1(\s[30] ));
  nano32aa1n06x5               g241(.a(new_n312), .b(new_n332), .c(new_n311), .d(new_n322), .out0(new_n337));
  aoai13aa1n03x5               g242(.a(new_n337), .b(new_n309), .c(new_n206), .d(new_n298), .o1(new_n338));
  xorc02aa1n02x5               g243(.a(\a[31] ), .b(\b[30] ), .out0(new_n339));
  inv000aa1d42x5               g244(.a(\a[30] ), .o1(new_n340));
  inv000aa1d42x5               g245(.a(\b[29] ), .o1(new_n341));
  oabi12aa1n02x5               g246(.a(new_n339), .b(\a[30] ), .c(\b[29] ), .out0(new_n342));
  oaoi13aa1n02x5               g247(.a(new_n342), .b(new_n329), .c(new_n340), .d(new_n341), .o1(new_n343));
  inv000aa1d42x5               g248(.a(new_n337), .o1(new_n344));
  oaoi03aa1n02x5               g249(.a(new_n340), .b(new_n341), .c(new_n329), .o1(new_n345));
  aoai13aa1n04x5               g250(.a(new_n345), .b(new_n344), .c(new_n302), .d(new_n299), .o1(new_n346));
  aoi022aa1n03x5               g251(.a(new_n346), .b(new_n339), .c(new_n338), .d(new_n343), .o1(\s[31] ));
  aoi022aa1n02x5               g252(.a(new_n103), .b(new_n102), .c(\a[1] ), .d(\b[0] ), .o1(new_n348));
  oaib12aa1n02x5               g253(.a(new_n348), .b(new_n103), .c(\a[2] ), .out0(new_n349));
  norb02aa1n02x5               g254(.a(new_n109), .b(new_n108), .out0(new_n350));
  aboi22aa1n03x5               g255(.a(new_n108), .b(new_n109), .c(new_n102), .d(new_n103), .out0(new_n351));
  aoi022aa1n02x5               g256(.a(new_n349), .b(new_n351), .c(new_n161), .d(new_n350), .o1(\s[3] ));
  obai22aa1n02x7               g257(.a(new_n107), .b(new_n106), .c(\a[3] ), .d(\b[2] ), .out0(new_n353));
  aoi012aa1n02x5               g258(.a(new_n353), .b(new_n161), .c(new_n350), .o1(new_n354));
  oaoi13aa1n02x5               g259(.a(new_n354), .b(new_n112), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  oai112aa1n02x5               g260(.a(new_n111), .b(new_n165), .c(new_n110), .d(new_n105), .o1(new_n356));
  aobi12aa1n02x5               g261(.a(new_n356), .b(new_n166), .c(new_n112), .out0(\s[5] ));
  oaoi03aa1n02x5               g262(.a(\a[5] ), .b(\b[4] ), .c(new_n163), .o1(new_n358));
  xorb03aa1n02x5               g263(.a(new_n358), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g264(.a(new_n167), .b(new_n114), .c(new_n358), .d(new_n113), .o1(new_n360));
  nanb02aa1n02x5               g265(.a(new_n164), .b(new_n358), .out0(new_n361));
  nona22aa1n02x4               g266(.a(new_n361), .b(new_n167), .c(new_n114), .out0(new_n362));
  nanp02aa1n02x5               g267(.a(new_n362), .b(new_n360), .o1(\s[7] ));
  xobna2aa1n03x5               g268(.a(new_n120), .b(new_n362), .c(new_n123), .out0(\s[8] ));
  xorb03aa1n02x5               g269(.a(new_n169), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


