// Benchmark "adder" written by ABC on Thu Jul 18 10:50:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n180, new_n181,
    new_n182, new_n183, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n323, new_n326,
    new_n328, new_n329, new_n330;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  aoi012aa1n09x5               g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  norp02aa1n09x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nand22aa1n12x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n02x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  ao0012aa1n03x5               g010(.a(new_n101), .b(new_n103), .c(new_n102), .o(new_n106));
  oabi12aa1n06x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .out0(new_n107));
  nand02aa1d28x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor002aa1n20x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand02aa1d24x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb03aa1n06x5               g015(.a(new_n109), .b(new_n110), .c(new_n108), .out0(new_n111));
  xnrc02aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .out0(new_n112));
  nor042aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor042aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nona22aa1n02x4               g020(.a(new_n115), .b(new_n114), .c(new_n113), .out0(new_n116));
  nor043aa1n03x5               g021(.a(new_n116), .b(new_n111), .c(new_n112), .o1(new_n117));
  oai022aa1d18x5               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  aoi013aa1n03x5               g023(.a(new_n109), .b(new_n118), .c(new_n110), .d(new_n108), .o1(new_n119));
  oaoi03aa1n09x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  tech160nm_fiaoi012aa1n05x5   g025(.a(new_n120), .b(new_n107), .c(new_n117), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .c(new_n121), .o1(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nor002aa1n06x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand22aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nano23aa1n06x5               g032(.a(new_n124), .b(new_n126), .c(new_n127), .d(new_n125), .out0(new_n128));
  inv040aa1n03x5               g033(.a(new_n128), .o1(new_n129));
  oai012aa1n06x5               g034(.a(new_n127), .b(new_n126), .c(new_n124), .o1(new_n130));
  oai012aa1n03x5               g035(.a(new_n130), .b(new_n121), .c(new_n129), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g037(.a(\a[12] ), .o1(new_n133));
  norp02aa1n06x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanp02aa1n06x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  aoi012aa1n03x5               g040(.a(new_n134), .b(new_n131), .c(new_n135), .o1(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[11] ), .c(new_n133), .out0(\s[12] ));
  norb02aa1n02x5               g042(.a(new_n135), .b(new_n134), .out0(new_n138));
  xorc02aa1n02x5               g043(.a(\a[12] ), .b(\b[11] ), .out0(new_n139));
  nano22aa1n03x7               g044(.a(new_n129), .b(new_n139), .c(new_n138), .out0(new_n140));
  aoai13aa1n03x5               g045(.a(new_n140), .b(new_n120), .c(new_n107), .d(new_n117), .o1(new_n141));
  inv000aa1d42x5               g046(.a(\b[11] ), .o1(new_n142));
  tech160nm_fiaoi012aa1n04x5   g047(.a(new_n134), .b(new_n133), .c(new_n142), .o1(new_n143));
  nand42aa1n02x5               g048(.a(new_n130), .b(new_n143), .o1(new_n144));
  aoai13aa1n04x5               g049(.a(\a[12] ), .b(\b[11] ), .c(\b[10] ), .d(\a[11] ), .o1(new_n145));
  oaib12aa1n06x5               g050(.a(new_n145), .b(new_n135), .c(\b[11] ), .out0(new_n146));
  oaib12aa1n02x5               g051(.a(new_n141), .b(new_n146), .c(new_n144), .out0(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n16x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nanp02aa1n04x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  aoi012aa1n02x5               g055(.a(new_n149), .b(new_n147), .c(new_n150), .o1(new_n151));
  xnrb03aa1n03x5               g056(.a(new_n151), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nand22aa1n09x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nona23aa1d18x5               g059(.a(new_n154), .b(new_n150), .c(new_n149), .d(new_n153), .out0(new_n155));
  oao003aa1n02x5               g060(.a(new_n133), .b(new_n142), .c(new_n135), .carry(new_n156));
  nano23aa1n06x5               g061(.a(new_n149), .b(new_n153), .c(new_n154), .d(new_n150), .out0(new_n157));
  nanp03aa1n02x5               g062(.a(new_n144), .b(new_n157), .c(new_n156), .o1(new_n158));
  tech160nm_fiaoi012aa1n03p5x5 g063(.a(new_n153), .b(new_n149), .c(new_n154), .o1(new_n159));
  oai112aa1n03x5               g064(.a(new_n158), .b(new_n159), .c(new_n141), .d(new_n155), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  xnrc02aa1n12x5               g067(.a(\b[14] ), .b(\a[15] ), .out0(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  xnrc02aa1n12x5               g069(.a(\b[15] ), .b(\a[16] ), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n162), .c(new_n160), .d(new_n164), .o1(new_n166));
  aoi112aa1n03x4               g071(.a(new_n162), .b(new_n165), .c(new_n160), .d(new_n164), .o1(new_n167));
  nanb02aa1n03x5               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  nona32aa1n02x4               g073(.a(new_n140), .b(new_n165), .c(new_n163), .d(new_n155), .out0(new_n169));
  aoi112aa1n03x5               g074(.a(new_n155), .b(new_n146), .c(new_n130), .d(new_n143), .o1(new_n170));
  inv000aa1n02x5               g075(.a(new_n159), .o1(new_n171));
  norp02aa1n24x5               g076(.a(new_n165), .b(new_n163), .o1(new_n172));
  inv000aa1d42x5               g077(.a(\a[16] ), .o1(new_n173));
  inv000aa1d42x5               g078(.a(\b[15] ), .o1(new_n174));
  tech160nm_fioaoi03aa1n02p5x5 g079(.a(new_n173), .b(new_n174), .c(new_n162), .o1(new_n175));
  inv000aa1n02x5               g080(.a(new_n175), .o1(new_n176));
  oaoi13aa1n12x5               g081(.a(new_n176), .b(new_n172), .c(new_n170), .d(new_n171), .o1(new_n177));
  oai012aa1n06x5               g082(.a(new_n177), .b(new_n121), .c(new_n169), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g084(.a(\a[18] ), .o1(new_n180));
  inv040aa1d30x5               g085(.a(\a[17] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\b[16] ), .o1(new_n182));
  oaoi03aa1n03x5               g087(.a(new_n181), .b(new_n182), .c(new_n178), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[17] ), .c(new_n180), .out0(\s[18] ));
  nanp03aa1n02x5               g089(.a(new_n128), .b(new_n138), .c(new_n139), .o1(new_n185));
  nano22aa1n03x7               g090(.a(new_n185), .b(new_n172), .c(new_n157), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n120), .c(new_n107), .d(new_n117), .o1(new_n187));
  xroi22aa1d06x4               g092(.a(new_n181), .b(\b[16] ), .c(new_n180), .d(\b[17] ), .out0(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\b[17] ), .o1(new_n190));
  oai022aa1d24x5               g095(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n191));
  oaib12aa1n18x5               g096(.a(new_n191), .b(new_n190), .c(\a[18] ), .out0(new_n192));
  aoai13aa1n04x5               g097(.a(new_n192), .b(new_n189), .c(new_n187), .d(new_n177), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n08x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nand02aa1n03x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  xnrc02aa1n02x5               g102(.a(\b[19] ), .b(\a[20] ), .out0(new_n198));
  aoai13aa1n03x5               g103(.a(new_n198), .b(new_n196), .c(new_n193), .d(new_n197), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n196), .b(new_n197), .out0(new_n200));
  nanb02aa1n03x5               g105(.a(new_n200), .b(new_n193), .out0(new_n201));
  nona22aa1n02x5               g106(.a(new_n201), .b(new_n198), .c(new_n196), .out0(new_n202));
  nand42aa1n02x5               g107(.a(new_n202), .b(new_n199), .o1(\s[20] ));
  nona22aa1n03x5               g108(.a(new_n188), .b(new_n200), .c(new_n198), .out0(new_n204));
  inv000aa1d42x5               g109(.a(\a[20] ), .o1(new_n205));
  inv000aa1d42x5               g110(.a(\b[19] ), .o1(new_n206));
  aoi012aa1n06x5               g111(.a(new_n196), .b(new_n205), .c(new_n206), .o1(new_n207));
  aoai13aa1n12x5               g112(.a(\a[20] ), .b(\b[19] ), .c(\b[18] ), .d(\a[19] ), .o1(new_n208));
  oaib12aa1n06x5               g113(.a(new_n208), .b(new_n197), .c(\b[19] ), .out0(new_n209));
  aoi012aa1n12x5               g114(.a(new_n209), .b(new_n192), .c(new_n207), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n204), .c(new_n187), .d(new_n177), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g118(.a(\b[20] ), .b(\a[21] ), .o1(new_n214));
  nand22aa1n03x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  nor042aa1n06x5               g121(.a(\b[21] ), .b(\a[22] ), .o1(new_n217));
  nand02aa1d08x5               g122(.a(\b[21] ), .b(\a[22] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n214), .c(new_n212), .d(new_n216), .o1(new_n220));
  inv040aa1n03x5               g125(.a(new_n204), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n216), .b(new_n210), .c(new_n178), .d(new_n221), .o1(new_n222));
  nona22aa1n03x5               g127(.a(new_n222), .b(new_n219), .c(new_n214), .out0(new_n223));
  nanp02aa1n03x5               g128(.a(new_n220), .b(new_n223), .o1(\s[22] ));
  nona23aa1n02x4               g129(.a(new_n218), .b(new_n215), .c(new_n214), .d(new_n217), .out0(new_n225));
  nona32aa1n03x5               g130(.a(new_n188), .b(new_n225), .c(new_n198), .d(new_n200), .out0(new_n226));
  nand42aa1n02x5               g131(.a(new_n192), .b(new_n207), .o1(new_n227));
  oao003aa1n03x5               g132(.a(new_n205), .b(new_n206), .c(new_n197), .carry(new_n228));
  nano23aa1n06x5               g133(.a(new_n214), .b(new_n217), .c(new_n218), .d(new_n215), .out0(new_n229));
  aoi012aa1d18x5               g134(.a(new_n217), .b(new_n214), .c(new_n218), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoi013aa1n02x4               g136(.a(new_n231), .b(new_n227), .c(new_n229), .d(new_n228), .o1(new_n232));
  aoai13aa1n04x5               g137(.a(new_n232), .b(new_n226), .c(new_n187), .d(new_n177), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  xorc02aa1n12x5               g140(.a(\a[23] ), .b(\b[22] ), .out0(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[23] ), .b(\a[24] ), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n235), .c(new_n233), .d(new_n236), .o1(new_n238));
  nand02aa1n02x5               g143(.a(new_n233), .b(new_n236), .o1(new_n239));
  nona22aa1n02x5               g144(.a(new_n239), .b(new_n237), .c(new_n235), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[24] ));
  norb02aa1n03x5               g146(.a(new_n236), .b(new_n237), .out0(new_n242));
  inv040aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  nona22aa1n03x5               g148(.a(new_n221), .b(new_n243), .c(new_n225), .out0(new_n244));
  nand23aa1n03x5               g149(.a(new_n227), .b(new_n229), .c(new_n228), .o1(new_n245));
  orn002aa1n02x5               g150(.a(\a[23] ), .b(\b[22] ), .o(new_n246));
  oao003aa1n02x5               g151(.a(\a[24] ), .b(\b[23] ), .c(new_n246), .carry(new_n247));
  aoai13aa1n12x5               g152(.a(new_n247), .b(new_n243), .c(new_n245), .d(new_n230), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n244), .c(new_n187), .d(new_n177), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  tech160nm_fixorc02aa1n05x5   g157(.a(\a[25] ), .b(\b[24] ), .out0(new_n253));
  xnrc02aa1n12x5               g158(.a(\b[25] ), .b(\a[26] ), .out0(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n252), .c(new_n250), .d(new_n253), .o1(new_n255));
  nand02aa1n02x5               g160(.a(new_n250), .b(new_n253), .o1(new_n256));
  nona22aa1n02x5               g161(.a(new_n256), .b(new_n254), .c(new_n252), .out0(new_n257));
  nanp02aa1n03x5               g162(.a(new_n257), .b(new_n255), .o1(\s[26] ));
  inv000aa1n03x5               g163(.a(new_n100), .o1(new_n259));
  nano23aa1n02x4               g164(.a(new_n101), .b(new_n103), .c(new_n104), .d(new_n102), .out0(new_n260));
  aoi012aa1n02x5               g165(.a(new_n106), .b(new_n260), .c(new_n259), .o1(new_n261));
  inv000aa1d42x5               g166(.a(\a[8] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(\b[7] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n108), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n109), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n110), .o1(new_n266));
  norp02aa1n02x5               g171(.a(new_n114), .b(new_n113), .o1(new_n267));
  oai013aa1n02x4               g172(.a(new_n265), .b(new_n267), .c(new_n266), .d(new_n264), .o1(new_n268));
  oaoi03aa1n02x5               g173(.a(new_n262), .b(new_n263), .c(new_n268), .o1(new_n269));
  oaib12aa1n03x5               g174(.a(new_n269), .b(new_n261), .c(new_n117), .out0(new_n270));
  inv000aa1n02x5               g175(.a(new_n172), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n175), .b(new_n271), .c(new_n158), .d(new_n159), .o1(new_n272));
  norb02aa1n06x5               g177(.a(new_n253), .b(new_n254), .out0(new_n273));
  nano22aa1n03x7               g178(.a(new_n226), .b(new_n242), .c(new_n273), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .d(new_n186), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n276));
  oab012aa1n02x4               g181(.a(new_n276), .b(\a[26] ), .c(\b[25] ), .out0(new_n277));
  aobi12aa1n12x5               g182(.a(new_n277), .b(new_n248), .c(new_n273), .out0(new_n278));
  tech160nm_fixorc02aa1n02p5x5 g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  xnbna2aa1n03x5               g184(.a(new_n279), .b(new_n275), .c(new_n278), .out0(\s[27] ));
  nand42aa1n03x5               g185(.a(new_n275), .b(new_n278), .o1(new_n281));
  norp02aa1n02x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  norp02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .o1(new_n283));
  nand42aa1n03x5               g188(.a(\b[27] ), .b(\a[28] ), .o1(new_n284));
  norb02aa1n06x4               g189(.a(new_n284), .b(new_n283), .out0(new_n285));
  inv040aa1n03x5               g190(.a(new_n285), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n282), .c(new_n281), .d(new_n279), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n242), .b(new_n231), .c(new_n210), .d(new_n229), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n273), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n277), .b(new_n289), .c(new_n288), .d(new_n247), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n279), .b(new_n290), .c(new_n178), .d(new_n274), .o1(new_n291));
  nona22aa1n02x5               g196(.a(new_n291), .b(new_n286), .c(new_n282), .out0(new_n292));
  nanp02aa1n03x5               g197(.a(new_n287), .b(new_n292), .o1(\s[28] ));
  norb02aa1n02x5               g198(.a(new_n279), .b(new_n286), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n290), .c(new_n178), .d(new_n274), .o1(new_n295));
  aoi012aa1n02x5               g200(.a(new_n283), .b(new_n282), .c(new_n284), .o1(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[28] ), .b(\a[29] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n295), .c(new_n296), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n294), .o1(new_n299));
  tech160nm_fiaoi012aa1n02p5x5 g204(.a(new_n299), .b(new_n275), .c(new_n278), .o1(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n297), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n298), .b(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n09x5               g208(.a(new_n297), .b(new_n279), .c(new_n285), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n290), .c(new_n178), .d(new_n274), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[29] ), .b(\a[30] ), .out0(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n307), .b(new_n305), .c(new_n306), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n304), .o1(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n309), .b(new_n275), .c(new_n278), .o1(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n307), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n308), .b(new_n311), .o1(\s[30] ));
  nano23aa1n06x5               g217(.a(new_n307), .b(new_n297), .c(new_n279), .d(new_n285), .out0(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n290), .c(new_n178), .d(new_n274), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n314), .c(new_n315), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n313), .o1(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n318), .b(new_n275), .c(new_n278), .o1(new_n319));
  nano22aa1n02x4               g224(.a(new_n319), .b(new_n315), .c(new_n316), .out0(new_n320));
  norp02aa1n03x5               g225(.a(new_n317), .b(new_n320), .o1(\s[31] ));
  xnrb03aa1n02x5               g226(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g227(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g229(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g230(.a(\a[5] ), .b(\b[4] ), .c(new_n261), .o1(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb03aa1n02x5               g232(.a(new_n115), .b(new_n261), .c(new_n114), .out0(new_n328));
  oabi12aa1n02x5               g233(.a(new_n111), .b(new_n328), .c(new_n118), .out0(new_n329));
  aoi122aa1n02x5               g234(.a(new_n113), .b(new_n265), .c(new_n110), .d(new_n326), .e(new_n108), .o1(new_n330));
  norb02aa1n02x5               g235(.a(new_n329), .b(new_n330), .out0(\s[7] ));
  xobna2aa1n03x5               g236(.a(new_n112), .b(new_n329), .c(new_n265), .out0(\s[8] ));
  xnrb03aa1n02x5               g237(.a(new_n121), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


