// Benchmark "adder" written by ABC on Thu Jul 18 14:49:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n330, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  norp02aa1n09x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  tech160nm_finand02aa1n05x5   g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nor022aa1n16x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  tech160nm_fiaoi012aa1n03p5x5 g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  nand02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n12x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor002aa1n06x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oaih12aa1n04x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n107));
  oai012aa1n12x5               g012(.a(new_n101), .b(new_n107), .c(new_n105), .o1(new_n108));
  orn002aa1n24x5               g013(.a(\a[7] ), .b(\b[6] ), .o(new_n109));
  nand22aa1n12x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n02x5               g015(.a(new_n109), .b(new_n110), .o1(new_n111));
  xnrc02aa1n03x5               g016(.a(\b[4] ), .b(\a[5] ), .out0(new_n112));
  nor042aa1d18x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor002aa1d24x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand42aa1n06x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nor043aa1n03x5               g022(.a(new_n117), .b(new_n112), .c(new_n111), .o1(new_n118));
  oaib12aa1n03x5               g023(.a(new_n116), .b(new_n115), .c(new_n109), .out0(new_n119));
  nor042aa1n09x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  oai122aa1n02x7               g025(.a(new_n114), .b(new_n113), .c(new_n120), .d(\b[7] ), .e(\a[8] ), .o1(new_n121));
  nanp03aa1n04x5               g026(.a(new_n109), .b(new_n110), .c(new_n116), .o1(new_n122));
  oai012aa1n06x5               g027(.a(new_n119), .b(new_n121), .c(new_n122), .o1(new_n123));
  inv040aa1n04x5               g028(.a(new_n123), .o1(new_n124));
  aob012aa1d15x5               g029(.a(new_n124), .b(new_n108), .c(new_n118), .out0(new_n125));
  nanp02aa1n24x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  tech160nm_fiaoi012aa1n05x5   g031(.a(new_n97), .b(new_n125), .c(new_n126), .o1(new_n127));
  xnrb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand02aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  oai022aa1n02x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  nor002aa1d32x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nano23aa1d15x5               g036(.a(new_n131), .b(new_n97), .c(new_n126), .d(new_n129), .out0(new_n132));
  aoi022aa1n06x5               g037(.a(new_n125), .b(new_n132), .c(new_n129), .d(new_n130), .o1(new_n133));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  inv020aa1n04x5               g039(.a(new_n134), .o1(new_n135));
  nanp02aa1n24x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n133), .b(new_n136), .c(new_n135), .out0(\s[11] ));
  oaoi03aa1n03x5               g042(.a(\a[11] ), .b(\b[10] ), .c(new_n133), .o1(new_n138));
  xorb03aa1n02x5               g043(.a(new_n138), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1d32x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nano23aa1n09x5               g046(.a(new_n134), .b(new_n140), .c(new_n141), .d(new_n136), .out0(new_n142));
  nand22aa1n12x5               g047(.a(new_n142), .b(new_n132), .o1(new_n143));
  inv040aa1d30x5               g048(.a(new_n143), .o1(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n123), .c(new_n108), .d(new_n118), .o1(new_n145));
  oai112aa1n06x5               g050(.a(new_n135), .b(new_n129), .c(new_n97), .d(new_n131), .o1(new_n146));
  nanb03aa1n12x5               g051(.a(new_n140), .b(new_n141), .c(new_n136), .out0(new_n147));
  aoi012aa1d18x5               g052(.a(new_n140), .b(new_n134), .c(new_n141), .o1(new_n148));
  oai012aa1d24x5               g053(.a(new_n148), .b(new_n146), .c(new_n147), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  xorc02aa1n12x5               g055(.a(\a[13] ), .b(\b[12] ), .out0(new_n151));
  xnbna2aa1n03x5               g056(.a(new_n151), .b(new_n145), .c(new_n150), .out0(\s[13] ));
  inv040aa1d32x5               g057(.a(\a[13] ), .o1(new_n153));
  inv040aa1d28x5               g058(.a(\b[12] ), .o1(new_n154));
  nand02aa1d24x5               g059(.a(new_n154), .b(new_n153), .o1(new_n155));
  aob012aa1n03x5               g060(.a(new_n151), .b(new_n145), .c(new_n150), .out0(new_n156));
  nor002aa1n10x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nanp02aa1n24x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  norb02aa1n03x5               g063(.a(new_n158), .b(new_n157), .out0(new_n159));
  xnbna2aa1n03x5               g064(.a(new_n159), .b(new_n156), .c(new_n155), .out0(\s[14] ));
  nand02aa1d28x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nano32aa1d15x5               g066(.a(new_n157), .b(new_n155), .c(new_n158), .d(new_n161), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  oaoi03aa1n09x5               g068(.a(\a[14] ), .b(\b[13] ), .c(new_n155), .o1(new_n164));
  inv000aa1n02x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n04x5               g070(.a(new_n165), .b(new_n163), .c(new_n145), .d(new_n150), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1d28x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nor002aa1n10x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand42aa1d28x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n168), .b(new_n172), .c(new_n166), .d(new_n169), .o1(new_n174));
  norb02aa1n03x4               g079(.a(new_n173), .b(new_n174), .out0(\s[16] ));
  nano23aa1d15x5               g080(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n176));
  nano32aa1d15x5               g081(.a(new_n143), .b(new_n176), .c(new_n151), .d(new_n159), .out0(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n123), .c(new_n108), .d(new_n118), .o1(new_n178));
  aoai13aa1n06x5               g083(.a(new_n176), .b(new_n164), .c(new_n149), .d(new_n162), .o1(new_n179));
  tech160nm_fiaoi012aa1n05x5   g084(.a(new_n170), .b(new_n168), .c(new_n171), .o1(new_n180));
  nand23aa1n06x5               g085(.a(new_n178), .b(new_n179), .c(new_n180), .o1(new_n181));
  xorb03aa1n03x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor002aa1n06x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  nand42aa1n10x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  tech160nm_fiaoi012aa1n05x5   g089(.a(new_n183), .b(new_n181), .c(new_n184), .o1(new_n185));
  xnrb03aa1n03x5               g090(.a(new_n185), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv000aa1n02x5               g091(.a(new_n176), .o1(new_n187));
  oai012aa1n02x7               g092(.a(new_n129), .b(\b[10] ), .c(\a[11] ), .o1(new_n188));
  oab012aa1n02x4               g093(.a(new_n188), .b(new_n131), .c(new_n97), .out0(new_n189));
  nano22aa1n02x4               g094(.a(new_n140), .b(new_n136), .c(new_n141), .out0(new_n190));
  inv020aa1n03x5               g095(.a(new_n148), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n162), .b(new_n191), .c(new_n189), .d(new_n190), .o1(new_n192));
  aoai13aa1n09x5               g097(.a(new_n180), .b(new_n187), .c(new_n192), .d(new_n165), .o1(new_n193));
  nor002aa1n04x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  nand42aa1n20x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nano23aa1n06x5               g100(.a(new_n183), .b(new_n194), .c(new_n195), .d(new_n184), .out0(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n193), .c(new_n125), .d(new_n177), .o1(new_n197));
  oa0012aa1n06x5               g102(.a(new_n195), .b(new_n194), .c(new_n183), .o(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  inv030aa1d32x5               g104(.a(\b[18] ), .o1(new_n200));
  nanb02aa1d36x5               g105(.a(\a[19] ), .b(new_n200), .out0(new_n201));
  nand02aa1d28x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1d10x5               g107(.a(new_n201), .b(new_n202), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n197), .c(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g111(.a(new_n204), .b(new_n198), .c(new_n181), .d(new_n196), .o1(new_n207));
  nor002aa1d32x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1d28x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  tech160nm_fiaoi012aa1n02p5x5 g115(.a(new_n210), .b(new_n207), .c(new_n201), .o1(new_n211));
  tech160nm_fiaoi012aa1n02p5x5 g116(.a(new_n203), .b(new_n197), .c(new_n199), .o1(new_n212));
  nano22aa1n02x4               g117(.a(new_n212), .b(new_n201), .c(new_n210), .out0(new_n213));
  norp02aa1n03x5               g118(.a(new_n211), .b(new_n213), .o1(\s[20] ));
  nona22aa1n09x5               g119(.a(new_n196), .b(new_n210), .c(new_n203), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n193), .c(new_n125), .d(new_n177), .o1(new_n217));
  oai022aa1d24x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  nand03aa1n12x5               g123(.a(new_n218), .b(new_n201), .c(new_n195), .o1(new_n219));
  nanb03aa1d18x5               g124(.a(new_n208), .b(new_n209), .c(new_n202), .out0(new_n220));
  nor042aa1n04x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  aoi012aa1n09x5               g126(.a(new_n208), .b(new_n221), .c(new_n209), .o1(new_n222));
  oai012aa1d24x5               g127(.a(new_n222), .b(new_n219), .c(new_n220), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  xnrc02aa1n12x5               g129(.a(\b[20] ), .b(\a[21] ), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n217), .c(new_n224), .out0(\s[21] ));
  nor042aa1d18x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  inv040aa1n08x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n226), .b(new_n223), .c(new_n181), .d(new_n216), .o1(new_n230));
  xnrc02aa1n12x5               g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  tech160nm_fiaoi012aa1n02p5x5 g136(.a(new_n231), .b(new_n230), .c(new_n229), .o1(new_n232));
  tech160nm_fiaoi012aa1n02p5x5 g137(.a(new_n225), .b(new_n217), .c(new_n224), .o1(new_n233));
  nano22aa1n02x4               g138(.a(new_n233), .b(new_n229), .c(new_n231), .out0(new_n234));
  norp02aa1n03x5               g139(.a(new_n232), .b(new_n234), .o1(\s[22] ));
  nor042aa1n06x5               g140(.a(new_n231), .b(new_n225), .o1(new_n236));
  norb02aa1n03x5               g141(.a(new_n236), .b(new_n215), .out0(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n193), .c(new_n125), .d(new_n177), .o1(new_n238));
  oao003aa1n02x5               g143(.a(\a[22] ), .b(\b[21] ), .c(new_n229), .carry(new_n239));
  inv030aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  aoi012aa1d24x5               g145(.a(new_n240), .b(new_n223), .c(new_n236), .o1(new_n241));
  xnrc02aa1n12x5               g146(.a(\b[22] ), .b(\a[23] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  xnbna2aa1n03x5               g148(.a(new_n243), .b(new_n238), .c(new_n241), .out0(\s[23] ));
  nor042aa1n06x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n241), .o1(new_n247));
  aoai13aa1n03x5               g152(.a(new_n243), .b(new_n247), .c(new_n181), .d(new_n237), .o1(new_n248));
  xnrc02aa1n03x5               g153(.a(\b[23] ), .b(\a[24] ), .out0(new_n249));
  tech160nm_fiaoi012aa1n02p5x5 g154(.a(new_n249), .b(new_n248), .c(new_n246), .o1(new_n250));
  tech160nm_fiaoi012aa1n02p5x5 g155(.a(new_n242), .b(new_n238), .c(new_n241), .o1(new_n251));
  nano22aa1n02x4               g156(.a(new_n251), .b(new_n246), .c(new_n249), .out0(new_n252));
  norp02aa1n03x5               g157(.a(new_n250), .b(new_n252), .o1(\s[24] ));
  nor042aa1n02x5               g158(.a(new_n249), .b(new_n242), .o1(new_n254));
  nano22aa1n03x7               g159(.a(new_n215), .b(new_n236), .c(new_n254), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n193), .c(new_n125), .d(new_n177), .o1(new_n256));
  oai012aa1n02x5               g161(.a(new_n195), .b(\b[18] ), .c(\a[19] ), .o1(new_n257));
  oab012aa1n02x5               g162(.a(new_n257), .b(new_n183), .c(new_n194), .out0(new_n258));
  nano22aa1n03x5               g163(.a(new_n208), .b(new_n202), .c(new_n209), .out0(new_n259));
  inv000aa1n02x5               g164(.a(new_n222), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n236), .b(new_n260), .c(new_n258), .d(new_n259), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n254), .o1(new_n262));
  oao003aa1n03x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n246), .carry(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n261), .d(new_n239), .o1(new_n264));
  inv030aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  xnrc02aa1n12x5               g170(.a(\b[24] ), .b(\a[25] ), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnbna2aa1n03x5               g172(.a(new_n267), .b(new_n256), .c(new_n265), .out0(\s[25] ));
  nor042aa1n03x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n267), .b(new_n264), .c(new_n181), .d(new_n255), .o1(new_n271));
  xnrc02aa1n12x5               g176(.a(\b[25] ), .b(\a[26] ), .out0(new_n272));
  tech160nm_fiaoi012aa1n02p5x5 g177(.a(new_n272), .b(new_n271), .c(new_n270), .o1(new_n273));
  tech160nm_fiaoi012aa1n03p5x5 g178(.a(new_n266), .b(new_n256), .c(new_n265), .o1(new_n274));
  nano22aa1n02x4               g179(.a(new_n274), .b(new_n270), .c(new_n272), .out0(new_n275));
  nor002aa1n02x5               g180(.a(new_n273), .b(new_n275), .o1(\s[26] ));
  norp02aa1n24x5               g181(.a(new_n272), .b(new_n266), .o1(new_n277));
  nano32aa1n03x7               g182(.a(new_n215), .b(new_n277), .c(new_n236), .d(new_n254), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n193), .c(new_n125), .d(new_n177), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .c(new_n270), .carry(new_n280));
  aobi12aa1n06x5               g185(.a(new_n280), .b(new_n264), .c(new_n277), .out0(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n279), .c(new_n281), .out0(\s[27] ));
  nor042aa1n03x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n254), .b(new_n240), .c(new_n223), .d(new_n236), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n277), .o1(new_n287));
  aoai13aa1n06x5               g192(.a(new_n280), .b(new_n287), .c(new_n286), .d(new_n263), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n282), .b(new_n288), .c(new_n181), .d(new_n278), .o1(new_n289));
  xnrc02aa1n12x5               g194(.a(\b[27] ), .b(\a[28] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n289), .c(new_n285), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n282), .o1(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n292), .b(new_n279), .c(new_n281), .o1(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n285), .c(new_n290), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n291), .b(new_n294), .o1(\s[28] ));
  xnrc02aa1n12x5               g200(.a(\b[28] ), .b(\a[29] ), .out0(new_n296));
  norb02aa1d21x5               g201(.a(new_n282), .b(new_n290), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n288), .c(new_n181), .d(new_n278), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n299));
  tech160nm_fiaoi012aa1n02p5x5 g204(.a(new_n296), .b(new_n298), .c(new_n299), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n297), .o1(new_n301));
  tech160nm_fiaoi012aa1n02p5x5 g206(.a(new_n301), .b(new_n279), .c(new_n281), .o1(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n296), .c(new_n299), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n300), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .out0(new_n306));
  norb03aa1n12x5               g211(.a(new_n282), .b(new_n296), .c(new_n290), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n288), .c(new_n181), .d(new_n278), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n299), .carry(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n307), .o1(new_n311));
  tech160nm_fiaoi012aa1n02p5x5 g216(.a(new_n311), .b(new_n279), .c(new_n281), .o1(new_n312));
  nano22aa1n03x5               g217(.a(new_n312), .b(new_n306), .c(new_n309), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n310), .b(new_n313), .o1(\s[30] ));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  norb02aa1n03x4               g220(.a(new_n307), .b(new_n306), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n288), .c(new_n181), .d(new_n278), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .carry(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n315), .b(new_n317), .c(new_n318), .o1(new_n319));
  inv020aa1n02x5               g224(.a(new_n316), .o1(new_n320));
  tech160nm_fiaoi012aa1n02p5x5 g225(.a(new_n320), .b(new_n279), .c(new_n281), .o1(new_n321));
  nano22aa1n03x5               g226(.a(new_n321), .b(new_n315), .c(new_n318), .out0(new_n322));
  norp02aa1n03x5               g227(.a(new_n319), .b(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g229(.a(\a[3] ), .b(\b[2] ), .c(new_n105), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoib12aa1n06x5               g232(.a(new_n120), .b(new_n108), .c(new_n112), .out0(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g234(.a(\a[6] ), .b(\b[5] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aobi12aa1n02x5               g236(.a(new_n109), .b(new_n330), .c(new_n110), .out0(new_n332));
  xnrb03aa1n03x5               g237(.a(new_n332), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g238(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


