// Benchmark "adder" written by ABC on Wed Jul 17 20:54:56 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n313,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n331, new_n332, new_n334, new_n335, new_n336, new_n338, new_n339,
    new_n340, new_n341, new_n343, new_n345, new_n346, new_n347, new_n349,
    new_n350, new_n352, new_n353, new_n354;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand42aa1d28x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand03aa1n04x5               g004(.a(new_n99), .b(\a[1] ), .c(\b[0] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nor002aa1d24x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nano22aa1d15x5               g007(.a(new_n102), .b(new_n99), .c(new_n101), .out0(new_n103));
  oai012aa1n12x5               g008(.a(new_n103), .b(new_n100), .c(new_n98), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nand02aa1d28x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb03aa1n03x5               g011(.a(new_n106), .b(new_n102), .c(new_n105), .out0(new_n107));
  nand42aa1d28x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nor002aa1n20x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  norb03aa1d15x5               g015(.a(new_n108), .b(new_n110), .c(new_n109), .out0(new_n111));
  nand02aa1d28x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand22aa1n02x5               g017(.a(new_n112), .b(new_n106), .o1(new_n113));
  nor002aa1n16x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1d28x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  norb02aa1n06x5               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  nand42aa1n16x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  oai012aa1d24x5               g022(.a(new_n117), .b(\b[5] ), .c(\a[6] ), .o1(new_n118));
  nona23aa1d18x5               g023(.a(new_n111), .b(new_n116), .c(new_n118), .d(new_n113), .out0(new_n119));
  oai012aa1n02x7               g024(.a(new_n108), .b(new_n114), .c(new_n110), .o1(new_n120));
  nano22aa1n03x5               g025(.a(new_n110), .b(new_n108), .c(new_n115), .out0(new_n121));
  nor002aa1d32x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  oai012aa1n12x5               g027(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .o1(new_n123));
  oab012aa1n06x5               g028(.a(new_n123), .b(new_n109), .c(new_n122), .out0(new_n124));
  aobi12aa1n06x5               g029(.a(new_n120), .b(new_n124), .c(new_n121), .out0(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n119), .c(new_n104), .d(new_n107), .o1(new_n126));
  nand42aa1d28x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  aoi012aa1n02x5               g032(.a(new_n97), .b(new_n126), .c(new_n127), .o1(new_n128));
  nor042aa1d18x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  norb02aa1n02x5               g036(.a(new_n127), .b(new_n97), .out0(new_n132));
  nanp02aa1n02x5               g037(.a(new_n126), .b(new_n132), .o1(new_n133));
  nor042aa1n04x5               g038(.a(new_n129), .b(new_n97), .o1(new_n134));
  nanp03aa1n02x5               g039(.a(new_n133), .b(new_n130), .c(new_n134), .o1(new_n135));
  oai012aa1n02x5               g040(.a(new_n135), .b(new_n128), .c(new_n131), .o1(\s[10] ));
  nano23aa1d15x5               g041(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n127), .out0(new_n137));
  nanp02aa1n02x5               g042(.a(new_n126), .b(new_n137), .o1(new_n138));
  oai012aa1n02x5               g043(.a(new_n130), .b(new_n129), .c(new_n97), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nanp02aa1n12x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norb02aa1n09x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n139), .out0(\s[11] ));
  inv040aa1n08x5               g048(.a(new_n140), .o1(new_n144));
  aob012aa1n03x5               g049(.a(new_n142), .b(new_n138), .c(new_n139), .out0(new_n145));
  nor002aa1d32x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n10x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n09x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  nona23aa1n02x4               g053(.a(new_n145), .b(new_n147), .c(new_n146), .d(new_n140), .out0(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n148), .c(new_n145), .d(new_n144), .o1(\s[12] ));
  nand23aa1d12x5               g055(.a(new_n137), .b(new_n142), .c(new_n148), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nanb03aa1d18x5               g057(.a(new_n146), .b(new_n147), .c(new_n141), .out0(new_n153));
  oaih12aa1n12x5               g058(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .o1(new_n154));
  oaoi03aa1n12x5               g059(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n155));
  inv000aa1n04x5               g060(.a(new_n155), .o1(new_n156));
  oai013aa1n09x5               g061(.a(new_n156), .b(new_n153), .c(new_n134), .d(new_n154), .o1(new_n157));
  nor002aa1d32x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand42aa1d28x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n159), .b(new_n158), .out0(new_n160));
  aoai13aa1n02x5               g065(.a(new_n160), .b(new_n157), .c(new_n126), .d(new_n152), .o1(new_n161));
  nano22aa1n02x4               g066(.a(new_n146), .b(new_n141), .c(new_n147), .out0(new_n162));
  oab012aa1n03x5               g067(.a(new_n154), .b(new_n97), .c(new_n129), .out0(new_n163));
  aoi112aa1n02x5               g068(.a(new_n155), .b(new_n160), .c(new_n163), .d(new_n162), .o1(new_n164));
  aobi12aa1n02x5               g069(.a(new_n164), .b(new_n126), .c(new_n152), .out0(new_n165));
  norb02aa1n02x5               g070(.a(new_n161), .b(new_n165), .out0(\s[13] ));
  inv030aa1n04x5               g071(.a(new_n158), .o1(new_n167));
  nor002aa1n06x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand42aa1d28x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  nona23aa1n02x4               g075(.a(new_n161), .b(new_n169), .c(new_n168), .d(new_n158), .out0(new_n171));
  aoai13aa1n02x5               g076(.a(new_n171), .b(new_n170), .c(new_n167), .d(new_n161), .o1(\s[14] ));
  nano23aa1d15x5               g077(.a(new_n158), .b(new_n168), .c(new_n169), .d(new_n159), .out0(new_n173));
  nanp03aa1n02x5               g078(.a(new_n126), .b(new_n152), .c(new_n173), .o1(new_n174));
  aoai13aa1n03x5               g079(.a(new_n173), .b(new_n155), .c(new_n163), .d(new_n162), .o1(new_n175));
  oaoi03aa1n12x5               g080(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(new_n175), .b(new_n177), .o1(new_n178));
  xorc02aa1n12x5               g083(.a(\a[15] ), .b(\b[14] ), .out0(new_n179));
  oaib12aa1n03x5               g084(.a(new_n179), .b(new_n178), .c(new_n174), .out0(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n176), .c(new_n157), .d(new_n173), .o1(new_n181));
  aobi12aa1n02x5               g086(.a(new_n180), .b(new_n181), .c(new_n174), .out0(\s[15] ));
  nor042aa1n06x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  inv020aa1n04x5               g088(.a(new_n183), .o1(new_n184));
  xorc02aa1n12x5               g089(.a(\a[16] ), .b(\b[15] ), .out0(new_n185));
  and002aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o(new_n186));
  oai022aa1n02x5               g091(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n187));
  nona22aa1n02x4               g092(.a(new_n180), .b(new_n186), .c(new_n187), .out0(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n185), .c(new_n180), .d(new_n184), .o1(\s[16] ));
  and002aa1n18x5               g094(.a(new_n185), .b(new_n179), .o(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n176), .c(new_n157), .d(new_n173), .o1(new_n191));
  nano32aa1d12x5               g096(.a(new_n151), .b(new_n185), .c(new_n173), .d(new_n179), .out0(new_n192));
  nanp02aa1n09x5               g097(.a(new_n126), .b(new_n192), .o1(new_n193));
  oaoi03aa1n02x5               g098(.a(\a[16] ), .b(\b[15] ), .c(new_n184), .o1(new_n194));
  inv000aa1n02x5               g099(.a(new_n194), .o1(new_n195));
  nand23aa1d12x5               g100(.a(new_n193), .b(new_n191), .c(new_n195), .o1(new_n196));
  tech160nm_fixorc02aa1n03p5x5 g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  aoi112aa1n02x5               g102(.a(new_n197), .b(new_n194), .c(new_n126), .d(new_n192), .o1(new_n198));
  aoi022aa1n02x5               g103(.a(new_n196), .b(new_n197), .c(new_n198), .d(new_n191), .o1(\s[17] ));
  norp02aa1n12x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  nor042aa1n06x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand02aa1d12x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nanb02aa1n06x5               g107(.a(new_n201), .b(new_n202), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n200), .c(new_n196), .d(new_n197), .o1(new_n204));
  nona22aa1n02x4               g109(.a(new_n202), .b(new_n201), .c(new_n200), .out0(new_n205));
  aoai13aa1n02x5               g110(.a(new_n204), .b(new_n205), .c(new_n197), .d(new_n196), .o1(\s[18] ));
  norb02aa1n06x5               g111(.a(new_n197), .b(new_n203), .out0(new_n207));
  oa0012aa1n02x5               g112(.a(new_n202), .b(new_n201), .c(new_n200), .o(new_n208));
  xorc02aa1n12x5               g113(.a(\a[19] ), .b(\b[18] ), .out0(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n208), .c(new_n196), .d(new_n207), .o1(new_n210));
  aoi112aa1n02x7               g115(.a(new_n209), .b(new_n208), .c(new_n196), .d(new_n207), .o1(new_n211));
  norb02aa1n03x4               g116(.a(new_n210), .b(new_n211), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g118(.a(\a[19] ), .o1(new_n214));
  inv000aa1d48x5               g119(.a(\b[18] ), .o1(new_n215));
  nand22aa1n04x5               g120(.a(new_n215), .b(new_n214), .o1(new_n216));
  nor042aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanp02aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  nano22aa1n02x4               g124(.a(new_n217), .b(new_n216), .c(new_n218), .out0(new_n220));
  nanp02aa1n03x5               g125(.a(new_n210), .b(new_n220), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n219), .c(new_n216), .d(new_n210), .o1(\s[20] ));
  and003aa1n06x5               g127(.a(new_n207), .b(new_n219), .c(new_n209), .o(new_n223));
  nanp02aa1n02x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  nano22aa1n03x7               g129(.a(new_n217), .b(new_n224), .c(new_n218), .out0(new_n225));
  oai012aa1n06x5               g130(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .o1(new_n226));
  oab012aa1n06x5               g131(.a(new_n226), .b(new_n200), .c(new_n201), .out0(new_n227));
  oaoi03aa1n03x5               g132(.a(\a[20] ), .b(\b[19] ), .c(new_n216), .o1(new_n228));
  tech160nm_fiao0012aa1n02p5x5 g133(.a(new_n228), .b(new_n227), .c(new_n225), .o(new_n229));
  nor042aa1d18x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nanp02aa1n04x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n229), .c(new_n196), .d(new_n223), .o1(new_n233));
  aoi112aa1n02x5               g138(.a(new_n228), .b(new_n232), .c(new_n227), .d(new_n225), .o1(new_n234));
  aobi12aa1n02x5               g139(.a(new_n234), .b(new_n196), .c(new_n223), .out0(new_n235));
  norb02aa1n03x4               g140(.a(new_n233), .b(new_n235), .out0(\s[21] ));
  inv000aa1d42x5               g141(.a(new_n230), .o1(new_n237));
  nor042aa1n06x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nand42aa1n16x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n238), .out0(new_n240));
  norb03aa1n02x5               g145(.a(new_n239), .b(new_n230), .c(new_n238), .out0(new_n241));
  nanp02aa1n03x5               g146(.a(new_n233), .b(new_n241), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n240), .c(new_n237), .d(new_n233), .o1(\s[22] ));
  nano23aa1n09x5               g148(.a(new_n230), .b(new_n238), .c(new_n239), .d(new_n231), .out0(new_n244));
  inv020aa1n03x5               g149(.a(new_n244), .o1(new_n245));
  nano32aa1n02x4               g150(.a(new_n245), .b(new_n207), .c(new_n209), .d(new_n219), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n244), .b(new_n228), .c(new_n227), .d(new_n225), .o1(new_n247));
  oai012aa1d24x5               g152(.a(new_n239), .b(new_n238), .c(new_n230), .o1(new_n248));
  nanp02aa1n02x5               g153(.a(new_n247), .b(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(new_n196), .d(new_n246), .o1(new_n251));
  nanb02aa1n02x5               g156(.a(new_n250), .b(new_n248), .out0(new_n252));
  aoi122aa1n02x7               g157(.a(new_n252), .b(new_n229), .c(new_n244), .d(new_n196), .e(new_n246), .o1(new_n253));
  norb02aa1n03x4               g158(.a(new_n251), .b(new_n253), .out0(\s[23] ));
  norp02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  tech160nm_fixorc02aa1n05x5   g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  oai022aa1n02x5               g162(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(\a[24] ), .c(\b[23] ), .o1(new_n259));
  nanp02aa1n03x5               g164(.a(new_n251), .b(new_n259), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n257), .c(new_n256), .d(new_n251), .o1(\s[24] ));
  nano22aa1n03x7               g166(.a(new_n245), .b(new_n250), .c(new_n257), .out0(new_n262));
  and002aa1n06x5               g167(.a(new_n223), .b(new_n262), .o(new_n263));
  and002aa1n02x5               g168(.a(new_n257), .b(new_n250), .o(new_n264));
  inv030aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  aob012aa1n02x5               g170(.a(new_n258), .b(\b[23] ), .c(\a[24] ), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n265), .c(new_n247), .d(new_n248), .o1(new_n267));
  tech160nm_fixorc02aa1n03p5x5 g172(.a(\a[25] ), .b(\b[24] ), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n267), .c(new_n196), .d(new_n263), .o1(new_n269));
  nanb02aa1n02x5               g174(.a(new_n268), .b(new_n266), .out0(new_n270));
  aoi122aa1n02x7               g175(.a(new_n270), .b(new_n249), .c(new_n264), .d(new_n196), .e(new_n263), .o1(new_n271));
  norb02aa1n03x4               g176(.a(new_n269), .b(new_n271), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  xorc02aa1n02x5               g179(.a(\a[26] ), .b(\b[25] ), .out0(new_n275));
  nanp02aa1n02x5               g180(.a(\b[25] ), .b(\a[26] ), .o1(new_n276));
  oai022aa1n02x5               g181(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n277));
  norb02aa1n02x5               g182(.a(new_n276), .b(new_n277), .out0(new_n278));
  nanp02aa1n03x5               g183(.a(new_n269), .b(new_n278), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n275), .c(new_n274), .d(new_n269), .o1(\s[26] ));
  and002aa1n02x5               g185(.a(new_n275), .b(new_n268), .o(new_n281));
  nand23aa1n06x5               g186(.a(new_n223), .b(new_n262), .c(new_n281), .o1(new_n282));
  inv040aa1n06x5               g187(.a(new_n282), .o1(new_n283));
  nand02aa1d08x5               g188(.a(new_n196), .b(new_n283), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n190), .o1(new_n285));
  tech160nm_fiaoi012aa1n04x5   g190(.a(new_n285), .b(new_n175), .c(new_n177), .o1(new_n286));
  aoi112aa1n03x5               g191(.a(new_n286), .b(new_n194), .c(new_n126), .d(new_n192), .o1(new_n287));
  aoi022aa1n09x5               g192(.a(new_n267), .b(new_n281), .c(new_n276), .d(new_n277), .o1(new_n288));
  tech160nm_fioai012aa1n04x5   g193(.a(new_n288), .b(new_n287), .c(new_n282), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[27] ), .b(\b[26] ), .out0(new_n290));
  aoi122aa1n02x5               g195(.a(new_n290), .b(new_n276), .c(new_n277), .d(new_n267), .e(new_n281), .o1(new_n291));
  aoi022aa1n02x5               g196(.a(new_n289), .b(new_n290), .c(new_n291), .d(new_n284), .o1(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  nand42aa1n02x5               g199(.a(new_n289), .b(new_n290), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .out0(new_n296));
  inv000aa1d42x5               g201(.a(new_n290), .o1(new_n297));
  oai022aa1d24x5               g202(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n298));
  aoi012aa1n02x5               g203(.a(new_n298), .b(\a[28] ), .c(\b[27] ), .o1(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n297), .c(new_n284), .d(new_n288), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n294), .o1(\s[28] ));
  and002aa1n06x5               g206(.a(new_n296), .b(new_n290), .o(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  inv000aa1d42x5               g208(.a(\b[27] ), .o1(new_n304));
  oaib12aa1n09x5               g209(.a(new_n298), .b(new_n304), .c(\a[28] ), .out0(new_n305));
  inv000aa1d42x5               g210(.a(new_n305), .o1(new_n306));
  tech160nm_fixorc02aa1n03p5x5 g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n307), .b(new_n306), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n303), .c(new_n284), .d(new_n288), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n307), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n289), .d(new_n302), .o1(new_n311));
  nanp02aa1n03x5               g216(.a(new_n311), .b(new_n309), .o1(\s[29] ));
  nanp02aa1n02x5               g217(.a(\b[0] ), .b(\a[1] ), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g219(.a(new_n310), .b(new_n290), .c(new_n296), .out0(new_n315));
  tech160nm_fioaoi03aa1n03p5x5 g220(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .o1(new_n316));
  xnrc02aa1n02x5               g221(.a(\b[29] ), .b(\a[30] ), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n316), .c(new_n289), .d(new_n315), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n315), .o1(new_n319));
  norp02aa1n02x5               g224(.a(new_n316), .b(new_n317), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n284), .d(new_n288), .o1(new_n321));
  nanp02aa1n03x5               g226(.a(new_n318), .b(new_n321), .o1(\s[30] ));
  nano32aa1n03x7               g227(.a(new_n317), .b(new_n307), .c(new_n296), .d(new_n290), .out0(new_n323));
  aoi012aa1n02x5               g228(.a(new_n320), .b(\a[30] ), .c(\b[29] ), .o1(new_n324));
  xnrc02aa1n02x5               g229(.a(\b[30] ), .b(\a[31] ), .out0(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n324), .c(new_n289), .d(new_n323), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n323), .o1(new_n327));
  norp02aa1n02x5               g232(.a(new_n324), .b(new_n325), .o1(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n327), .c(new_n284), .d(new_n288), .o1(new_n329));
  nanp02aa1n03x5               g234(.a(new_n326), .b(new_n329), .o1(\s[31] ));
  oai012aa1n02x5               g235(.a(new_n99), .b(new_n98), .c(new_n313), .o1(new_n331));
  oaib12aa1n02x5               g236(.a(new_n331), .b(new_n102), .c(new_n101), .out0(new_n332));
  and002aa1n02x5               g237(.a(new_n104), .b(new_n332), .o(\s[3] ));
  inv000aa1d42x5               g238(.a(new_n102), .o1(new_n334));
  nanp02aa1n02x5               g239(.a(new_n104), .b(new_n107), .o1(new_n335));
  norb02aa1n02x5               g240(.a(new_n106), .b(new_n105), .out0(new_n336));
  aoai13aa1n02x5               g241(.a(new_n335), .b(new_n336), .c(new_n104), .d(new_n334), .o1(\s[4] ));
  nano22aa1n02x4               g242(.a(new_n109), .b(new_n106), .c(new_n117), .out0(new_n338));
  nanp02aa1n03x5               g243(.a(new_n335), .b(new_n338), .o1(new_n339));
  inv000aa1d42x5               g244(.a(new_n109), .o1(new_n340));
  aoi022aa1n02x5               g245(.a(new_n335), .b(new_n106), .c(new_n117), .d(new_n340), .o1(new_n341));
  norb02aa1n02x5               g246(.a(new_n339), .b(new_n341), .out0(\s[5] ));
  norb02aa1n02x5               g247(.a(new_n112), .b(new_n122), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n339), .c(new_n340), .out0(\s[6] ));
  and003aa1n02x5               g249(.a(new_n339), .b(new_n340), .c(new_n343), .o(new_n345));
  aoi112aa1n03x5               g250(.a(new_n345), .b(new_n123), .c(\a[7] ), .d(\b[6] ), .o1(new_n346));
  aoi012aa1n02x5               g251(.a(new_n345), .b(\a[6] ), .c(\b[5] ), .o1(new_n347));
  oab012aa1n02x4               g252(.a(new_n346), .b(new_n347), .c(new_n116), .out0(\s[7] ));
  norb03aa1n02x5               g253(.a(new_n108), .b(new_n114), .c(new_n110), .out0(new_n349));
  obai22aa1n02x7               g254(.a(new_n108), .b(new_n110), .c(new_n346), .d(new_n114), .out0(new_n350));
  oaib12aa1n02x5               g255(.a(new_n350), .b(new_n346), .c(new_n349), .out0(\s[8] ));
  aoi012aa1n02x5               g256(.a(new_n119), .b(new_n104), .c(new_n107), .o1(new_n352));
  oaib12aa1n02x5               g257(.a(new_n120), .b(new_n97), .c(new_n127), .out0(new_n353));
  aoi012aa1n02x5               g258(.a(new_n353), .b(new_n124), .c(new_n121), .o1(new_n354));
  aboi22aa1n03x5               g259(.a(new_n352), .b(new_n354), .c(new_n126), .d(new_n132), .out0(\s[9] ));
endmodule


