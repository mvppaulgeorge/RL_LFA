// Benchmark "adder" written by ABC on Wed Jul 17 20:25:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n305, new_n308, new_n310, new_n312;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  and002aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o(new_n98));
  inv040aa1d30x5               g003(.a(\a[3] ), .o1(new_n99));
  inv040aa1d32x5               g004(.a(\b[2] ), .o1(new_n100));
  tech160nm_finand02aa1n03p5x5 g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  tech160nm_finand02aa1n03p5x5 g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand22aa1n03x5               g007(.a(new_n101), .b(new_n102), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand42aa1n08x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand42aa1n20x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  aoi012aa1n12x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[4] ), .o1(new_n108));
  aboi22aa1n06x5               g013(.a(\b[3] ), .b(new_n108), .c(new_n99), .d(new_n100), .out0(new_n109));
  oaoi13aa1n12x5               g014(.a(new_n98), .b(new_n109), .c(new_n107), .d(new_n103), .o1(new_n110));
  nor022aa1n08x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  tech160nm_finand02aa1n03p5x5 g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nor022aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n113), .b(new_n112), .c(new_n114), .d(new_n111), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  tech160nm_fixnrc02aa1n02p5x5 g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nor043aa1n04x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  oai012aa1n02x5               g023(.a(new_n112), .b(new_n114), .c(new_n111), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[5] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[4] ), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  oaib12aa1n09x5               g028(.a(new_n119), .b(new_n115), .c(new_n123), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n127), .b(new_n126), .c(new_n97), .out0(\s[10] ));
  aobi12aa1n06x5               g033(.a(new_n127), .b(new_n126), .c(new_n97), .out0(new_n129));
  nor042aa1n12x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nand42aa1d28x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  oaoi03aa1n12x5               g037(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n133));
  tech160nm_fioai012aa1n04x5   g038(.a(new_n132), .b(new_n129), .c(new_n133), .o1(new_n134));
  norp03aa1n02x5               g039(.a(new_n129), .b(new_n132), .c(new_n133), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n130), .o1(new_n137));
  nor042aa1n06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand42aa1n16x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n138), .b(new_n139), .out0(new_n140));
  nand43aa1n02x5               g045(.a(new_n134), .b(new_n137), .c(new_n140), .o1(new_n141));
  tech160nm_fiaoi012aa1n03p5x5 g046(.a(new_n140), .b(new_n134), .c(new_n137), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(\s[12] ));
  nano23aa1d15x5               g048(.a(new_n130), .b(new_n138), .c(new_n139), .d(new_n131), .out0(new_n144));
  nand23aa1d12x5               g049(.a(new_n144), .b(new_n125), .c(new_n127), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  aoai13aa1n06x5               g051(.a(new_n146), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n147));
  aoi112aa1n02x5               g052(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n148));
  aoi112aa1n03x5               g053(.a(new_n148), .b(new_n138), .c(new_n144), .d(new_n133), .o1(new_n149));
  xnrc02aa1n12x5               g054(.a(\b[12] ), .b(\a[13] ), .out0(new_n150));
  xobna2aa1n03x5               g055(.a(new_n150), .b(new_n147), .c(new_n149), .out0(\s[13] ));
  orn002aa1n03x5               g056(.a(\a[13] ), .b(\b[12] ), .o(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n150), .c(new_n147), .d(new_n149), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xnrc02aa1n02x5               g059(.a(\b[13] ), .b(\a[14] ), .out0(new_n155));
  norp02aa1n02x5               g060(.a(new_n155), .b(new_n150), .o1(new_n156));
  inv000aa1n02x5               g061(.a(new_n156), .o1(new_n157));
  oao003aa1n03x5               g062(.a(\a[14] ), .b(\b[13] ), .c(new_n152), .carry(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n157), .c(new_n147), .d(new_n149), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n06x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nand42aa1n06x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  norp02aa1n06x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nand42aa1n04x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n165), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  nano23aa1n02x4               g073(.a(new_n161), .b(new_n163), .c(new_n164), .d(new_n162), .out0(new_n169));
  nona22aa1n03x5               g074(.a(new_n169), .b(new_n155), .c(new_n150), .out0(new_n170));
  nor042aa1n09x5               g075(.a(new_n170), .b(new_n145), .o1(new_n171));
  aoai13aa1n12x5               g076(.a(new_n171), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n172));
  nand22aa1n03x5               g077(.a(new_n144), .b(new_n133), .o1(new_n173));
  nona22aa1n03x5               g078(.a(new_n173), .b(new_n148), .c(new_n138), .out0(new_n174));
  nona23aa1n03x5               g079(.a(new_n164), .b(new_n162), .c(new_n161), .d(new_n163), .out0(new_n175));
  nor043aa1n02x5               g080(.a(new_n175), .b(new_n155), .c(new_n150), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n163), .b(new_n161), .c(new_n164), .o1(new_n177));
  tech160nm_fioai012aa1n04x5   g082(.a(new_n177), .b(new_n158), .c(new_n175), .o1(new_n178));
  aoi012aa1n12x5               g083(.a(new_n178), .b(new_n174), .c(new_n176), .o1(new_n179));
  xorc02aa1n02x5               g084(.a(\a[17] ), .b(\b[16] ), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n172), .c(new_n179), .out0(\s[17] ));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  nand02aa1n03x5               g088(.a(new_n183), .b(new_n182), .o1(new_n184));
  oai012aa1n02x5               g089(.a(new_n109), .b(new_n107), .c(new_n103), .o1(new_n185));
  oaib12aa1n02x5               g090(.a(new_n185), .b(new_n108), .c(\b[3] ), .out0(new_n186));
  inv000aa1n02x5               g091(.a(new_n124), .o1(new_n187));
  oaib12aa1n06x5               g092(.a(new_n187), .b(new_n186), .c(new_n118), .out0(new_n188));
  oabi12aa1n03x5               g093(.a(new_n178), .b(new_n149), .c(new_n170), .out0(new_n189));
  aoai13aa1n02x5               g094(.a(new_n180), .b(new_n189), .c(new_n188), .d(new_n171), .o1(new_n190));
  nor002aa1d24x5               g095(.a(\b[17] ), .b(\a[18] ), .o1(new_n191));
  nanp02aa1n12x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nanb02aa1n12x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  xobna2aa1n03x5               g098(.a(new_n193), .b(new_n190), .c(new_n184), .out0(\s[18] ));
  nanp02aa1n02x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  nano22aa1d15x5               g100(.a(new_n193), .b(new_n184), .c(new_n195), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n192), .b(new_n191), .c(new_n182), .d(new_n183), .o1(new_n198));
  aoai13aa1n04x5               g103(.a(new_n198), .b(new_n197), .c(new_n172), .d(new_n179), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nanp02aa1n04x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nor042aa1n06x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand02aa1n06x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  norb02aa1n02x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  aoi112aa1n02x5               g111(.a(new_n206), .b(new_n202), .c(new_n199), .d(new_n203), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n206), .b(new_n202), .c(new_n199), .d(new_n203), .o1(new_n208));
  norb02aa1n02x7               g113(.a(new_n208), .b(new_n207), .out0(\s[20] ));
  nano23aa1n09x5               g114(.a(new_n202), .b(new_n204), .c(new_n205), .d(new_n203), .out0(new_n210));
  nanp02aa1n02x5               g115(.a(new_n196), .b(new_n210), .o1(new_n211));
  nona23aa1n09x5               g116(.a(new_n205), .b(new_n203), .c(new_n202), .d(new_n204), .out0(new_n212));
  aoi012aa1n09x5               g117(.a(new_n204), .b(new_n202), .c(new_n205), .o1(new_n213));
  oai012aa1n18x5               g118(.a(new_n213), .b(new_n212), .c(new_n198), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n04x5               g120(.a(new_n215), .b(new_n211), .c(new_n172), .d(new_n179), .o1(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  xorc02aa1n02x5               g123(.a(\a[21] ), .b(\b[20] ), .out0(new_n219));
  xorc02aa1n02x5               g124(.a(\a[22] ), .b(\b[21] ), .out0(new_n220));
  aoi112aa1n02x5               g125(.a(new_n218), .b(new_n220), .c(new_n216), .d(new_n219), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n220), .b(new_n218), .c(new_n216), .d(new_n219), .o1(new_n222));
  norb02aa1n02x7               g127(.a(new_n222), .b(new_n221), .out0(\s[22] ));
  inv000aa1d42x5               g128(.a(\a[21] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\a[22] ), .o1(new_n225));
  xroi22aa1d06x4               g130(.a(new_n224), .b(\b[20] ), .c(new_n225), .d(\b[21] ), .out0(new_n226));
  nanp03aa1n03x5               g131(.a(new_n226), .b(new_n196), .c(new_n210), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\b[21] ), .o1(new_n228));
  oaoi03aa1n09x5               g133(.a(new_n225), .b(new_n228), .c(new_n218), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoi012aa1n02x5               g135(.a(new_n230), .b(new_n214), .c(new_n226), .o1(new_n231));
  aoai13aa1n04x5               g136(.a(new_n231), .b(new_n227), .c(new_n172), .d(new_n179), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  xorc02aa1n03x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  xorc02aa1n02x5               g140(.a(\a[24] ), .b(\b[23] ), .out0(new_n236));
  aoi112aa1n02x5               g141(.a(new_n234), .b(new_n236), .c(new_n232), .d(new_n235), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n234), .c(new_n232), .d(new_n235), .o1(new_n238));
  norb02aa1n02x7               g143(.a(new_n238), .b(new_n237), .out0(\s[24] ));
  nanp02aa1n09x5               g144(.a(new_n172), .b(new_n179), .o1(new_n240));
  and002aa1n09x5               g145(.a(new_n236), .b(new_n235), .o(new_n241));
  inv000aa1n02x5               g146(.a(new_n241), .o1(new_n242));
  norp02aa1n02x5               g147(.a(new_n227), .b(new_n242), .o1(new_n243));
  inv040aa1n02x5               g148(.a(new_n198), .o1(new_n244));
  inv020aa1n03x5               g149(.a(new_n213), .o1(new_n245));
  aoai13aa1n06x5               g150(.a(new_n226), .b(new_n245), .c(new_n210), .d(new_n244), .o1(new_n246));
  orn002aa1n02x5               g151(.a(\a[23] ), .b(\b[22] ), .o(new_n247));
  oao003aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .c(new_n247), .carry(new_n248));
  aoai13aa1n04x5               g153(.a(new_n248), .b(new_n242), .c(new_n246), .d(new_n229), .o1(new_n249));
  tech160nm_fixorc02aa1n05x5   g154(.a(\a[25] ), .b(\b[24] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(new_n240), .d(new_n243), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(new_n250), .b(new_n249), .c(new_n240), .d(new_n243), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(\s[25] ));
  nor042aa1n03x5               g158(.a(\b[24] ), .b(\a[25] ), .o1(new_n254));
  tech160nm_fixorc02aa1n05x5   g159(.a(\a[26] ), .b(\b[25] ), .out0(new_n255));
  nona22aa1n02x5               g160(.a(new_n251), .b(new_n255), .c(new_n254), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n254), .o1(new_n257));
  aobi12aa1n06x5               g162(.a(new_n255), .b(new_n251), .c(new_n257), .out0(new_n258));
  norb02aa1n03x4               g163(.a(new_n256), .b(new_n258), .out0(\s[26] ));
  and002aa1n06x5               g164(.a(new_n255), .b(new_n250), .o(new_n260));
  nano22aa1n03x7               g165(.a(new_n227), .b(new_n241), .c(new_n260), .out0(new_n261));
  aoai13aa1n04x5               g166(.a(new_n261), .b(new_n189), .c(new_n188), .d(new_n171), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[26] ), .b(\b[25] ), .c(new_n257), .carry(new_n263));
  aobi12aa1n06x5               g168(.a(new_n263), .b(new_n249), .c(new_n260), .out0(new_n264));
  xorc02aa1n12x5               g169(.a(\a[27] ), .b(\b[26] ), .out0(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n264), .c(new_n262), .out0(\s[27] ));
  norp02aa1n02x5               g171(.a(\b[26] ), .b(\a[27] ), .o1(new_n267));
  inv040aa1n03x5               g172(.a(new_n267), .o1(new_n268));
  aobi12aa1n02x7               g173(.a(new_n265), .b(new_n264), .c(new_n262), .out0(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[27] ), .b(\a[28] ), .out0(new_n270));
  nano22aa1n03x5               g175(.a(new_n269), .b(new_n268), .c(new_n270), .out0(new_n271));
  aobi12aa1n06x5               g176(.a(new_n261), .b(new_n172), .c(new_n179), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n241), .b(new_n230), .c(new_n214), .d(new_n226), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n260), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n263), .b(new_n274), .c(new_n273), .d(new_n248), .o1(new_n275));
  oaih12aa1n02x5               g180(.a(new_n265), .b(new_n275), .c(new_n272), .o1(new_n276));
  tech160nm_fiaoi012aa1n02p5x5 g181(.a(new_n270), .b(new_n276), .c(new_n268), .o1(new_n277));
  norp02aa1n03x5               g182(.a(new_n277), .b(new_n271), .o1(\s[28] ));
  xnrc02aa1n02x5               g183(.a(\b[28] ), .b(\a[29] ), .out0(new_n279));
  norb02aa1n02x5               g184(.a(new_n265), .b(new_n270), .out0(new_n280));
  oaih12aa1n02x5               g185(.a(new_n280), .b(new_n275), .c(new_n272), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[28] ), .b(\b[27] ), .c(new_n268), .carry(new_n282));
  tech160nm_fiaoi012aa1n02p5x5 g187(.a(new_n279), .b(new_n281), .c(new_n282), .o1(new_n283));
  aobi12aa1n03x5               g188(.a(new_n280), .b(new_n264), .c(new_n262), .out0(new_n284));
  nano22aa1n03x5               g189(.a(new_n284), .b(new_n279), .c(new_n282), .out0(new_n285));
  norp02aa1n03x5               g190(.a(new_n283), .b(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g191(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g192(.a(new_n265), .b(new_n279), .c(new_n270), .out0(new_n288));
  oaih12aa1n02x5               g193(.a(new_n288), .b(new_n275), .c(new_n272), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[29] ), .b(\b[28] ), .c(new_n282), .carry(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[29] ), .b(\a[30] ), .out0(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  aobi12aa1n03x5               g197(.a(new_n288), .b(new_n264), .c(new_n262), .out0(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n291), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[30] ));
  xnrc02aa1n02x5               g200(.a(\b[30] ), .b(\a[31] ), .out0(new_n296));
  norb02aa1n02x5               g201(.a(new_n288), .b(new_n291), .out0(new_n297));
  aobi12aa1n02x7               g202(.a(new_n297), .b(new_n264), .c(new_n262), .out0(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n290), .carry(new_n299));
  nano22aa1n03x5               g204(.a(new_n298), .b(new_n296), .c(new_n299), .out0(new_n300));
  oaih12aa1n02x5               g205(.a(new_n297), .b(new_n275), .c(new_n272), .o1(new_n301));
  tech160nm_fiaoi012aa1n02p5x5 g206(.a(new_n296), .b(new_n301), .c(new_n299), .o1(new_n302));
  norp02aa1n03x5               g207(.a(new_n302), .b(new_n300), .o1(\s[31] ));
  xnbna2aa1n03x5               g208(.a(new_n107), .b(new_n101), .c(new_n102), .out0(\s[3] ));
  oaoi03aa1n02x5               g209(.a(\a[3] ), .b(\b[2] ), .c(new_n107), .o1(new_n305));
  xorb03aa1n02x5               g210(.a(new_n305), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g211(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g212(.a(new_n120), .b(new_n121), .c(new_n110), .o1(new_n308));
  xnrb03aa1n02x5               g213(.a(new_n308), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g214(.a(\a[6] ), .b(\b[5] ), .c(new_n308), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g216(.a(new_n114), .b(new_n310), .c(new_n113), .o1(new_n312));
  xnrb03aa1n02x5               g217(.a(new_n312), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g218(.a(new_n188), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


