// Benchmark "adder" written by ABC on Thu Jul 18 05:05:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n311, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n333, new_n335, new_n336, new_n337, new_n339,
    new_n340, new_n341, new_n342, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n351, new_n353, new_n354, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixnrc02aa1n04x5   g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\a[9] ), .b(new_n98), .out0(new_n99));
  oai112aa1n06x5               g004(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n100));
  nand22aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand22aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  techfinor002aa1n02p5x5       g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  aoi113aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n100), .d(new_n103), .e(new_n101), .o1(new_n105));
  nand22aa1n12x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  inv000aa1n02x5               g011(.a(new_n106), .o1(new_n107));
  oai022aa1d18x5               g012(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n108));
  nor002aa1n02x5               g013(.a(new_n108), .b(new_n107), .o1(new_n109));
  xorc02aa1n12x5               g014(.a(\a[6] ), .b(\b[5] ), .out0(new_n110));
  inv000aa1d42x5               g015(.a(\b[3] ), .o1(new_n111));
  obai22aa1d24x5               g016(.a(\a[4] ), .b(new_n111), .c(\b[4] ), .d(\a[5] ), .out0(new_n112));
  nand42aa1d28x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nand02aa1d08x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nano22aa1n03x7               g019(.a(new_n112), .b(new_n113), .c(new_n114), .out0(new_n115));
  nand23aa1n02x5               g020(.a(new_n115), .b(new_n109), .c(new_n110), .o1(new_n116));
  nor042aa1d18x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  inv000aa1n06x5               g022(.a(new_n117), .o1(new_n118));
  oaoi03aa1n02x5               g023(.a(\a[6] ), .b(\b[5] ), .c(new_n118), .o1(new_n119));
  nor042aa1n02x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nor002aa1n20x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nano23aa1n03x7               g026(.a(new_n121), .b(new_n120), .c(new_n114), .d(new_n106), .out0(new_n122));
  aoi022aa1n06x5               g027(.a(new_n122), .b(new_n119), .c(new_n108), .d(new_n114), .o1(new_n123));
  oai012aa1n18x5               g028(.a(new_n123), .b(new_n116), .c(new_n105), .o1(new_n124));
  oaib12aa1n09x5               g029(.a(new_n124), .b(new_n98), .c(\a[9] ), .out0(new_n125));
  xobna2aa1n03x5               g030(.a(new_n97), .b(new_n125), .c(new_n99), .out0(\s[10] ));
  nand42aa1n04x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nor002aa1d32x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n127), .b(new_n128), .out0(new_n129));
  oai022aa1d18x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  aboi22aa1n03x5               g035(.a(new_n130), .b(new_n125), .c(\b[9] ), .d(\a[10] ), .out0(new_n131));
  aoi022aa1d24x5               g036(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n128), .out0(new_n133));
  oaib12aa1n06x5               g038(.a(new_n133), .b(new_n130), .c(new_n125), .out0(new_n134));
  oa0012aa1n03x5               g039(.a(new_n134), .b(new_n131), .c(new_n129), .o(\s[11] ));
  inv000aa1d42x5               g040(.a(new_n128), .o1(new_n136));
  nor002aa1n06x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanp02aa1n12x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  nor042aa1n02x5               g044(.a(new_n137), .b(new_n128), .o1(new_n140));
  nanp03aa1n02x5               g045(.a(new_n134), .b(new_n138), .c(new_n140), .o1(new_n141));
  aoai13aa1n03x5               g046(.a(new_n141), .b(new_n139), .c(new_n136), .d(new_n134), .o1(\s[12] ));
  nano23aa1n06x5               g047(.a(new_n137), .b(new_n128), .c(new_n138), .d(new_n127), .out0(new_n143));
  xorc02aa1n12x5               g048(.a(\a[9] ), .b(\b[8] ), .out0(new_n144));
  nanb03aa1d24x5               g049(.a(new_n97), .b(new_n143), .c(new_n144), .out0(new_n145));
  inv000aa1n02x5               g050(.a(new_n145), .o1(new_n146));
  nand02aa1d06x5               g051(.a(new_n124), .b(new_n146), .o1(new_n147));
  aob012aa1n03x5               g052(.a(new_n140), .b(new_n130), .c(new_n132), .out0(new_n148));
  nanp02aa1n02x5               g053(.a(new_n148), .b(new_n138), .o1(new_n149));
  xorc02aa1n12x5               g054(.a(\a[13] ), .b(\b[12] ), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n147), .c(new_n149), .out0(\s[13] ));
  inv040aa1d32x5               g056(.a(\a[13] ), .o1(new_n152));
  inv000aa1d42x5               g057(.a(\b[12] ), .o1(new_n153));
  nanp02aa1n04x5               g058(.a(new_n153), .b(new_n152), .o1(new_n154));
  nand02aa1d06x5               g059(.a(new_n147), .b(new_n149), .o1(new_n155));
  nand42aa1n02x5               g060(.a(new_n155), .b(new_n150), .o1(new_n156));
  tech160nm_fixorc02aa1n03p5x5 g061(.a(\a[14] ), .b(\b[13] ), .out0(new_n157));
  nand42aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  oai022aa1n09x5               g063(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n159));
  nanb03aa1n03x5               g064(.a(new_n159), .b(new_n156), .c(new_n158), .out0(new_n160));
  aoai13aa1n03x5               g065(.a(new_n160), .b(new_n157), .c(new_n154), .d(new_n156), .o1(\s[14] ));
  and002aa1n02x5               g066(.a(new_n157), .b(new_n150), .o(new_n162));
  oaoi03aa1n02x5               g067(.a(\a[14] ), .b(\b[13] ), .c(new_n154), .o1(new_n163));
  nor042aa1n09x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand42aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n163), .c(new_n155), .d(new_n162), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n167), .b(new_n163), .c(new_n155), .d(new_n162), .o1(new_n169));
  norb02aa1n03x4               g074(.a(new_n168), .b(new_n169), .out0(\s[15] ));
  inv000aa1d42x5               g075(.a(new_n164), .o1(new_n171));
  nor042aa1n06x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand02aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  inv000aa1d42x5               g079(.a(new_n172), .o1(new_n175));
  oai112aa1n02x5               g080(.a(new_n175), .b(new_n173), .c(\b[14] ), .d(\a[15] ), .o1(new_n176));
  nanb02aa1n03x5               g081(.a(new_n176), .b(new_n168), .out0(new_n177));
  aoai13aa1n03x5               g082(.a(new_n177), .b(new_n174), .c(new_n171), .d(new_n168), .o1(\s[16] ));
  nano23aa1n03x7               g083(.a(new_n164), .b(new_n172), .c(new_n173), .d(new_n165), .out0(new_n179));
  nano32aa1d12x5               g084(.a(new_n145), .b(new_n179), .c(new_n150), .d(new_n157), .out0(new_n180));
  nanp02aa1n09x5               g085(.a(new_n124), .b(new_n180), .o1(new_n181));
  nano22aa1n03x5               g086(.a(new_n172), .b(new_n165), .c(new_n173), .out0(new_n182));
  oai022aa1n02x7               g087(.a(new_n152), .b(new_n153), .c(\b[13] ), .d(\a[14] ), .o1(new_n183));
  oaih12aa1n02x5               g088(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .o1(new_n184));
  nano23aa1n02x5               g089(.a(new_n183), .b(new_n184), .c(new_n154), .d(new_n138), .out0(new_n185));
  nand03aa1n02x5               g090(.a(new_n185), .b(new_n148), .c(new_n182), .o1(new_n186));
  aoi022aa1n02x7               g091(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n187));
  aoai13aa1n02x5               g092(.a(new_n187), .b(new_n164), .c(new_n159), .d(new_n158), .o1(new_n188));
  nand23aa1n09x5               g093(.a(new_n186), .b(new_n175), .c(new_n188), .o1(new_n189));
  nanb02aa1n12x5               g094(.a(new_n189), .b(new_n181), .out0(new_n190));
  xorc02aa1n12x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  nano32aa1n02x4               g096(.a(new_n191), .b(new_n186), .c(new_n188), .d(new_n175), .out0(new_n192));
  aoi022aa1n02x5               g097(.a(new_n190), .b(new_n191), .c(new_n181), .d(new_n192), .o1(\s[17] ));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  nanb02aa1d36x5               g099(.a(\b[16] ), .b(new_n194), .out0(new_n195));
  aoai13aa1n06x5               g100(.a(new_n191), .b(new_n189), .c(new_n124), .d(new_n180), .o1(new_n196));
  nor042aa1n04x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nand22aa1n04x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  norb02aa1n06x4               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  nano22aa1n02x4               g104(.a(new_n197), .b(new_n195), .c(new_n198), .out0(new_n200));
  nanp02aa1n02x5               g105(.a(new_n196), .b(new_n200), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n201), .b(new_n199), .c(new_n195), .d(new_n196), .o1(\s[18] ));
  and002aa1n02x5               g107(.a(new_n191), .b(new_n199), .o(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n189), .c(new_n124), .d(new_n180), .o1(new_n204));
  oaoi03aa1n12x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n195), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  nor002aa1d32x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand42aa1n20x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n06x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n204), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n08x5               g116(.a(new_n207), .o1(new_n212));
  aob012aa1n03x5               g117(.a(new_n209), .b(new_n204), .c(new_n206), .out0(new_n213));
  nor002aa1n10x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand42aa1n20x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  norb02aa1n06x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  norb03aa1n02x5               g121(.a(new_n215), .b(new_n207), .c(new_n214), .out0(new_n217));
  nand42aa1n02x5               g122(.a(new_n213), .b(new_n217), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n216), .c(new_n212), .d(new_n213), .o1(\s[20] ));
  nano23aa1n09x5               g124(.a(new_n207), .b(new_n214), .c(new_n215), .d(new_n208), .out0(new_n220));
  nand23aa1n04x5               g125(.a(new_n220), .b(new_n191), .c(new_n199), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoi112aa1n09x5               g127(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n223));
  oai112aa1n04x5               g128(.a(new_n209), .b(new_n216), .c(new_n223), .d(new_n197), .o1(new_n224));
  oaoi03aa1n09x5               g129(.a(\a[20] ), .b(\b[19] ), .c(new_n212), .o1(new_n225));
  inv030aa1n02x5               g130(.a(new_n225), .o1(new_n226));
  nanp02aa1n02x5               g131(.a(new_n224), .b(new_n226), .o1(new_n227));
  nor002aa1n16x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  nand42aa1n06x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  norb02aa1n09x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  aoai13aa1n04x5               g135(.a(new_n230), .b(new_n227), .c(new_n190), .d(new_n222), .o1(new_n231));
  nona22aa1n02x4               g136(.a(new_n224), .b(new_n225), .c(new_n230), .out0(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n190), .c(new_n222), .o1(new_n233));
  norb02aa1n03x4               g138(.a(new_n231), .b(new_n233), .out0(\s[21] ));
  inv000aa1n02x5               g139(.a(new_n228), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[21] ), .b(\a[22] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  oai022aa1n02x5               g142(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(\a[22] ), .c(\b[21] ), .o1(new_n239));
  nanp02aa1n03x5               g144(.a(new_n231), .b(new_n239), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n237), .c(new_n235), .d(new_n231), .o1(\s[22] ));
  nanb02aa1n12x5               g146(.a(new_n236), .b(new_n230), .out0(new_n242));
  nano32aa1n02x4               g147(.a(new_n242), .b(new_n220), .c(new_n199), .d(new_n191), .out0(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n189), .c(new_n124), .d(new_n180), .o1(new_n244));
  aob012aa1n03x5               g149(.a(new_n238), .b(\b[21] ), .c(\a[22] ), .out0(new_n245));
  aoai13aa1n12x5               g150(.a(new_n245), .b(new_n242), .c(new_n224), .d(new_n226), .o1(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[23] ), .b(\b[22] ), .out0(new_n248));
  aob012aa1n03x5               g153(.a(new_n248), .b(new_n244), .c(new_n247), .out0(new_n249));
  nano22aa1n03x7               g154(.a(new_n236), .b(new_n235), .c(new_n229), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n225), .c(new_n220), .d(new_n205), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n248), .o1(new_n252));
  and003aa1n02x5               g157(.a(new_n251), .b(new_n252), .c(new_n245), .o(new_n253));
  aobi12aa1n02x7               g158(.a(new_n249), .b(new_n253), .c(new_n244), .out0(\s[23] ));
  nor022aa1n16x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  inv040aa1n15x5               g160(.a(new_n255), .o1(new_n256));
  xorc02aa1n02x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  oai022aa1n02x5               g162(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(\a[24] ), .c(\b[23] ), .o1(new_n259));
  aoai13aa1n02x5               g164(.a(new_n259), .b(new_n252), .c(new_n244), .d(new_n247), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n257), .c(new_n249), .d(new_n256), .o1(\s[24] ));
  nand42aa1n03x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  tech160nm_fixnrc02aa1n05x5   g167(.a(\b[23] ), .b(\a[24] ), .out0(new_n263));
  nano22aa1n09x5               g168(.a(new_n263), .b(new_n256), .c(new_n262), .out0(new_n264));
  nano22aa1n02x5               g169(.a(new_n221), .b(new_n250), .c(new_n264), .out0(new_n265));
  inv000aa1d42x5               g170(.a(new_n264), .o1(new_n266));
  oaoi03aa1n02x5               g171(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n266), .c(new_n251), .d(new_n245), .o1(new_n269));
  tech160nm_fixorc02aa1n03p5x5 g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n269), .c(new_n190), .d(new_n265), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(new_n270), .b(new_n267), .c(new_n246), .d(new_n264), .o1(new_n272));
  aobi12aa1n02x5               g177(.a(new_n272), .b(new_n190), .c(new_n265), .out0(new_n273));
  norb02aa1n03x4               g178(.a(new_n271), .b(new_n273), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  tech160nm_fixorc02aa1n02p5x5 g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  nanp02aa1n02x5               g182(.a(\b[25] ), .b(\a[26] ), .o1(new_n278));
  oai022aa1n02x5               g183(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n279));
  norb02aa1n02x5               g184(.a(new_n278), .b(new_n279), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n271), .b(new_n280), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n277), .c(new_n276), .d(new_n271), .o1(\s[26] ));
  and002aa1n02x5               g187(.a(new_n277), .b(new_n270), .o(new_n283));
  nano32aa1d12x5               g188(.a(new_n221), .b(new_n283), .c(new_n250), .d(new_n264), .out0(new_n284));
  aoai13aa1n12x5               g189(.a(new_n284), .b(new_n189), .c(new_n124), .d(new_n180), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n283), .b(new_n267), .c(new_n246), .d(new_n264), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(new_n279), .b(new_n278), .o1(new_n287));
  nand23aa1n06x5               g192(.a(new_n285), .b(new_n286), .c(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  aoi122aa1n02x5               g194(.a(new_n289), .b(new_n278), .c(new_n279), .d(new_n269), .e(new_n283), .o1(new_n290));
  aoi022aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n288), .d(new_n289), .o1(\s[27] ));
  nor002aa1n03x5               g196(.a(\b[26] ), .b(\a[27] ), .o1(new_n292));
  nor042aa1n03x5               g197(.a(\b[27] ), .b(\a[28] ), .o1(new_n293));
  and002aa1n12x5               g198(.a(\b[27] ), .b(\a[28] ), .o(new_n294));
  norp02aa1n02x5               g199(.a(new_n294), .b(new_n293), .o1(new_n295));
  inv000aa1n03x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n292), .c(new_n288), .d(new_n289), .o1(new_n297));
  aoi022aa1n03x5               g202(.a(new_n269), .b(new_n283), .c(new_n278), .d(new_n279), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n289), .o1(new_n299));
  norp03aa1n02x5               g204(.a(new_n294), .b(new_n293), .c(new_n292), .o1(new_n300));
  aoai13aa1n02x5               g205(.a(new_n300), .b(new_n299), .c(new_n298), .d(new_n285), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n297), .b(new_n301), .o1(\s[28] ));
  norb02aa1n03x5               g207(.a(new_n289), .b(new_n296), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n288), .b(new_n303), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n303), .o1(new_n305));
  aoib12aa1n06x5               g210(.a(new_n293), .b(new_n292), .c(new_n294), .out0(new_n306));
  aoai13aa1n02x7               g211(.a(new_n306), .b(new_n305), .c(new_n298), .d(new_n285), .o1(new_n307));
  xorc02aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .out0(new_n308));
  norb02aa1n02x5               g213(.a(new_n306), .b(new_n308), .out0(new_n309));
  aoi022aa1n03x5               g214(.a(new_n307), .b(new_n308), .c(new_n304), .d(new_n309), .o1(\s[29] ));
  nanp02aa1n02x5               g215(.a(\b[0] ), .b(\a[1] ), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g217(.a(new_n308), .b(new_n289), .c(new_n295), .o1(new_n313));
  nanb02aa1n03x5               g218(.a(new_n313), .b(new_n288), .out0(new_n314));
  xorc02aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .out0(new_n315));
  norp02aa1n02x5               g220(.a(\b[28] ), .b(\a[29] ), .o1(new_n316));
  aoi012aa1n02x5               g221(.a(new_n306), .b(\a[29] ), .c(\b[28] ), .o1(new_n317));
  norp03aa1n02x5               g222(.a(new_n317), .b(new_n315), .c(new_n316), .o1(new_n318));
  tech160nm_fioaoi03aa1n03p5x5 g223(.a(\a[29] ), .b(\b[28] ), .c(new_n306), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n319), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n313), .c(new_n298), .d(new_n285), .o1(new_n321));
  aoi022aa1n03x5               g226(.a(new_n321), .b(new_n315), .c(new_n314), .d(new_n318), .o1(\s[30] ));
  nand03aa1n02x5               g227(.a(new_n303), .b(new_n308), .c(new_n315), .o1(new_n323));
  nanb02aa1n03x5               g228(.a(new_n323), .b(new_n288), .out0(new_n324));
  xorc02aa1n02x5               g229(.a(\a[31] ), .b(\b[30] ), .out0(new_n325));
  inv000aa1d42x5               g230(.a(\a[30] ), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\b[29] ), .o1(new_n327));
  oabi12aa1n02x5               g232(.a(new_n325), .b(\a[30] ), .c(\b[29] ), .out0(new_n328));
  oaoi13aa1n02x5               g233(.a(new_n328), .b(new_n319), .c(new_n326), .d(new_n327), .o1(new_n329));
  tech160nm_fioaoi03aa1n02p5x5 g234(.a(new_n326), .b(new_n327), .c(new_n319), .o1(new_n330));
  aoai13aa1n02x7               g235(.a(new_n330), .b(new_n323), .c(new_n298), .d(new_n285), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n331), .b(new_n325), .c(new_n324), .d(new_n329), .o1(\s[31] ));
  nanb02aa1n02x5               g237(.a(new_n102), .b(new_n103), .out0(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n100), .c(new_n101), .out0(\s[3] ));
  inv000aa1n06x5               g239(.a(new_n105), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[4] ), .b(\b[3] ), .out0(new_n336));
  aoi113aa1n02x5               g241(.a(new_n336), .b(new_n102), .c(new_n100), .d(new_n103), .e(new_n101), .o1(new_n337));
  aoi012aa1n02x5               g242(.a(new_n337), .b(new_n335), .c(new_n336), .o1(\s[4] ));
  inv000aa1d42x5               g243(.a(new_n113), .o1(new_n339));
  nona22aa1d18x5               g244(.a(new_n335), .b(new_n112), .c(new_n339), .out0(new_n340));
  inv000aa1d42x5               g245(.a(new_n340), .o1(new_n341));
  oaib12aa1n02x5               g246(.a(new_n335), .b(new_n111), .c(\a[4] ), .out0(new_n342));
  oaoi13aa1n02x5               g247(.a(new_n341), .b(new_n342), .c(new_n117), .d(new_n339), .o1(\s[5] ));
  xnbna2aa1n03x5               g248(.a(new_n110), .b(new_n340), .c(new_n118), .out0(\s[6] ));
  and002aa1n02x5               g249(.a(\b[5] ), .b(\a[6] ), .o(new_n345));
  nand23aa1n04x5               g250(.a(new_n340), .b(new_n110), .c(new_n118), .o1(new_n346));
  nona32aa1n03x5               g251(.a(new_n346), .b(new_n345), .c(new_n121), .d(new_n107), .out0(new_n347));
  inv000aa1d42x5               g252(.a(new_n121), .o1(new_n348));
  aboi22aa1n03x5               g253(.a(new_n345), .b(new_n346), .c(new_n106), .d(new_n348), .out0(new_n349));
  norb02aa1n02x5               g254(.a(new_n347), .b(new_n349), .out0(\s[7] ));
  norb02aa1n02x5               g255(.a(new_n114), .b(new_n120), .out0(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n351), .b(new_n347), .c(new_n348), .out0(\s[8] ));
  inv000aa1d42x5               g257(.a(new_n144), .o1(new_n353));
  aoi122aa1n02x5               g258(.a(new_n353), .b(new_n108), .c(new_n114), .d(new_n122), .e(new_n119), .o1(new_n354));
  oai012aa1n02x5               g259(.a(new_n354), .b(new_n116), .c(new_n105), .o1(new_n355));
  aob012aa1n02x5               g260(.a(new_n355), .b(new_n124), .c(new_n353), .out0(\s[9] ));
endmodule


