// Benchmark "adder" written by ABC on Wed Jul 17 17:28:54 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n318, new_n319,
    new_n321, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d28x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor002aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  tech160nm_fioai012aa1n04x5   g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand02aa1d04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norp02aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  aoi012aa1n02x5               g013(.a(new_n104), .b(new_n106), .c(new_n105), .o1(new_n109));
  tech160nm_fioai012aa1n05x5   g014(.a(new_n109), .b(new_n108), .c(new_n103), .o1(new_n110));
  xorc02aa1n02x5               g015(.a(\a[5] ), .b(\b[4] ), .out0(new_n111));
  nanp02aa1n12x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  inv000aa1n02x5               g017(.a(new_n112), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  orn002aa1n02x5               g020(.a(\a[7] ), .b(\b[6] ), .o(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n115), .c(new_n113), .d(new_n114), .out0(new_n117));
  tech160nm_fixorc02aa1n02p5x5 g022(.a(\a[6] ), .b(\b[5] ), .out0(new_n118));
  nano22aa1n03x7               g023(.a(new_n117), .b(new_n111), .c(new_n118), .out0(new_n119));
  nanp02aa1n03x5               g024(.a(new_n119), .b(new_n110), .o1(new_n120));
  orn002aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .o(new_n121));
  nanp02aa1n02x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  nanp03aa1n02x5               g028(.a(new_n123), .b(new_n115), .c(new_n122), .o1(new_n124));
  aoi013aa1n06x4               g029(.a(new_n113), .b(new_n124), .c(new_n116), .d(new_n121), .o1(new_n125));
  inv000aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  tech160nm_fixnrc02aa1n05x5   g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n99), .b(new_n127), .c(new_n120), .d(new_n126), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n16x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1d28x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  nanb02aa1n02x5               g037(.a(new_n132), .b(new_n128), .out0(new_n133));
  aoai13aa1n12x5               g038(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n134));
  nand02aa1d28x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor042aa1n12x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  inv040aa1n02x5               g043(.a(new_n134), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n135), .o1(new_n140));
  nona32aa1n02x4               g045(.a(new_n133), .b(new_n136), .c(new_n140), .d(new_n139), .out0(new_n141));
  nor042aa1n06x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand22aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  aob012aa1n02x5               g049(.a(new_n144), .b(new_n141), .c(new_n135), .out0(new_n145));
  nona22aa1n02x4               g050(.a(new_n141), .b(new_n144), .c(new_n140), .out0(new_n146));
  nanp02aa1n02x5               g051(.a(new_n145), .b(new_n146), .o1(\s[12] ));
  nano23aa1d15x5               g052(.a(new_n142), .b(new_n136), .c(new_n143), .d(new_n135), .out0(new_n148));
  nona22aa1d18x5               g053(.a(new_n148), .b(new_n127), .c(new_n132), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n125), .c(new_n119), .d(new_n110), .o1(new_n151));
  nona23aa1n09x5               g056(.a(new_n135), .b(new_n143), .c(new_n142), .d(new_n136), .out0(new_n152));
  ao0012aa1n03x5               g057(.a(new_n142), .b(new_n136), .c(new_n143), .o(new_n153));
  oabi12aa1n18x5               g058(.a(new_n153), .b(new_n152), .c(new_n134), .out0(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n151), .b(new_n155), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nand42aa1n06x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nor042aa1n04x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  aoi012aa1n02x5               g064(.a(new_n159), .b(new_n156), .c(new_n158), .o1(new_n160));
  xnrb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand42aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nano23aa1d15x5               g068(.a(new_n162), .b(new_n159), .c(new_n163), .d(new_n158), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  oaih12aa1n06x5               g070(.a(new_n163), .b(new_n162), .c(new_n159), .o1(new_n166));
  aoai13aa1n04x5               g071(.a(new_n166), .b(new_n165), .c(new_n151), .d(new_n155), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand02aa1n06x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nor042aa1n03x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nanp02aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(new_n173), .b(new_n170), .c(new_n167), .d(new_n169), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n173), .b(new_n170), .c(new_n167), .d(new_n169), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[16] ));
  nano23aa1d15x5               g081(.a(new_n171), .b(new_n170), .c(new_n172), .d(new_n169), .out0(new_n177));
  nano22aa1d15x5               g082(.a(new_n149), .b(new_n164), .c(new_n177), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n125), .c(new_n119), .d(new_n110), .o1(new_n179));
  inv000aa1d42x5               g084(.a(new_n166), .o1(new_n180));
  aoai13aa1n12x5               g085(.a(new_n177), .b(new_n180), .c(new_n154), .d(new_n164), .o1(new_n181));
  aoi012aa1n02x5               g086(.a(new_n171), .b(new_n170), .c(new_n172), .o1(new_n182));
  nanp03aa1d12x5               g087(.a(new_n179), .b(new_n181), .c(new_n182), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[18] ), .o1(new_n185));
  inv040aa1d32x5               g090(.a(\a[17] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[16] ), .o1(new_n187));
  tech160nm_fioaoi03aa1n03p5x5 g092(.a(new_n186), .b(new_n187), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  nand42aa1n04x5               g094(.a(new_n120), .b(new_n126), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n177), .o1(new_n191));
  aoai13aa1n04x5               g096(.a(new_n164), .b(new_n153), .c(new_n148), .d(new_n139), .o1(new_n192));
  aoai13aa1n06x5               g097(.a(new_n182), .b(new_n191), .c(new_n192), .d(new_n166), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n186), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n194), .b(new_n193), .c(new_n190), .d(new_n178), .o1(new_n195));
  oai022aa1n02x7               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oaib12aa1n12x5               g101(.a(new_n196), .b(new_n185), .c(\b[17] ), .out0(new_n197));
  nand02aa1n08x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nor042aa1d18x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g108(.a(new_n187), .b(new_n186), .o1(new_n204));
  oaoi03aa1n12x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n205));
  aoai13aa1n09x5               g110(.a(new_n201), .b(new_n205), .c(new_n183), .d(new_n194), .o1(new_n206));
  nor042aa1n04x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nand02aa1n16x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nanb02aa1n02x5               g113(.a(new_n207), .b(new_n208), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nona22aa1n03x5               g115(.a(new_n206), .b(new_n210), .c(new_n199), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n199), .o1(new_n212));
  tech160nm_fiaoi012aa1n05x5   g117(.a(new_n209), .b(new_n206), .c(new_n212), .o1(new_n213));
  norb02aa1n03x4               g118(.a(new_n211), .b(new_n213), .out0(\s[20] ));
  nano23aa1n09x5               g119(.a(new_n207), .b(new_n199), .c(new_n208), .d(new_n198), .out0(new_n215));
  nand02aa1d04x5               g120(.a(new_n194), .b(new_n215), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n193), .c(new_n190), .d(new_n178), .o1(new_n218));
  nona23aa1n09x5               g123(.a(new_n198), .b(new_n208), .c(new_n207), .d(new_n199), .out0(new_n219));
  aoi012aa1n12x5               g124(.a(new_n207), .b(new_n199), .c(new_n208), .o1(new_n220));
  oai012aa1d24x5               g125(.a(new_n220), .b(new_n219), .c(new_n197), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  tech160nm_finand02aa1n05x5   g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nor042aa1n06x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  norb02aa1n02x7               g129(.a(new_n223), .b(new_n224), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n218), .c(new_n222), .out0(\s[21] ));
  inv000aa1n06x5               g131(.a(new_n224), .o1(new_n227));
  inv000aa1n02x5               g132(.a(new_n225), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n218), .c(new_n222), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[21] ), .b(\a[22] ), .out0(new_n230));
  nano22aa1n02x4               g135(.a(new_n229), .b(new_n227), .c(new_n230), .out0(new_n231));
  aoai13aa1n03x5               g136(.a(new_n225), .b(new_n221), .c(new_n183), .d(new_n217), .o1(new_n232));
  aoi012aa1n03x5               g137(.a(new_n230), .b(new_n232), .c(new_n227), .o1(new_n233));
  norp02aa1n03x5               g138(.a(new_n233), .b(new_n231), .o1(\s[22] ));
  nona32aa1n09x5               g139(.a(new_n183), .b(new_n230), .c(new_n228), .d(new_n216), .out0(new_n235));
  nano22aa1n03x7               g140(.a(new_n230), .b(new_n223), .c(new_n227), .out0(new_n236));
  oao003aa1n06x5               g141(.a(\a[22] ), .b(\b[21] ), .c(new_n227), .carry(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(new_n221), .c(new_n236), .o1(new_n239));
  tech160nm_fixnrc02aa1n05x5   g144(.a(\b[22] ), .b(\a[23] ), .out0(new_n240));
  xobna2aa1n03x5               g145(.a(new_n240), .b(new_n235), .c(new_n239), .out0(\s[23] ));
  and002aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o(new_n242));
  xorc02aa1n12x5               g147(.a(\a[24] ), .b(\b[23] ), .out0(new_n243));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(new_n244), .b(new_n238), .c(new_n221), .d(new_n236), .o1(new_n245));
  aoai13aa1n02x7               g150(.a(new_n243), .b(new_n242), .c(new_n235), .d(new_n245), .o1(new_n246));
  aoi112aa1n06x5               g151(.a(new_n243), .b(new_n242), .c(new_n235), .d(new_n245), .o1(new_n247));
  nanb02aa1n03x5               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  norb02aa1n02x5               g153(.a(new_n243), .b(new_n240), .out0(new_n249));
  inv020aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  nano32aa1n02x4               g155(.a(new_n250), .b(new_n194), .c(new_n236), .d(new_n215), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n193), .c(new_n190), .d(new_n178), .o1(new_n252));
  inv020aa1n03x5               g157(.a(new_n220), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n236), .b(new_n253), .c(new_n215), .d(new_n205), .o1(new_n254));
  orn002aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .o(new_n255));
  oao003aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n255), .carry(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n250), .c(new_n254), .d(new_n237), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[24] ), .b(\a[25] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n252), .c(new_n258), .out0(\s[25] ));
  nor042aa1n03x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoi012aa1n02x7               g168(.a(new_n259), .b(new_n252), .c(new_n258), .o1(new_n264));
  xnrc02aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  nano22aa1n03x7               g170(.a(new_n264), .b(new_n263), .c(new_n265), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n260), .b(new_n257), .c(new_n183), .d(new_n251), .o1(new_n267));
  aoi012aa1n03x5               g172(.a(new_n265), .b(new_n267), .c(new_n263), .o1(new_n268));
  nor002aa1n02x5               g173(.a(new_n268), .b(new_n266), .o1(\s[26] ));
  nor042aa1n02x5               g174(.a(new_n265), .b(new_n259), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  nano23aa1n06x5               g176(.a(new_n216), .b(new_n271), .c(new_n249), .d(new_n236), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n193), .c(new_n190), .d(new_n178), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n274));
  aobi12aa1n12x5               g179(.a(new_n274), .b(new_n257), .c(new_n270), .out0(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  norb02aa1n02x5               g182(.a(new_n277), .b(new_n276), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n273), .c(new_n275), .out0(\s[27] ));
  inv000aa1n06x5               g184(.a(new_n276), .o1(new_n280));
  xnrc02aa1n02x5               g185(.a(\b[27] ), .b(\a[28] ), .out0(new_n281));
  aobi12aa1n06x5               g186(.a(new_n277), .b(new_n273), .c(new_n275), .out0(new_n282));
  nano22aa1n03x7               g187(.a(new_n282), .b(new_n280), .c(new_n281), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n249), .b(new_n238), .c(new_n221), .d(new_n236), .o1(new_n284));
  aoai13aa1n04x5               g189(.a(new_n274), .b(new_n271), .c(new_n284), .d(new_n256), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n277), .b(new_n285), .c(new_n183), .d(new_n272), .o1(new_n286));
  aoi012aa1n03x5               g191(.a(new_n281), .b(new_n286), .c(new_n280), .o1(new_n287));
  nor002aa1n02x5               g192(.a(new_n287), .b(new_n283), .o1(\s[28] ));
  nano22aa1n02x4               g193(.a(new_n281), .b(new_n280), .c(new_n277), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n285), .c(new_n183), .d(new_n272), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[28] ), .b(\a[29] ), .out0(new_n292));
  aoi012aa1n03x5               g197(.a(new_n292), .b(new_n290), .c(new_n291), .o1(new_n293));
  aobi12aa1n06x5               g198(.a(new_n289), .b(new_n273), .c(new_n275), .out0(new_n294));
  nano22aa1n03x7               g199(.a(new_n294), .b(new_n291), .c(new_n292), .out0(new_n295));
  norp02aa1n03x5               g200(.a(new_n293), .b(new_n295), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g202(.a(new_n278), .b(new_n292), .c(new_n281), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n285), .c(new_n183), .d(new_n272), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n300));
  xnrc02aa1n02x5               g205(.a(\b[29] ), .b(\a[30] ), .out0(new_n301));
  aoi012aa1n03x5               g206(.a(new_n301), .b(new_n299), .c(new_n300), .o1(new_n302));
  aobi12aa1n06x5               g207(.a(new_n298), .b(new_n273), .c(new_n275), .out0(new_n303));
  nano22aa1n03x7               g208(.a(new_n303), .b(new_n300), .c(new_n301), .out0(new_n304));
  nor002aa1n02x5               g209(.a(new_n302), .b(new_n304), .o1(\s[30] ));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  norb03aa1n02x5               g211(.a(new_n289), .b(new_n301), .c(new_n292), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n285), .c(new_n183), .d(new_n272), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n309));
  aoi012aa1n03x5               g214(.a(new_n306), .b(new_n308), .c(new_n309), .o1(new_n310));
  aobi12aa1n06x5               g215(.a(new_n307), .b(new_n273), .c(new_n275), .out0(new_n311));
  nano22aa1n03x7               g216(.a(new_n311), .b(new_n306), .c(new_n309), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n310), .b(new_n312), .o1(\s[31] ));
  xnrb03aa1n02x5               g218(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g219(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g221(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai112aa1n02x5               g222(.a(new_n109), .b(new_n111), .c(new_n108), .d(new_n103), .o1(new_n318));
  aob012aa1n02x5               g223(.a(new_n318), .b(\b[4] ), .c(\a[5] ), .out0(new_n319));
  xnrc02aa1n02x5               g224(.a(new_n319), .b(new_n118), .out0(\s[6] ));
  aob012aa1n02x5               g225(.a(new_n122), .b(new_n319), .c(new_n118), .out0(new_n321));
  xnbna2aa1n03x5               g226(.a(new_n321), .b(new_n115), .c(new_n116), .out0(\s[7] ));
  oaoi03aa1n02x5               g227(.a(\a[7] ), .b(\b[6] ), .c(new_n321), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g229(.a(new_n127), .b(new_n120), .c(new_n126), .out0(\s[9] ));
endmodule


