// Benchmark "adder" written by ABC on Wed Jul 17 19:03:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n337, new_n340,
    new_n341, new_n342, new_n344, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  oa0022aa1n06x5               g003(.a(\a[6] ), .b(\b[5] ), .c(\a[5] ), .d(\b[4] ), .o(new_n99));
  inv040aa1d32x5               g004(.a(\a[7] ), .o1(new_n100));
  inv030aa1d32x5               g005(.a(\b[6] ), .o1(new_n101));
  nand42aa1n04x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nand42aa1n02x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  aoi022aa1d24x5               g008(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n104));
  nanp03aa1n02x5               g009(.a(new_n104), .b(new_n102), .c(new_n103), .o1(new_n105));
  oaoi03aa1n03x5               g010(.a(\a[8] ), .b(\b[7] ), .c(new_n102), .o1(new_n106));
  oab012aa1n04x5               g011(.a(new_n106), .b(new_n105), .c(new_n99), .out0(new_n107));
  and002aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .o(new_n108));
  nano32aa1n03x7               g013(.a(new_n108), .b(new_n104), .c(new_n102), .d(new_n103), .out0(new_n109));
  and002aa1n12x5               g014(.a(\b[0] ), .b(\a[1] ), .o(new_n110));
  oaoi03aa1n09x5               g015(.a(\a[2] ), .b(\b[1] ), .c(new_n110), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nand22aa1n06x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  norp02aa1n24x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  nand02aa1n03x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  tech160nm_fiaoi012aa1n05x5   g021(.a(new_n112), .b(new_n114), .c(new_n113), .o1(new_n117));
  inv000aa1n02x5               g022(.a(new_n117), .o1(new_n118));
  aoai13aa1n06x5               g023(.a(new_n109), .b(new_n118), .c(new_n116), .d(new_n111), .o1(new_n119));
  nand02aa1d10x5               g024(.a(new_n119), .b(new_n107), .o1(new_n120));
  oaoi03aa1n09x5               g025(.a(new_n97), .b(new_n98), .c(new_n120), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\a[10] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[9] ), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n123), .b(new_n122), .o1(new_n124));
  nand02aa1d24x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n121), .b(new_n125), .c(new_n124), .out0(\s[10] ));
  nand02aa1d28x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nor002aa1d32x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  norb02aa1d21x5               g033(.a(new_n127), .b(new_n128), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  nand02aa1d04x5               g035(.a(new_n121), .b(new_n124), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n130), .b(new_n131), .c(new_n125), .out0(\s[11] ));
  inv000aa1d42x5               g037(.a(new_n128), .o1(new_n133));
  inv040aa1n02x5               g038(.a(new_n125), .o1(new_n134));
  nona22aa1n03x5               g039(.a(new_n131), .b(new_n130), .c(new_n134), .out0(new_n135));
  nor002aa1n02x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1d28x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aobi12aa1n03x5               g043(.a(new_n138), .b(new_n135), .c(new_n133), .out0(new_n139));
  aoi112aa1n02x7               g044(.a(new_n130), .b(new_n134), .c(new_n121), .d(new_n124), .o1(new_n140));
  norp03aa1n02x5               g045(.a(new_n140), .b(new_n138), .c(new_n128), .o1(new_n141));
  nor002aa1n02x5               g046(.a(new_n139), .b(new_n141), .o1(\s[12] ));
  oai022aa1d24x5               g047(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n143));
  nanb03aa1d24x5               g048(.a(new_n128), .b(new_n125), .c(new_n127), .out0(new_n144));
  nano22aa1n03x7               g049(.a(new_n144), .b(new_n137), .c(new_n143), .out0(new_n145));
  tech160nm_fiaoi012aa1n05x5   g050(.a(new_n136), .b(new_n128), .c(new_n137), .o1(new_n146));
  inv000aa1n03x5               g051(.a(new_n146), .o1(new_n147));
  nor002aa1n02x5               g052(.a(new_n145), .b(new_n147), .o1(new_n148));
  oabi12aa1n02x5               g053(.a(new_n106), .b(new_n99), .c(new_n105), .out0(new_n149));
  inv000aa1d42x5               g054(.a(\a[1] ), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\b[0] ), .o1(new_n151));
  nor002aa1n02x5               g056(.a(\b[1] ), .b(\a[2] ), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(\b[1] ), .b(\a[2] ), .o1(new_n153));
  oaoi13aa1n09x5               g058(.a(new_n152), .b(new_n153), .c(new_n150), .d(new_n151), .o1(new_n154));
  nona23aa1n03x5               g059(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n155));
  tech160nm_fioai012aa1n03p5x5 g060(.a(new_n117), .b(new_n155), .c(new_n154), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[8] ), .b(\a[9] ), .o1(new_n157));
  nano22aa1n03x7               g062(.a(new_n144), .b(new_n157), .c(new_n137), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n149), .c(new_n156), .d(new_n109), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(new_n159), .b(new_n148), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n16x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand02aa1d28x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n162), .b(new_n160), .c(new_n163), .o1(new_n164));
  xnrb03aa1n03x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n09x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanp02aa1n12x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nona23aa1d18x5               g072(.a(new_n167), .b(new_n163), .c(new_n162), .d(new_n166), .out0(new_n168));
  oa0012aa1n02x5               g073(.a(new_n167), .b(new_n166), .c(new_n162), .o(new_n169));
  inv000aa1n02x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n168), .c(new_n159), .d(new_n148), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n09x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nor042aa1n12x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand22aa1n12x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  norb02aa1n09x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  aoi112aa1n02x5               g082(.a(new_n173), .b(new_n177), .c(new_n171), .d(new_n174), .o1(new_n178));
  aoai13aa1n03x5               g083(.a(new_n177), .b(new_n173), .c(new_n171), .d(new_n174), .o1(new_n179));
  norb02aa1n03x4               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  tech160nm_fiaoi012aa1n02p5x5 g085(.a(new_n149), .b(new_n156), .c(new_n109), .o1(new_n181));
  norb02aa1n06x4               g086(.a(new_n174), .b(new_n173), .out0(new_n182));
  nano22aa1n03x7               g087(.a(new_n168), .b(new_n182), .c(new_n177), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n143), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n137), .o1(new_n185));
  nona22aa1n02x4               g090(.a(new_n129), .b(new_n185), .c(new_n134), .out0(new_n186));
  nano32aa1n03x7               g091(.a(new_n186), .b(new_n146), .c(new_n184), .d(new_n157), .out0(new_n187));
  nanp02aa1n02x5               g092(.a(new_n187), .b(new_n183), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n175), .o1(new_n189));
  inv000aa1n02x5               g094(.a(new_n173), .o1(new_n190));
  oai112aa1n03x5               g095(.a(new_n167), .b(new_n174), .c(new_n166), .d(new_n162), .o1(new_n191));
  aob012aa1n06x5               g096(.a(new_n176), .b(new_n191), .c(new_n190), .out0(new_n192));
  nona23aa1n06x5               g097(.a(new_n129), .b(new_n143), .c(new_n185), .d(new_n134), .out0(new_n193));
  nano23aa1n03x7               g098(.a(new_n162), .b(new_n166), .c(new_n167), .d(new_n163), .out0(new_n194));
  nand23aa1n03x5               g099(.a(new_n194), .b(new_n182), .c(new_n177), .o1(new_n195));
  tech160nm_fiaoi012aa1n02p5x5 g100(.a(new_n195), .b(new_n193), .c(new_n146), .o1(new_n196));
  nano22aa1n03x7               g101(.a(new_n196), .b(new_n192), .c(new_n189), .out0(new_n197));
  tech160nm_fioai012aa1n05x5   g102(.a(new_n197), .b(new_n181), .c(new_n188), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nano32aa1n06x5               g104(.a(new_n195), .b(new_n193), .c(new_n158), .d(new_n146), .out0(new_n200));
  oaih12aa1n12x5               g105(.a(new_n183), .b(new_n145), .c(new_n147), .o1(new_n201));
  nand23aa1d12x5               g106(.a(new_n201), .b(new_n189), .c(new_n192), .o1(new_n202));
  aoi012aa1n06x5               g107(.a(new_n202), .b(new_n120), .c(new_n200), .o1(new_n203));
  oaoi03aa1n03x5               g108(.a(\a[17] ), .b(\b[16] ), .c(new_n203), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv000aa1d42x5               g110(.a(\a[17] ), .o1(new_n206));
  inv020aa1n04x5               g111(.a(\a[18] ), .o1(new_n207));
  xroi22aa1d06x4               g112(.a(new_n206), .b(\b[16] ), .c(new_n207), .d(\b[17] ), .out0(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n202), .c(new_n120), .d(new_n200), .o1(new_n209));
  inv040aa1d28x5               g114(.a(\b[17] ), .o1(new_n210));
  oai022aa1d24x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  oaib12aa1n18x5               g116(.a(new_n211), .b(new_n210), .c(\a[18] ), .out0(new_n212));
  xorc02aa1n12x5               g117(.a(\a[19] ), .b(\b[18] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g120(.a(\a[19] ), .o1(new_n216));
  nanb02aa1n09x5               g121(.a(\b[18] ), .b(new_n216), .out0(new_n217));
  inv030aa1n02x5               g122(.a(new_n213), .o1(new_n218));
  aoi012aa1n03x5               g123(.a(new_n218), .b(new_n209), .c(new_n212), .o1(new_n219));
  xnrc02aa1n03x5               g124(.a(\b[19] ), .b(\a[20] ), .out0(new_n220));
  nano22aa1n03x5               g125(.a(new_n219), .b(new_n217), .c(new_n220), .out0(new_n221));
  aoi012aa1n06x5               g126(.a(new_n188), .b(new_n119), .c(new_n107), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n212), .o1(new_n223));
  oaoi13aa1n03x5               g128(.a(new_n223), .b(new_n208), .c(new_n222), .d(new_n202), .o1(new_n224));
  oaoi13aa1n02x7               g129(.a(new_n220), .b(new_n217), .c(new_n224), .d(new_n218), .o1(new_n225));
  nor002aa1n02x5               g130(.a(new_n225), .b(new_n221), .o1(\s[20] ));
  inv040aa1d30x5               g131(.a(\a[21] ), .o1(new_n227));
  nona22aa1d18x5               g132(.a(new_n208), .b(new_n218), .c(new_n220), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  norp02aa1n02x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  inv000aa1n02x5               g135(.a(new_n230), .o1(new_n231));
  and002aa1n02x5               g136(.a(\b[18] ), .b(\a[19] ), .o(new_n232));
  and002aa1n02x5               g137(.a(\b[19] ), .b(\a[20] ), .o(new_n233));
  nand22aa1n03x5               g138(.a(new_n212), .b(new_n217), .o1(new_n234));
  nona22aa1n09x5               g139(.a(new_n234), .b(new_n233), .c(new_n232), .out0(new_n235));
  nanp02aa1n02x5               g140(.a(new_n235), .b(new_n231), .o1(new_n236));
  oaoi13aa1n06x5               g141(.a(new_n236), .b(new_n229), .c(new_n222), .d(new_n202), .o1(new_n237));
  xorb03aa1n02x5               g142(.a(new_n237), .b(\b[20] ), .c(new_n227), .out0(\s[21] ));
  nanb02aa1n02x5               g143(.a(\b[20] ), .b(new_n227), .out0(new_n239));
  inv000aa1n02x5               g144(.a(new_n236), .o1(new_n240));
  xorc02aa1n12x5               g145(.a(\a[21] ), .b(\b[20] ), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  oaoi13aa1n02x7               g147(.a(new_n242), .b(new_n240), .c(new_n203), .d(new_n228), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[22] ), .b(\b[21] ), .out0(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  nano22aa1n03x5               g150(.a(new_n243), .b(new_n239), .c(new_n245), .out0(new_n246));
  oaoi13aa1n03x5               g151(.a(new_n245), .b(new_n239), .c(new_n237), .d(new_n242), .o1(new_n247));
  norp02aa1n03x5               g152(.a(new_n247), .b(new_n246), .o1(\s[22] ));
  inv000aa1d42x5               g153(.a(\a[23] ), .o1(new_n249));
  inv020aa1n04x5               g154(.a(\a[22] ), .o1(new_n250));
  xroi22aa1d06x4               g155(.a(new_n227), .b(\b[20] ), .c(new_n250), .d(\b[21] ), .out0(new_n251));
  nano32aa1n03x7               g156(.a(new_n220), .b(new_n251), .c(new_n208), .d(new_n213), .out0(new_n252));
  nand42aa1n02x5               g157(.a(\b[21] ), .b(\a[22] ), .o1(new_n253));
  aoi112aa1n06x5               g158(.a(new_n233), .b(new_n232), .c(new_n212), .d(new_n217), .o1(new_n254));
  oaih12aa1n02x5               g159(.a(new_n251), .b(new_n254), .c(new_n230), .o1(new_n255));
  oai022aa1d18x5               g160(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n256));
  aob012aa1n03x5               g161(.a(new_n255), .b(new_n256), .c(new_n253), .out0(new_n257));
  oaoi13aa1n04x5               g162(.a(new_n257), .b(new_n252), .c(new_n222), .d(new_n202), .o1(new_n258));
  xorb03aa1n02x5               g163(.a(new_n258), .b(\b[22] ), .c(new_n249), .out0(\s[23] ));
  inv020aa1n03x5               g164(.a(\b[22] ), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(new_n260), .b(new_n249), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n252), .b(new_n202), .c(new_n120), .d(new_n200), .o1(new_n262));
  tech160nm_fixnrc02aa1n03p5x5 g167(.a(\b[22] ), .b(\a[23] ), .out0(new_n263));
  aoib12aa1n03x5               g168(.a(new_n263), .b(new_n262), .c(new_n257), .out0(new_n264));
  xnrc02aa1n03x5               g169(.a(\b[23] ), .b(\a[24] ), .out0(new_n265));
  nano22aa1n03x5               g170(.a(new_n264), .b(new_n261), .c(new_n265), .out0(new_n266));
  oaoi13aa1n02x5               g171(.a(new_n265), .b(new_n261), .c(new_n258), .d(new_n263), .o1(new_n267));
  norp02aa1n03x5               g172(.a(new_n267), .b(new_n266), .o1(\s[24] ));
  nona22aa1n12x5               g173(.a(new_n251), .b(new_n263), .c(new_n265), .out0(new_n269));
  nor042aa1n04x5               g174(.a(new_n228), .b(new_n269), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n202), .c(new_n120), .d(new_n200), .o1(new_n271));
  norp02aa1n02x5               g176(.a(\b[23] ), .b(\a[24] ), .o1(new_n272));
  oai112aa1n03x5               g177(.a(new_n256), .b(new_n253), .c(new_n260), .d(new_n249), .o1(new_n273));
  aoi022aa1n02x5               g178(.a(new_n273), .b(new_n261), .c(\a[24] ), .d(\b[23] ), .o1(new_n274));
  nor042aa1n06x5               g179(.a(new_n274), .b(new_n272), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n275), .b(new_n269), .c(new_n235), .d(new_n231), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  xnrc02aa1n12x5               g182(.a(\b[24] ), .b(\a[25] ), .out0(new_n278));
  xobna2aa1n03x5               g183(.a(new_n278), .b(new_n271), .c(new_n277), .out0(\s[25] ));
  nor042aa1n03x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  tech160nm_fiaoi012aa1n02p5x5 g186(.a(new_n278), .b(new_n271), .c(new_n277), .o1(new_n282));
  xnrc02aa1n06x5               g187(.a(\b[25] ), .b(\a[26] ), .out0(new_n283));
  nano22aa1n02x4               g188(.a(new_n282), .b(new_n281), .c(new_n283), .out0(new_n284));
  oaoi13aa1n03x5               g189(.a(new_n276), .b(new_n270), .c(new_n222), .d(new_n202), .o1(new_n285));
  oaoi13aa1n03x5               g190(.a(new_n283), .b(new_n281), .c(new_n285), .d(new_n278), .o1(new_n286));
  norp02aa1n03x5               g191(.a(new_n286), .b(new_n284), .o1(\s[26] ));
  nor022aa1n04x5               g192(.a(new_n283), .b(new_n278), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  nor043aa1d12x5               g194(.a(new_n228), .b(new_n269), .c(new_n289), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n202), .c(new_n120), .d(new_n200), .o1(new_n291));
  oao003aa1n02x5               g196(.a(\a[26] ), .b(\b[25] ), .c(new_n281), .carry(new_n292));
  aobi12aa1n06x5               g197(.a(new_n292), .b(new_n276), .c(new_n288), .out0(new_n293));
  xorc02aa1n12x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(new_n291), .out0(\s[27] ));
  nor042aa1n03x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  inv040aa1n03x5               g201(.a(new_n296), .o1(new_n297));
  aobi12aa1n02x7               g202(.a(new_n294), .b(new_n293), .c(new_n291), .out0(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[27] ), .b(\a[28] ), .out0(new_n299));
  nano22aa1n03x5               g204(.a(new_n298), .b(new_n297), .c(new_n299), .out0(new_n300));
  nand22aa1n03x5               g205(.a(new_n244), .b(new_n241), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[23] ), .b(\b[22] ), .out0(new_n302));
  xorc02aa1n02x5               g207(.a(\a[24] ), .b(\b[23] ), .out0(new_n303));
  nano22aa1n03x7               g208(.a(new_n301), .b(new_n302), .c(new_n303), .out0(new_n304));
  oai012aa1n04x7               g209(.a(new_n304), .b(new_n254), .c(new_n230), .o1(new_n305));
  aoai13aa1n06x5               g210(.a(new_n292), .b(new_n289), .c(new_n305), .d(new_n275), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n294), .b(new_n306), .c(new_n198), .d(new_n290), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n299), .b(new_n307), .c(new_n297), .o1(new_n308));
  norp02aa1n03x5               g213(.a(new_n308), .b(new_n300), .o1(\s[28] ));
  norb02aa1n02x5               g214(.a(new_n294), .b(new_n299), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n198), .d(new_n290), .o1(new_n311));
  oao003aa1n03x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n297), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[28] ), .b(\a[29] ), .out0(new_n313));
  tech160nm_fiaoi012aa1n02p5x5 g218(.a(new_n313), .b(new_n311), .c(new_n312), .o1(new_n314));
  aobi12aa1n02x7               g219(.a(new_n310), .b(new_n293), .c(new_n291), .out0(new_n315));
  nano22aa1n03x5               g220(.a(new_n315), .b(new_n312), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[29] ));
  xnrb03aa1n02x5               g222(.a(new_n110), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g223(.a(new_n294), .b(new_n313), .c(new_n299), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n306), .c(new_n198), .d(new_n290), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .carry(new_n321));
  xnrc02aa1n02x5               g226(.a(\b[29] ), .b(\a[30] ), .out0(new_n322));
  tech160nm_fiaoi012aa1n02p5x5 g227(.a(new_n322), .b(new_n320), .c(new_n321), .o1(new_n323));
  aobi12aa1n02x7               g228(.a(new_n319), .b(new_n293), .c(new_n291), .out0(new_n324));
  nano22aa1n03x5               g229(.a(new_n324), .b(new_n321), .c(new_n322), .out0(new_n325));
  norp02aa1n03x5               g230(.a(new_n323), .b(new_n325), .o1(\s[30] ));
  xnrc02aa1n02x5               g231(.a(\b[30] ), .b(\a[31] ), .out0(new_n327));
  norb02aa1n02x5               g232(.a(new_n319), .b(new_n322), .out0(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n306), .c(new_n198), .d(new_n290), .o1(new_n329));
  oao003aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n330));
  tech160nm_fiaoi012aa1n02p5x5 g235(.a(new_n327), .b(new_n329), .c(new_n330), .o1(new_n331));
  aobi12aa1n02x7               g236(.a(new_n328), .b(new_n293), .c(new_n291), .out0(new_n332));
  nano22aa1n03x5               g237(.a(new_n332), .b(new_n327), .c(new_n330), .out0(new_n333));
  norp02aa1n03x5               g238(.a(new_n331), .b(new_n333), .o1(\s[31] ));
  xnrb03aa1n02x5               g239(.a(new_n154), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g240(.a(new_n112), .o1(new_n336));
  aoi122aa1n02x5               g241(.a(new_n114), .b(new_n336), .c(new_n113), .d(new_n111), .e(new_n115), .o1(new_n337));
  aoi012aa1n02x5               g242(.a(new_n337), .b(new_n336), .c(new_n156), .o1(\s[4] ));
  xorb03aa1n02x5               g243(.a(new_n156), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  xorc02aa1n02x5               g244(.a(\a[5] ), .b(\b[4] ), .out0(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n118), .c(new_n116), .d(new_n111), .o1(new_n341));
  oai012aa1n02x5               g246(.a(new_n341), .b(\b[4] ), .c(\a[5] ), .o1(new_n342));
  xorb03aa1n02x5               g247(.a(new_n342), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi022aa1n02x5               g248(.a(new_n341), .b(new_n99), .c(\a[6] ), .d(\b[5] ), .o1(new_n344));
  xorb03aa1n02x5               g249(.a(new_n344), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g250(.a(new_n100), .b(new_n101), .c(new_n344), .o1(new_n346));
  xnrb03aa1n02x5               g251(.a(new_n346), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g252(.a(new_n120), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


