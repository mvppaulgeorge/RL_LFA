// Benchmark "adder" written by ABC on Wed Jul 17 19:34:24 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n329, new_n330, new_n332,
    new_n333, new_n335, new_n336, new_n337, new_n338, new_n340, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  orn002aa1n02x5               g004(.a(\a[2] ), .b(\b[1] ), .o(new_n100));
  nanp02aa1n04x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n06x5               g006(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(new_n102));
  xnrc02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .out0(new_n103));
  inv000aa1d42x5               g008(.a(\a[3] ), .o1(new_n104));
  inv000aa1d42x5               g009(.a(\b[2] ), .o1(new_n105));
  and002aa1n24x5               g010(.a(\b[3] ), .b(\a[4] ), .o(new_n106));
  nor002aa1n03x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  aoi112aa1n06x5               g012(.a(new_n106), .b(new_n107), .c(new_n104), .d(new_n105), .o1(new_n108));
  aoai13aa1n06x5               g013(.a(new_n108), .b(new_n103), .c(new_n100), .d(new_n102), .o1(new_n109));
  norp02aa1n04x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  norp02aa1n04x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nand42aa1n06x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nona22aa1n09x5               g017(.a(new_n112), .b(new_n111), .c(new_n110), .out0(new_n113));
  nor042aa1d18x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  oab012aa1n04x5               g019(.a(new_n114), .b(\a[8] ), .c(\b[7] ), .out0(new_n115));
  aoi022aa1n09x5               g020(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n116));
  aoi022aa1n06x5               g021(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n117));
  nano32aa1n03x7               g022(.a(new_n113), .b(new_n117), .c(new_n115), .d(new_n116), .out0(new_n118));
  nand42aa1n06x5               g023(.a(new_n118), .b(new_n109), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n114), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  and002aa1n03x5               g026(.a(\b[6] ), .b(\a[7] ), .o(new_n122));
  aoi112aa1n06x5               g027(.a(new_n122), .b(new_n114), .c(\a[6] ), .d(\b[5] ), .o1(new_n123));
  xorc02aa1n12x5               g028(.a(\a[8] ), .b(\b[7] ), .out0(new_n124));
  aoi013aa1n09x5               g029(.a(new_n121), .b(new_n113), .c(new_n123), .d(new_n124), .o1(new_n125));
  xnrc02aa1n12x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n99), .b(new_n126), .c(new_n119), .d(new_n125), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n16x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand22aa1n09x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1d24x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(new_n127), .b(new_n132), .o1(new_n133));
  aoai13aa1n12x5               g038(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n134));
  nor042aa1n12x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand02aa1n03x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  inv000aa1d42x5               g043(.a(new_n135), .o1(new_n139));
  inv040aa1n02x5               g044(.a(new_n134), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n137), .b(new_n140), .c(new_n127), .d(new_n132), .o1(new_n141));
  nor042aa1n03x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1n03x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  aoi012aa1n02x5               g049(.a(new_n144), .b(new_n141), .c(new_n139), .o1(new_n145));
  aobi12aa1n02x5               g050(.a(new_n137), .b(new_n133), .c(new_n134), .out0(new_n146));
  nano22aa1n02x4               g051(.a(new_n146), .b(new_n139), .c(new_n144), .out0(new_n147));
  norp02aa1n02x5               g052(.a(new_n147), .b(new_n145), .o1(\s[12] ));
  nano23aa1n06x5               g053(.a(new_n135), .b(new_n142), .c(new_n143), .d(new_n136), .out0(new_n149));
  nona22aa1n02x4               g054(.a(new_n149), .b(new_n126), .c(new_n131), .out0(new_n150));
  tech160nm_fiaoi012aa1n04x5   g055(.a(new_n142), .b(new_n135), .c(new_n143), .o1(new_n151));
  aobi12aa1n06x5               g056(.a(new_n151), .b(new_n149), .c(new_n140), .out0(new_n152));
  aoai13aa1n03x5               g057(.a(new_n152), .b(new_n150), .c(new_n119), .d(new_n125), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n12x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n155), .b(new_n153), .c(new_n156), .o1(new_n157));
  xnrb03aa1n02x5               g062(.a(new_n157), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nanp02aa1n02x5               g063(.a(new_n102), .b(new_n100), .o1(new_n159));
  xorc02aa1n02x5               g064(.a(\a[3] ), .b(\b[2] ), .out0(new_n160));
  aobi12aa1n06x5               g065(.a(new_n108), .b(new_n160), .c(new_n159), .out0(new_n161));
  norb03aa1n03x5               g066(.a(new_n112), .b(new_n110), .c(new_n111), .out0(new_n162));
  nanp02aa1n02x5               g067(.a(new_n117), .b(new_n116), .o1(new_n163));
  nanb03aa1n09x5               g068(.a(new_n163), .b(new_n162), .c(new_n115), .out0(new_n164));
  oai012aa1d24x5               g069(.a(new_n125), .b(new_n161), .c(new_n164), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n143), .b(new_n136), .c(new_n135), .d(new_n142), .out0(new_n166));
  nor043aa1n02x5               g071(.a(new_n166), .b(new_n131), .c(new_n126), .o1(new_n167));
  oai012aa1n02x7               g072(.a(new_n151), .b(new_n166), .c(new_n134), .o1(new_n168));
  nor042aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand42aa1n06x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nona23aa1n09x5               g075(.a(new_n170), .b(new_n156), .c(new_n155), .d(new_n169), .out0(new_n171));
  inv040aa1n06x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n165), .d(new_n167), .o1(new_n173));
  oa0012aa1n06x5               g078(.a(new_n170), .b(new_n169), .c(new_n155), .o(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  orn002aa1n24x5               g080(.a(\a[15] ), .b(\b[14] ), .o(new_n176));
  nand02aa1d28x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand02aa1d16x5               g082(.a(new_n176), .b(new_n177), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n173), .c(new_n175), .out0(\s[15] ));
  aoai13aa1n02x5               g085(.a(new_n179), .b(new_n174), .c(new_n153), .d(new_n172), .o1(new_n181));
  xnrc02aa1n12x5               g086(.a(\b[15] ), .b(\a[16] ), .out0(new_n182));
  tech160nm_fiaoi012aa1n02p5x5 g087(.a(new_n182), .b(new_n181), .c(new_n176), .o1(new_n183));
  tech160nm_fiaoi012aa1n02p5x5 g088(.a(new_n178), .b(new_n173), .c(new_n175), .o1(new_n184));
  nano22aa1n02x4               g089(.a(new_n184), .b(new_n176), .c(new_n182), .out0(new_n185));
  norp02aa1n02x5               g090(.a(new_n185), .b(new_n183), .o1(\s[16] ));
  nor043aa1n02x5               g091(.a(new_n171), .b(new_n178), .c(new_n182), .o1(new_n187));
  nand02aa1n02x5               g092(.a(new_n187), .b(new_n167), .o1(new_n188));
  orn002aa1n02x5               g093(.a(\a[16] ), .b(\b[15] ), .o(new_n189));
  and002aa1n02x5               g094(.a(\b[15] ), .b(\a[16] ), .o(new_n190));
  oai112aa1n02x7               g095(.a(new_n170), .b(new_n177), .c(new_n169), .d(new_n155), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n189), .b(new_n190), .c(new_n191), .d(new_n176), .o1(new_n192));
  aoi012aa1n06x5               g097(.a(new_n192), .b(new_n168), .c(new_n187), .o1(new_n193));
  aoai13aa1n12x5               g098(.a(new_n193), .b(new_n188), .c(new_n119), .d(new_n125), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g100(.a(\a[18] ), .o1(new_n196));
  inv040aa1d32x5               g101(.a(\a[17] ), .o1(new_n197));
  inv040aa1d28x5               g102(.a(\b[16] ), .o1(new_n198));
  oaoi03aa1n03x5               g103(.a(new_n197), .b(new_n198), .c(new_n194), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[17] ), .c(new_n196), .out0(\s[18] ));
  nona22aa1n09x5               g105(.a(new_n172), .b(new_n178), .c(new_n182), .out0(new_n201));
  nor042aa1n06x5               g106(.a(new_n201), .b(new_n150), .o1(new_n202));
  oabi12aa1n18x5               g107(.a(new_n192), .b(new_n201), .c(new_n152), .out0(new_n203));
  xroi22aa1d04x5               g108(.a(new_n197), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n203), .c(new_n165), .d(new_n202), .o1(new_n205));
  nand02aa1d16x5               g110(.a(new_n198), .b(new_n197), .o1(new_n206));
  oaoi03aa1n12x5               g111(.a(\a[18] ), .b(\b[17] ), .c(new_n206), .o1(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  nor002aa1d32x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand42aa1n06x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nanb02aa1n02x5               g115(.a(new_n209), .b(new_n210), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n205), .c(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n03x5               g119(.a(new_n209), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n212), .b(new_n207), .c(new_n194), .d(new_n204), .o1(new_n216));
  nor042aa1n03x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand42aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoi012aa1n03x5               g124(.a(new_n219), .b(new_n216), .c(new_n215), .o1(new_n220));
  tech160nm_fiaoi012aa1n05x5   g125(.a(new_n211), .b(new_n205), .c(new_n208), .o1(new_n221));
  nano22aa1n02x4               g126(.a(new_n221), .b(new_n215), .c(new_n219), .out0(new_n222));
  nor002aa1n02x5               g127(.a(new_n220), .b(new_n222), .o1(\s[20] ));
  nano23aa1d15x5               g128(.a(new_n209), .b(new_n217), .c(new_n218), .d(new_n210), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  norb02aa1n02x5               g130(.a(new_n204), .b(new_n225), .out0(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n203), .c(new_n165), .d(new_n202), .o1(new_n227));
  tech160nm_fioaoi03aa1n04x5   g132(.a(\a[20] ), .b(\b[19] ), .c(new_n215), .o1(new_n228));
  aoi012aa1d24x5               g133(.a(new_n228), .b(new_n224), .c(new_n207), .o1(new_n229));
  nor042aa1n06x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand42aa1n03x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  nanb02aa1n02x5               g136(.a(new_n230), .b(new_n231), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n227), .c(new_n229), .out0(\s[21] ));
  inv000aa1d42x5               g139(.a(new_n230), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n229), .o1(new_n236));
  aoai13aa1n03x5               g141(.a(new_n233), .b(new_n236), .c(new_n194), .d(new_n226), .o1(new_n237));
  nor002aa1n03x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nand02aa1n04x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nanb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(new_n240));
  aoi012aa1n03x5               g145(.a(new_n240), .b(new_n237), .c(new_n235), .o1(new_n241));
  aoi012aa1n03x5               g146(.a(new_n232), .b(new_n227), .c(new_n229), .o1(new_n242));
  nano22aa1n03x5               g147(.a(new_n242), .b(new_n235), .c(new_n240), .out0(new_n243));
  norp02aa1n03x5               g148(.a(new_n241), .b(new_n243), .o1(\s[22] ));
  nano23aa1n03x7               g149(.a(new_n230), .b(new_n238), .c(new_n239), .d(new_n231), .out0(new_n245));
  and003aa1n02x5               g150(.a(new_n204), .b(new_n245), .c(new_n224), .o(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n203), .c(new_n165), .d(new_n202), .o1(new_n247));
  nona23aa1n09x5               g152(.a(new_n239), .b(new_n231), .c(new_n230), .d(new_n238), .out0(new_n248));
  oaoi03aa1n02x5               g153(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .o1(new_n249));
  oab012aa1n06x5               g154(.a(new_n249), .b(new_n229), .c(new_n248), .out0(new_n250));
  orn002aa1n24x5               g155(.a(\a[23] ), .b(\b[22] ), .o(new_n251));
  nanp02aa1n06x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  nand22aa1n09x5               g157(.a(new_n251), .b(new_n252), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n247), .c(new_n250), .out0(\s[23] ));
  inv040aa1n03x5               g160(.a(new_n250), .o1(new_n256));
  aoai13aa1n06x5               g161(.a(new_n254), .b(new_n256), .c(new_n194), .d(new_n246), .o1(new_n257));
  xnrc02aa1n02x5               g162(.a(\b[23] ), .b(\a[24] ), .out0(new_n258));
  aoi012aa1n02x7               g163(.a(new_n258), .b(new_n257), .c(new_n251), .o1(new_n259));
  aoi012aa1n03x5               g164(.a(new_n253), .b(new_n247), .c(new_n250), .o1(new_n260));
  nano22aa1n02x4               g165(.a(new_n260), .b(new_n251), .c(new_n258), .out0(new_n261));
  norp02aa1n03x5               g166(.a(new_n259), .b(new_n261), .o1(\s[24] ));
  nona22aa1n06x5               g167(.a(new_n245), .b(new_n258), .c(new_n253), .out0(new_n263));
  nano22aa1n03x7               g168(.a(new_n263), .b(new_n204), .c(new_n224), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n203), .c(new_n165), .d(new_n202), .o1(new_n265));
  norp02aa1n02x5               g170(.a(\b[23] ), .b(\a[24] ), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n252), .b(new_n238), .c(new_n230), .d(new_n239), .o1(new_n267));
  aoi022aa1n02x5               g172(.a(new_n267), .b(new_n251), .c(\a[24] ), .d(\b[23] ), .o1(new_n268));
  nor042aa1n04x5               g173(.a(new_n268), .b(new_n266), .o1(new_n269));
  oai012aa1d24x5               g174(.a(new_n269), .b(new_n229), .c(new_n263), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  xnrc02aa1n12x5               g176(.a(\b[24] ), .b(\a[25] ), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  xnbna2aa1n03x5               g178(.a(new_n273), .b(new_n265), .c(new_n271), .out0(\s[25] ));
  nor042aa1n03x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n273), .b(new_n270), .c(new_n194), .d(new_n264), .o1(new_n277));
  xnrc02aa1n12x5               g182(.a(\b[25] ), .b(\a[26] ), .out0(new_n278));
  aoi012aa1n03x5               g183(.a(new_n278), .b(new_n277), .c(new_n276), .o1(new_n279));
  aoi012aa1n02x7               g184(.a(new_n272), .b(new_n265), .c(new_n271), .o1(new_n280));
  nano22aa1n02x4               g185(.a(new_n280), .b(new_n276), .c(new_n278), .out0(new_n281));
  nor002aa1n02x5               g186(.a(new_n279), .b(new_n281), .o1(\s[26] ));
  nor042aa1n12x5               g187(.a(new_n278), .b(new_n272), .o1(new_n283));
  nano32aa1n03x7               g188(.a(new_n263), .b(new_n204), .c(new_n283), .d(new_n224), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n203), .c(new_n165), .d(new_n202), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .c(new_n276), .carry(new_n286));
  aobi12aa1n18x5               g191(.a(new_n286), .b(new_n270), .c(new_n283), .out0(new_n287));
  xorc02aa1n02x5               g192(.a(\a[27] ), .b(\b[26] ), .out0(new_n288));
  xnbna2aa1n03x5               g193(.a(new_n288), .b(new_n285), .c(new_n287), .out0(\s[27] ));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  inv040aa1n03x5               g195(.a(new_n290), .o1(new_n291));
  norp03aa1n03x5               g196(.a(new_n248), .b(new_n253), .c(new_n258), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n228), .c(new_n207), .d(new_n224), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n283), .o1(new_n294));
  aoai13aa1n04x5               g199(.a(new_n286), .b(new_n294), .c(new_n293), .d(new_n269), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n288), .b(new_n295), .c(new_n194), .d(new_n284), .o1(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[27] ), .b(\a[28] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n296), .c(new_n291), .o1(new_n298));
  aobi12aa1n02x7               g203(.a(new_n288), .b(new_n285), .c(new_n287), .out0(new_n299));
  nano22aa1n03x5               g204(.a(new_n299), .b(new_n291), .c(new_n297), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n298), .b(new_n300), .o1(\s[28] ));
  norb02aa1n02x5               g206(.a(new_n288), .b(new_n297), .out0(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n295), .c(new_n194), .d(new_n284), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n291), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[28] ), .b(\a[29] ), .out0(new_n305));
  aoi012aa1n02x5               g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  aobi12aa1n02x7               g211(.a(new_n302), .b(new_n285), .c(new_n287), .out0(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n304), .c(new_n305), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n306), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g215(.a(new_n288), .b(new_n305), .c(new_n297), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n295), .c(new_n194), .d(new_n284), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[29] ), .b(\a[30] ), .out0(new_n314));
  aoi012aa1n02x7               g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  aobi12aa1n03x5               g220(.a(new_n311), .b(new_n285), .c(new_n287), .out0(new_n316));
  nano22aa1n03x5               g221(.a(new_n316), .b(new_n313), .c(new_n314), .out0(new_n317));
  norp02aa1n03x5               g222(.a(new_n315), .b(new_n317), .o1(\s[30] ));
  xnrc02aa1n02x5               g223(.a(\b[30] ), .b(\a[31] ), .out0(new_n319));
  nona32aa1n02x4               g224(.a(new_n288), .b(new_n314), .c(new_n305), .d(new_n297), .out0(new_n320));
  inv000aa1d42x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n295), .c(new_n194), .d(new_n284), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n323));
  aoi012aa1n03x5               g228(.a(new_n319), .b(new_n322), .c(new_n323), .o1(new_n324));
  tech160nm_fiaoi012aa1n05x5   g229(.a(new_n320), .b(new_n285), .c(new_n287), .o1(new_n325));
  nano22aa1n03x5               g230(.a(new_n325), .b(new_n319), .c(new_n323), .out0(new_n326));
  norp02aa1n03x5               g231(.a(new_n324), .b(new_n326), .o1(\s[31] ));
  xnbna2aa1n03x5               g232(.a(new_n160), .b(new_n100), .c(new_n102), .out0(\s[3] ));
  norp02aa1n02x5               g233(.a(new_n106), .b(new_n107), .o1(new_n329));
  oaoi03aa1n02x5               g234(.a(new_n104), .b(new_n105), .c(new_n159), .o1(new_n330));
  oai012aa1n02x5               g235(.a(new_n109), .b(new_n330), .c(new_n329), .o1(\s[4] ));
  inv000aa1d42x5               g236(.a(new_n106), .o1(new_n332));
  xnrc02aa1n02x5               g237(.a(\b[4] ), .b(\a[5] ), .out0(new_n333));
  xnbna2aa1n03x5               g238(.a(new_n333), .b(new_n109), .c(new_n332), .out0(\s[5] ));
  norb02aa1n02x5               g239(.a(new_n112), .b(new_n111), .out0(new_n335));
  nona22aa1n02x4               g240(.a(new_n109), .b(new_n333), .c(new_n106), .out0(new_n336));
  norb02aa1n02x5               g241(.a(new_n336), .b(new_n110), .out0(new_n337));
  nanp02aa1n02x5               g242(.a(new_n336), .b(new_n162), .o1(new_n338));
  oai012aa1n02x5               g243(.a(new_n338), .b(new_n337), .c(new_n335), .o1(\s[6] ));
  norp02aa1n02x5               g244(.a(new_n122), .b(new_n114), .o1(new_n340));
  xobna2aa1n03x5               g245(.a(new_n340), .b(new_n338), .c(new_n112), .out0(\s[7] ));
  nanp02aa1n02x5               g246(.a(new_n338), .b(new_n123), .o1(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n124), .b(new_n342), .c(new_n120), .out0(\s[8] ));
  xobna2aa1n03x5               g248(.a(new_n126), .b(new_n119), .c(new_n125), .out0(\s[9] ));
endmodule


