// Benchmark "adder" written by ABC on Wed Jul 17 16:54:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n329, new_n331, new_n333,
    new_n335, new_n336, new_n339;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1d06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n12x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n09x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor002aa1d32x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1d32x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n06x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  inv000aa1d42x5               g012(.a(\a[3] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[2] ), .o1(new_n109));
  aoai13aa1n06x5               g014(.a(new_n104), .b(new_n103), .c(new_n108), .d(new_n109), .o1(new_n110));
  oai012aa1n12x5               g015(.a(new_n110), .b(new_n107), .c(new_n102), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n24x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  norp02aa1n09x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nona23aa1n02x5               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  nanp02aa1n12x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1n06x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanb02aa1n12x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  xorc02aa1n12x5               g024(.a(\a[5] ), .b(\b[4] ), .out0(new_n120));
  norb03aa1n09x5               g025(.a(new_n120), .b(new_n116), .c(new_n119), .out0(new_n121));
  inv000aa1d42x5               g026(.a(new_n112), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n113), .o1(new_n123));
  inv000aa1n02x5               g028(.a(new_n114), .o1(new_n124));
  nor042aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  aoai13aa1n04x5               g030(.a(new_n115), .b(new_n118), .c(new_n125), .d(new_n117), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n122), .b(new_n123), .c(new_n126), .d(new_n124), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n121), .d(new_n111), .o1(new_n129));
  xobna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  nand42aa1n04x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor002aa1d32x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nanb02aa1n12x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  oai022aa1d24x5               g038(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n134), .b(new_n129), .out0(new_n135));
  aob012aa1n02x5               g040(.a(new_n135), .b(\b[9] ), .c(\a[10] ), .out0(new_n136));
  inv040aa1n09x5               g041(.a(new_n132), .o1(new_n137));
  aoi022aa1d24x5               g042(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n138));
  nand42aa1n16x5               g043(.a(new_n138), .b(new_n137), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  aoi022aa1n02x5               g045(.a(new_n136), .b(new_n133), .c(new_n135), .d(new_n140), .o1(\s[11] ));
  inv000aa1n03x5               g046(.a(new_n102), .o1(new_n142));
  nano23aa1n06x5               g047(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n143));
  aobi12aa1n06x5               g048(.a(new_n110), .b(new_n143), .c(new_n142), .out0(new_n144));
  nanb02aa1n03x5               g049(.a(new_n112), .b(new_n113), .out0(new_n145));
  norb02aa1n02x7               g050(.a(new_n115), .b(new_n114), .out0(new_n146));
  nona23aa1n03x5               g051(.a(new_n120), .b(new_n146), .c(new_n145), .d(new_n119), .out0(new_n147));
  nand42aa1n02x5               g052(.a(new_n126), .b(new_n124), .o1(new_n148));
  tech160nm_fiaoi012aa1n03p5x5 g053(.a(new_n112), .b(new_n148), .c(new_n113), .o1(new_n149));
  tech160nm_fioai012aa1n05x5   g054(.a(new_n149), .b(new_n144), .c(new_n147), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n140), .b(new_n134), .c(new_n150), .d(new_n128), .o1(new_n151));
  nor042aa1n04x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  nand02aa1n04x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  norb02aa1n06x5               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  xnbna2aa1n03x5               g059(.a(new_n154), .b(new_n151), .c(new_n137), .out0(\s[12] ));
  nona23aa1d24x5               g060(.a(new_n154), .b(new_n128), .c(new_n97), .d(new_n133), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n03x5               g062(.a(new_n157), .b(new_n127), .c(new_n121), .d(new_n111), .o1(new_n158));
  oaoi03aa1n12x5               g063(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .o1(new_n159));
  nanb03aa1n09x5               g064(.a(new_n152), .b(new_n134), .c(new_n153), .out0(new_n160));
  oabi12aa1n18x5               g065(.a(new_n159), .b(new_n160), .c(new_n139), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nanp02aa1n03x5               g067(.a(new_n158), .b(new_n162), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1d18x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand22aa1n09x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n165), .b(new_n163), .c(new_n166), .o1(new_n167));
  xnrb03aa1n03x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1d18x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1d28x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nona23aa1d18x5               g075(.a(new_n170), .b(new_n166), .c(new_n165), .d(new_n169), .out0(new_n171));
  inv000aa1n02x5               g076(.a(new_n171), .o1(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n161), .c(new_n150), .d(new_n157), .o1(new_n173));
  aoi012aa1n02x5               g078(.a(new_n169), .b(new_n165), .c(new_n170), .o1(new_n174));
  nor042aa1n04x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nand02aa1n06x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  xobna2aa1n03x5               g082(.a(new_n177), .b(new_n173), .c(new_n174), .out0(\s[15] ));
  aoai13aa1n04x5               g083(.a(new_n174), .b(new_n171), .c(new_n158), .d(new_n162), .o1(new_n179));
  nor042aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanp02aa1n02x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nanb02aa1n03x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n175), .c(new_n179), .d(new_n176), .o1(new_n183));
  aoi112aa1n03x5               g088(.a(new_n175), .b(new_n182), .c(new_n179), .d(new_n176), .o1(new_n184));
  nanb02aa1n03x5               g089(.a(new_n184), .b(new_n183), .out0(\s[16] ));
  nano23aa1n03x7               g090(.a(new_n175), .b(new_n180), .c(new_n181), .d(new_n176), .out0(new_n186));
  nano22aa1d15x5               g091(.a(new_n156), .b(new_n172), .c(new_n186), .out0(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n127), .c(new_n111), .d(new_n121), .o1(new_n188));
  norp03aa1n06x5               g093(.a(new_n171), .b(new_n177), .c(new_n182), .o1(new_n189));
  aoai13aa1n02x5               g094(.a(new_n176), .b(new_n169), .c(new_n165), .d(new_n170), .o1(new_n190));
  aboi22aa1n03x5               g095(.a(new_n175), .b(new_n190), .c(\a[16] ), .d(\b[15] ), .out0(new_n191));
  aoi112aa1n09x5               g096(.a(new_n180), .b(new_n191), .c(new_n161), .d(new_n189), .o1(new_n192));
  nor002aa1d32x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  nand42aa1d28x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n188), .c(new_n192), .out0(\s[17] ));
  inv000aa1d42x5               g101(.a(\a[18] ), .o1(new_n197));
  nanp02aa1n06x5               g102(.a(new_n188), .b(new_n192), .o1(new_n198));
  tech160nm_fiaoi012aa1n05x5   g103(.a(new_n193), .b(new_n198), .c(new_n195), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[17] ), .c(new_n197), .out0(\s[18] ));
  nanp02aa1n03x5               g105(.a(new_n161), .b(new_n189), .o1(new_n201));
  nona22aa1n03x5               g106(.a(new_n201), .b(new_n191), .c(new_n180), .out0(new_n202));
  nor002aa1n20x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand42aa1d28x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nano23aa1d15x5               g109(.a(new_n193), .b(new_n203), .c(new_n204), .d(new_n194), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n202), .c(new_n150), .d(new_n187), .o1(new_n206));
  oa0012aa1n02x5               g111(.a(new_n204), .b(new_n203), .c(new_n193), .o(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  nor042aa1d18x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand22aa1n04x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  norb02aa1n09x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n206), .c(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g118(.a(new_n206), .b(new_n208), .o1(new_n214));
  nor042aa1d18x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nand02aa1d28x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nanb02aa1n03x5               g121(.a(new_n215), .b(new_n216), .out0(new_n217));
  aoai13aa1n02x5               g122(.a(new_n217), .b(new_n209), .c(new_n214), .d(new_n210), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n211), .b(new_n207), .c(new_n198), .d(new_n205), .o1(new_n219));
  nona22aa1n02x5               g124(.a(new_n219), .b(new_n217), .c(new_n209), .out0(new_n220));
  nanp02aa1n03x5               g125(.a(new_n218), .b(new_n220), .o1(\s[20] ));
  nanb03aa1d18x5               g126(.a(new_n217), .b(new_n205), .c(new_n211), .out0(new_n222));
  nanb03aa1n06x5               g127(.a(new_n215), .b(new_n216), .c(new_n210), .out0(new_n223));
  orn002aa1n03x5               g128(.a(\a[19] ), .b(\b[18] ), .o(new_n224));
  oai112aa1n06x5               g129(.a(new_n224), .b(new_n204), .c(new_n203), .d(new_n193), .o1(new_n225));
  aoi012aa1n12x5               g130(.a(new_n215), .b(new_n209), .c(new_n216), .o1(new_n226));
  oai012aa1n18x5               g131(.a(new_n226), .b(new_n225), .c(new_n223), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n04x5               g133(.a(new_n228), .b(new_n222), .c(new_n188), .d(new_n192), .o1(new_n229));
  nor002aa1n20x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand42aa1n16x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n222), .o1(new_n233));
  aoi112aa1n03x4               g138(.a(new_n232), .b(new_n227), .c(new_n198), .d(new_n233), .o1(new_n234));
  aoi012aa1n03x5               g139(.a(new_n234), .b(new_n229), .c(new_n232), .o1(\s[21] ));
  nor002aa1n06x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  nand42aa1n16x5               g141(.a(\b[21] ), .b(\a[22] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n239), .b(new_n230), .c(new_n229), .d(new_n232), .o1(new_n240));
  nand02aa1n02x5               g145(.a(new_n229), .b(new_n232), .o1(new_n241));
  nona22aa1n02x5               g146(.a(new_n241), .b(new_n239), .c(new_n230), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n242), .b(new_n240), .o1(\s[22] ));
  nano23aa1n09x5               g148(.a(new_n230), .b(new_n236), .c(new_n237), .d(new_n231), .out0(new_n244));
  nanb02aa1n03x5               g149(.a(new_n222), .b(new_n244), .out0(new_n245));
  nano22aa1n03x7               g150(.a(new_n215), .b(new_n210), .c(new_n216), .out0(new_n246));
  tech160nm_fioai012aa1n03p5x5 g151(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .o1(new_n247));
  oab012aa1n06x5               g152(.a(new_n247), .b(new_n193), .c(new_n203), .out0(new_n248));
  inv000aa1n06x5               g153(.a(new_n226), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n244), .b(new_n249), .c(new_n248), .d(new_n246), .o1(new_n250));
  oa0012aa1n02x5               g155(.a(new_n237), .b(new_n236), .c(new_n230), .o(new_n251));
  inv000aa1n03x5               g156(.a(new_n251), .o1(new_n252));
  nanp02aa1n02x5               g157(.a(new_n250), .b(new_n252), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n245), .c(new_n188), .d(new_n192), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[23] ), .b(\b[22] ), .out0(new_n258));
  tech160nm_fixnrc02aa1n05x5   g163(.a(\b[23] ), .b(\a[24] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n260));
  nand02aa1n02x5               g165(.a(new_n255), .b(new_n258), .o1(new_n261));
  nona22aa1n02x5               g166(.a(new_n261), .b(new_n259), .c(new_n257), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n262), .b(new_n260), .o1(\s[24] ));
  norb02aa1n06x4               g168(.a(new_n258), .b(new_n259), .out0(new_n264));
  nanb03aa1n03x5               g169(.a(new_n222), .b(new_n264), .c(new_n244), .out0(new_n265));
  inv030aa1n02x5               g170(.a(new_n264), .o1(new_n266));
  orn002aa1n02x5               g171(.a(\a[23] ), .b(\b[22] ), .o(new_n267));
  oao003aa1n02x5               g172(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .carry(new_n268));
  aoai13aa1n12x5               g173(.a(new_n268), .b(new_n266), .c(new_n250), .d(new_n252), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n265), .c(new_n188), .d(new_n192), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n276));
  nand02aa1n02x5               g181(.a(new_n271), .b(new_n274), .o1(new_n277));
  nona22aa1n02x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .out0(new_n278));
  nand42aa1n02x5               g183(.a(new_n278), .b(new_n276), .o1(\s[26] ));
  norb02aa1n06x4               g184(.a(new_n274), .b(new_n275), .out0(new_n280));
  inv030aa1n02x5               g185(.a(new_n280), .o1(new_n281));
  nano23aa1n06x5               g186(.a(new_n281), .b(new_n222), .c(new_n264), .d(new_n244), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n202), .c(new_n150), .d(new_n187), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(\b[25] ), .b(\a[26] ), .o1(new_n284));
  oai022aa1n02x5               g189(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n285));
  aoi022aa1n12x5               g190(.a(new_n269), .b(new_n280), .c(new_n284), .d(new_n285), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[27] ), .b(\b[26] ), .out0(new_n287));
  xnbna2aa1n03x5               g192(.a(new_n287), .b(new_n286), .c(new_n283), .out0(\s[27] ));
  nand42aa1n03x5               g193(.a(new_n286), .b(new_n283), .o1(new_n289));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  xnrc02aa1n12x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n289), .d(new_n287), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n264), .b(new_n251), .c(new_n227), .d(new_n244), .o1(new_n293));
  nanp02aa1n02x5               g198(.a(new_n285), .b(new_n284), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n281), .c(new_n293), .d(new_n268), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n287), .b(new_n295), .c(new_n198), .d(new_n282), .o1(new_n296));
  nona22aa1n02x5               g201(.a(new_n296), .b(new_n291), .c(new_n290), .out0(new_n297));
  nanp02aa1n03x5               g202(.a(new_n292), .b(new_n297), .o1(\s[28] ));
  norb02aa1n03x5               g203(.a(new_n287), .b(new_n291), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n295), .c(new_n198), .d(new_n282), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n299), .o1(new_n301));
  orn002aa1n02x5               g206(.a(\a[27] ), .b(\b[26] ), .o(new_n302));
  oao003aa1n03x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n302), .carry(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n301), .c(new_n286), .d(new_n283), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n303), .b(new_n305), .out0(new_n306));
  aoi022aa1n03x5               g211(.a(new_n304), .b(new_n305), .c(new_n300), .d(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d18x5               g213(.a(new_n291), .b(new_n287), .c(new_n305), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n295), .c(new_n198), .d(new_n282), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n309), .o1(new_n311));
  oaoi03aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .o1(new_n312));
  inv000aa1n03x5               g217(.a(new_n312), .o1(new_n313));
  aoai13aa1n02x7               g218(.a(new_n313), .b(new_n311), .c(new_n286), .d(new_n283), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .out0(new_n315));
  and002aa1n02x5               g220(.a(\b[28] ), .b(\a[29] ), .o(new_n316));
  oabi12aa1n02x5               g221(.a(new_n315), .b(\a[29] ), .c(\b[28] ), .out0(new_n317));
  oab012aa1n02x4               g222(.a(new_n317), .b(new_n303), .c(new_n316), .out0(new_n318));
  aoi022aa1n03x5               g223(.a(new_n314), .b(new_n315), .c(new_n310), .d(new_n318), .o1(\s[30] ));
  nand03aa1n02x5               g224(.a(new_n299), .b(new_n305), .c(new_n315), .o1(new_n320));
  nanb02aa1n02x5               g225(.a(new_n320), .b(new_n289), .out0(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  aoai13aa1n02x7               g229(.a(new_n323), .b(new_n320), .c(new_n286), .d(new_n283), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n321), .b(new_n324), .c(new_n325), .d(new_n322), .o1(\s[31] ));
  xorb03aa1n02x5               g231(.a(new_n102), .b(\b[2] ), .c(new_n108), .out0(\s[3] ));
  norb02aa1n02x5               g232(.a(new_n104), .b(new_n103), .out0(new_n328));
  aoi112aa1n02x5               g233(.a(new_n105), .b(new_n328), .c(new_n142), .d(new_n106), .o1(new_n329));
  aoib12aa1n02x5               g234(.a(new_n329), .b(new_n111), .c(new_n103), .out0(\s[4] ));
  nanp02aa1n02x5               g235(.a(new_n143), .b(new_n142), .o1(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n120), .b(new_n331), .c(new_n110), .out0(\s[5] ));
  oaoi03aa1n02x5               g237(.a(\a[5] ), .b(\b[4] ), .c(new_n144), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g239(.a(new_n146), .b(new_n118), .c(new_n333), .d(new_n117), .o1(new_n335));
  aoi112aa1n02x5               g240(.a(new_n118), .b(new_n146), .c(new_n333), .d(new_n117), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n335), .b(new_n336), .out0(\s[7] ));
  xobna2aa1n03x5               g242(.a(new_n145), .b(new_n335), .c(new_n124), .out0(\s[8] ));
  aoi112aa1n02x5               g243(.a(new_n127), .b(new_n128), .c(new_n121), .d(new_n111), .o1(new_n339));
  aoi012aa1n02x5               g244(.a(new_n339), .b(new_n150), .c(new_n128), .o1(\s[9] ));
endmodule


