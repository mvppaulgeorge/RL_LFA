// Benchmark "adder" written by ABC on Thu Jul 18 03:42:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n316, new_n317,
    new_n319, new_n320, new_n322, new_n324, new_n325, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  inv000aa1d42x5               g002(.a(\a[3] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[4] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[2] ), .o1(new_n100));
  aboi22aa1n09x5               g005(.a(\b[3] ), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n101));
  tech160nm_fixnrc02aa1n04x5   g006(.a(\b[2] ), .b(\a[3] ), .out0(new_n102));
  nanp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n04x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  oai012aa1n04x7               g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n101), .b(new_n102), .c(new_n106), .o1(new_n107));
  nor042aa1d18x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(new_n108), .o1(new_n109));
  nand02aa1n03x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  oai112aa1n02x5               g015(.a(new_n109), .b(new_n110), .c(\b[7] ), .d(\a[8] ), .o1(new_n111));
  inv040aa1d30x5               g016(.a(\a[5] ), .o1(new_n112));
  aoi022aa1d24x5               g017(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  oaib12aa1n03x5               g018(.a(new_n113), .b(\b[4] ), .c(new_n112), .out0(new_n114));
  nand42aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  orn002aa1n02x7               g020(.a(\a[7] ), .b(\b[6] ), .o(new_n116));
  nand02aa1d08x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nand23aa1n03x5               g022(.a(new_n116), .b(new_n115), .c(new_n117), .o1(new_n118));
  nor043aa1n03x5               g023(.a(new_n111), .b(new_n118), .c(new_n114), .o1(new_n119));
  nand02aa1n04x5               g024(.a(new_n119), .b(new_n107), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\a[8] ), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\b[7] ), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n117), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[4] ), .o1(new_n125));
  aoai13aa1n06x5               g030(.a(new_n110), .b(new_n108), .c(new_n112), .d(new_n125), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n123), .b(new_n124), .c(new_n126), .d(new_n116), .o1(new_n127));
  nand42aa1n02x5               g032(.a(new_n127), .b(new_n115), .o1(new_n128));
  xnrc02aa1n12x5               g033(.a(\b[8] ), .b(\a[9] ), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n97), .b(new_n129), .c(new_n128), .d(new_n120), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  aoi022aa1n09x5               g036(.a(new_n127), .b(new_n115), .c(new_n119), .d(new_n107), .o1(new_n132));
  tech160nm_fixnrc02aa1n04x5   g037(.a(\b[9] ), .b(\a[10] ), .out0(new_n133));
  oaoi13aa1n06x5               g038(.a(new_n133), .b(new_n97), .c(new_n132), .d(new_n129), .o1(new_n134));
  oaoi03aa1n12x5               g039(.a(\a[10] ), .b(\b[9] ), .c(new_n97), .o1(new_n135));
  nor002aa1n16x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand42aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  tech160nm_fioai012aa1n05x5   g043(.a(new_n138), .b(new_n134), .c(new_n135), .o1(new_n139));
  norp03aa1n02x5               g044(.a(new_n134), .b(new_n135), .c(new_n138), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(\s[11] ));
  oai012aa1n02x5               g046(.a(new_n139), .b(\b[10] ), .c(\a[11] ), .o1(new_n142));
  nor022aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1d06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  aoib12aa1n02x5               g050(.a(new_n136), .b(new_n144), .c(new_n143), .out0(new_n146));
  aoi022aa1n02x5               g051(.a(new_n142), .b(new_n145), .c(new_n139), .d(new_n146), .o1(\s[12] ));
  nona23aa1d18x5               g052(.a(new_n144), .b(new_n137), .c(new_n136), .d(new_n143), .out0(new_n148));
  nor043aa1d12x5               g053(.a(new_n148), .b(new_n133), .c(new_n129), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoi012aa1n06x5               g055(.a(new_n143), .b(new_n136), .c(new_n144), .o1(new_n151));
  oaib12aa1n06x5               g056(.a(new_n151), .b(new_n148), .c(new_n135), .out0(new_n152));
  oabi12aa1n06x5               g057(.a(new_n152), .b(new_n132), .c(new_n150), .out0(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n03x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  inv040aa1n03x5               g060(.a(new_n155), .o1(new_n156));
  tech160nm_fixnrc02aa1n02p5x5 g061(.a(\b[12] ), .b(\a[13] ), .out0(new_n157));
  nanb02aa1n02x5               g062(.a(new_n157), .b(new_n153), .out0(new_n158));
  tech160nm_fixnrc02aa1n04x5   g063(.a(\b[13] ), .b(\a[14] ), .out0(new_n159));
  xobna2aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n156), .out0(\s[14] ));
  nor042aa1n06x5               g065(.a(new_n159), .b(new_n157), .o1(new_n161));
  oaoi03aa1n02x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n162));
  xorc02aa1n02x5               g067(.a(\a[15] ), .b(\b[14] ), .out0(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n162), .c(new_n153), .d(new_n161), .o1(new_n164));
  aoi112aa1n02x5               g069(.a(new_n163), .b(new_n162), .c(new_n153), .d(new_n161), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(\s[15] ));
  inv000aa1d42x5               g071(.a(\a[15] ), .o1(new_n167));
  oaib12aa1n02x5               g072(.a(new_n164), .b(\b[14] ), .c(new_n167), .out0(new_n168));
  xorc02aa1n02x5               g073(.a(\a[16] ), .b(\b[15] ), .out0(new_n169));
  aoib12aa1n02x5               g074(.a(new_n169), .b(new_n167), .c(\b[14] ), .out0(new_n170));
  aoi022aa1n02x5               g075(.a(new_n168), .b(new_n169), .c(new_n164), .d(new_n170), .o1(\s[16] ));
  inv040aa1d32x5               g076(.a(\a[16] ), .o1(new_n172));
  xroi22aa1d06x4               g077(.a(new_n167), .b(\b[14] ), .c(new_n172), .d(\b[15] ), .out0(new_n173));
  nand23aa1n09x5               g078(.a(new_n149), .b(new_n161), .c(new_n173), .o1(new_n174));
  aoai13aa1n04x5               g079(.a(new_n173), .b(new_n162), .c(new_n152), .d(new_n161), .o1(new_n175));
  aoi112aa1n02x5               g080(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n176));
  aoib12aa1n02x5               g081(.a(new_n176), .b(new_n172), .c(\b[15] ), .out0(new_n177));
  oai112aa1n06x5               g082(.a(new_n175), .b(new_n177), .c(new_n174), .d(new_n132), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g084(.a(\a[17] ), .o1(new_n180));
  nanb02aa1n12x5               g085(.a(\b[16] ), .b(new_n180), .out0(new_n181));
  aoi012aa1n12x5               g086(.a(new_n174), .b(new_n128), .c(new_n120), .o1(new_n182));
  inv030aa1n02x5               g087(.a(new_n162), .o1(new_n183));
  inv000aa1n02x5               g088(.a(new_n173), .o1(new_n184));
  nano23aa1n09x5               g089(.a(new_n136), .b(new_n143), .c(new_n144), .d(new_n137), .out0(new_n185));
  inv030aa1n02x5               g090(.a(new_n151), .o1(new_n186));
  aoai13aa1n06x5               g091(.a(new_n161), .b(new_n186), .c(new_n185), .d(new_n135), .o1(new_n187));
  aoai13aa1n09x5               g092(.a(new_n177), .b(new_n184), .c(new_n187), .d(new_n183), .o1(new_n188));
  tech160nm_fixorc02aa1n05x5   g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  oai012aa1n03x5               g094(.a(new_n189), .b(new_n188), .c(new_n182), .o1(new_n190));
  xorc02aa1n12x5               g095(.a(\a[18] ), .b(\b[17] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n190), .c(new_n181), .out0(\s[18] ));
  inv000aa1d42x5               g097(.a(\a[18] ), .o1(new_n193));
  xroi22aa1d04x5               g098(.a(new_n180), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n194));
  oai012aa1n06x5               g099(.a(new_n194), .b(new_n188), .c(new_n182), .o1(new_n195));
  oai022aa1n04x5               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oaib12aa1n09x5               g101(.a(new_n196), .b(new_n193), .c(\b[17] ), .out0(new_n197));
  nor002aa1d32x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand42aa1n20x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n12x5               g108(.a(\a[18] ), .b(\b[17] ), .c(new_n181), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n201), .b(new_n204), .c(new_n178), .d(new_n194), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n198), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n206), .b(new_n200), .c(new_n195), .d(new_n197), .o1(new_n207));
  nor042aa1n06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand42aa1d28x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoib12aa1n02x5               g115(.a(new_n198), .b(new_n209), .c(new_n208), .out0(new_n211));
  aoi022aa1n03x5               g116(.a(new_n207), .b(new_n210), .c(new_n205), .d(new_n211), .o1(\s[20] ));
  nano23aa1n09x5               g117(.a(new_n198), .b(new_n208), .c(new_n209), .d(new_n199), .out0(new_n213));
  nand23aa1n06x5               g118(.a(new_n213), .b(new_n189), .c(new_n191), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  tech160nm_fioai012aa1n05x5   g120(.a(new_n215), .b(new_n188), .c(new_n182), .o1(new_n216));
  nona23aa1d18x5               g121(.a(new_n209), .b(new_n199), .c(new_n198), .d(new_n208), .out0(new_n217));
  aoi012aa1d18x5               g122(.a(new_n208), .b(new_n198), .c(new_n209), .o1(new_n218));
  oai012aa1d24x5               g123(.a(new_n218), .b(new_n217), .c(new_n197), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  xorc02aa1n02x5               g125(.a(\a[21] ), .b(\b[20] ), .out0(new_n221));
  xnbna2aa1n03x5               g126(.a(new_n221), .b(new_n216), .c(new_n220), .out0(\s[21] ));
  aoai13aa1n03x5               g127(.a(new_n221), .b(new_n219), .c(new_n178), .d(new_n215), .o1(new_n223));
  nor042aa1d18x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n221), .o1(new_n226));
  aoai13aa1n02x5               g131(.a(new_n225), .b(new_n226), .c(new_n216), .d(new_n220), .o1(new_n227));
  xorc02aa1n02x5               g132(.a(\a[22] ), .b(\b[21] ), .out0(new_n228));
  norp02aa1n02x5               g133(.a(new_n228), .b(new_n224), .o1(new_n229));
  aoi022aa1n03x5               g134(.a(new_n227), .b(new_n228), .c(new_n223), .d(new_n229), .o1(\s[22] ));
  nanp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  tech160nm_fixnrc02aa1n02p5x5 g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  nano22aa1n06x5               g137(.a(new_n232), .b(new_n225), .c(new_n231), .out0(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n214), .out0(new_n234));
  tech160nm_fioai012aa1n05x5   g139(.a(new_n234), .b(new_n188), .c(new_n182), .o1(new_n235));
  oao003aa1n12x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .carry(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  tech160nm_fiaoi012aa1n03p5x5 g142(.a(new_n237), .b(new_n219), .c(new_n233), .o1(new_n238));
  xorc02aa1n12x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xnbna2aa1n03x5               g144(.a(new_n239), .b(new_n235), .c(new_n238), .out0(\s[23] ));
  inv000aa1n02x5               g145(.a(new_n238), .o1(new_n241));
  aoai13aa1n02x7               g146(.a(new_n239), .b(new_n241), .c(new_n178), .d(new_n234), .o1(new_n242));
  nor042aa1n06x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n239), .o1(new_n245));
  aoai13aa1n02x5               g150(.a(new_n244), .b(new_n245), .c(new_n235), .d(new_n238), .o1(new_n246));
  tech160nm_fixorc02aa1n04x5   g151(.a(\a[24] ), .b(\b[23] ), .out0(new_n247));
  norp02aa1n02x5               g152(.a(new_n247), .b(new_n243), .o1(new_n248));
  aoi022aa1n02x5               g153(.a(new_n246), .b(new_n247), .c(new_n242), .d(new_n248), .o1(\s[24] ));
  nano32aa1n03x7               g154(.a(new_n214), .b(new_n247), .c(new_n233), .d(new_n239), .out0(new_n250));
  tech160nm_fioai012aa1n05x5   g155(.a(new_n250), .b(new_n188), .c(new_n182), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n218), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n233), .b(new_n252), .c(new_n213), .d(new_n204), .o1(new_n253));
  and002aa1n12x5               g158(.a(new_n247), .b(new_n239), .o(new_n254));
  inv000aa1n06x5               g159(.a(new_n254), .o1(new_n255));
  oao003aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n244), .carry(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n255), .c(new_n253), .d(new_n236), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[25] ), .b(\b[24] ), .out0(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n251), .c(new_n258), .out0(\s[25] ));
  aoai13aa1n03x5               g165(.a(new_n259), .b(new_n257), .c(new_n178), .d(new_n250), .o1(new_n261));
  nor042aa1n03x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n259), .o1(new_n264));
  aoai13aa1n02x5               g169(.a(new_n263), .b(new_n264), .c(new_n251), .d(new_n258), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  norp02aa1n02x5               g171(.a(new_n266), .b(new_n262), .o1(new_n267));
  aoi022aa1n03x5               g172(.a(new_n265), .b(new_n266), .c(new_n261), .d(new_n267), .o1(\s[26] ));
  and002aa1n12x5               g173(.a(new_n266), .b(new_n259), .o(new_n269));
  inv020aa1n03x5               g174(.a(new_n269), .o1(new_n270));
  nano23aa1n06x5               g175(.a(new_n270), .b(new_n214), .c(new_n254), .d(new_n233), .out0(new_n271));
  oai012aa1n09x5               g176(.a(new_n271), .b(new_n188), .c(new_n182), .o1(new_n272));
  oao003aa1n02x5               g177(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n273));
  aobi12aa1n12x5               g178(.a(new_n273), .b(new_n257), .c(new_n269), .out0(new_n274));
  xorc02aa1n12x5               g179(.a(\a[27] ), .b(\b[26] ), .out0(new_n275));
  xnbna2aa1n06x5               g180(.a(new_n275), .b(new_n274), .c(new_n272), .out0(\s[27] ));
  aoai13aa1n03x5               g181(.a(new_n254), .b(new_n237), .c(new_n219), .d(new_n233), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n273), .b(new_n270), .c(new_n277), .d(new_n256), .o1(new_n278));
  aoai13aa1n02x7               g183(.a(new_n275), .b(new_n278), .c(new_n178), .d(new_n271), .o1(new_n279));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1n03x5               g185(.a(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n275), .o1(new_n282));
  aoai13aa1n03x5               g187(.a(new_n281), .b(new_n282), .c(new_n274), .d(new_n272), .o1(new_n283));
  xorc02aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .out0(new_n284));
  norp02aa1n02x5               g189(.a(new_n284), .b(new_n280), .o1(new_n285));
  aoi022aa1n03x5               g190(.a(new_n283), .b(new_n284), .c(new_n279), .d(new_n285), .o1(\s[28] ));
  and002aa1n02x5               g191(.a(new_n284), .b(new_n275), .o(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n278), .c(new_n178), .d(new_n271), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n287), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n281), .carry(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n289), .c(new_n274), .d(new_n272), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .out0(new_n292));
  norb02aa1n02x5               g197(.a(new_n290), .b(new_n292), .out0(new_n293));
  aoi022aa1n03x5               g198(.a(new_n291), .b(new_n292), .c(new_n288), .d(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g200(.a(new_n282), .b(new_n284), .c(new_n292), .out0(new_n296));
  aoai13aa1n04x5               g201(.a(new_n296), .b(new_n278), .c(new_n178), .d(new_n271), .o1(new_n297));
  inv000aa1n02x5               g202(.a(new_n296), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n274), .d(new_n272), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  norb02aa1n02x5               g206(.a(new_n299), .b(new_n301), .out0(new_n302));
  aoi022aa1n03x5               g207(.a(new_n300), .b(new_n301), .c(new_n297), .d(new_n302), .o1(\s[30] ));
  xorc02aa1n02x5               g208(.a(\a[31] ), .b(\b[30] ), .out0(new_n304));
  nano32aa1d12x5               g209(.a(new_n282), .b(new_n301), .c(new_n284), .d(new_n292), .out0(new_n305));
  aoai13aa1n04x5               g210(.a(new_n305), .b(new_n278), .c(new_n178), .d(new_n271), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n305), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n307), .c(new_n274), .d(new_n272), .o1(new_n309));
  and002aa1n02x5               g214(.a(\b[29] ), .b(\a[30] ), .o(new_n310));
  oabi12aa1n02x5               g215(.a(new_n304), .b(\a[30] ), .c(\b[29] ), .out0(new_n311));
  oab012aa1n02x4               g216(.a(new_n311), .b(new_n299), .c(new_n310), .out0(new_n312));
  aoi022aa1n03x5               g217(.a(new_n309), .b(new_n304), .c(new_n306), .d(new_n312), .o1(\s[31] ));
  xorb03aa1n02x5               g218(.a(new_n106), .b(\b[2] ), .c(new_n98), .out0(\s[3] ));
  norp02aa1n02x5               g219(.a(new_n102), .b(new_n106), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[4] ), .b(\b[3] ), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n316), .b(new_n98), .c(new_n100), .o1(new_n317));
  aboi22aa1n03x5               g222(.a(new_n315), .b(new_n317), .c(new_n107), .d(new_n316), .out0(\s[4] ));
  xnrc02aa1n02x5               g223(.a(\b[4] ), .b(\a[5] ), .out0(new_n319));
  oaib12aa1n02x5               g224(.a(new_n107), .b(new_n99), .c(\b[3] ), .out0(new_n320));
  aboi22aa1n03x5               g225(.a(new_n114), .b(new_n107), .c(new_n320), .d(new_n319), .out0(\s[5] ));
  obai22aa1n02x7               g226(.a(new_n107), .b(new_n114), .c(\a[5] ), .d(\b[4] ), .out0(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  xorc02aa1n02x5               g228(.a(\a[7] ), .b(\b[6] ), .out0(new_n324));
  aoai13aa1n02x5               g229(.a(new_n324), .b(new_n108), .c(new_n322), .d(new_n110), .o1(new_n325));
  aoi112aa1n02x5               g230(.a(new_n324), .b(new_n108), .c(new_n322), .d(new_n110), .o1(new_n326));
  norb02aa1n02x5               g231(.a(new_n325), .b(new_n326), .out0(\s[7] ));
  xorc02aa1n02x5               g232(.a(\a[8] ), .b(\b[7] ), .out0(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n325), .c(new_n116), .out0(\s[8] ));
  xobna2aa1n03x5               g234(.a(new_n129), .b(new_n128), .c(new_n120), .out0(\s[9] ));
endmodule


