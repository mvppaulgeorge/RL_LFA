// Benchmark "adder" written by ABC on Wed Jul 17 14:42:57 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n337,
    new_n338, new_n339, new_n340, new_n342, new_n343, new_n345, new_n347,
    new_n348, new_n349, new_n351, new_n352, new_n353, new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  inv020aa1d32x5               g002(.a(\a[2] ), .o1(new_n98));
  inv040aa1d32x5               g003(.a(\b[1] ), .o1(new_n99));
  nand02aa1d16x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oao003aa1n09x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n101));
  nor042aa1d18x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand42aa1d28x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n24x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano23aa1n06x5               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  inv040aa1d30x5               g011(.a(\a[3] ), .o1(new_n107));
  inv040aa1d32x5               g012(.a(\b[2] ), .o1(new_n108));
  aoai13aa1n04x5               g013(.a(new_n103), .b(new_n102), .c(new_n107), .d(new_n108), .o1(new_n109));
  aobi12aa1d24x5               g014(.a(new_n109), .b(new_n106), .c(new_n101), .out0(new_n110));
  nand42aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor022aa1n16x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanb02aa1n12x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nor002aa1d32x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand02aa1d20x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanb02aa1d36x5               g020(.a(new_n114), .b(new_n115), .out0(new_n116));
  xnrc02aa1n12x5               g021(.a(\b[5] ), .b(\a[6] ), .out0(new_n117));
  inv000aa1d42x5               g022(.a(new_n117), .o1(new_n118));
  xorc02aa1n12x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nona23aa1d18x5               g024(.a(new_n118), .b(new_n119), .c(new_n116), .d(new_n113), .out0(new_n120));
  nona23aa1n02x5               g025(.a(new_n111), .b(new_n115), .c(new_n114), .d(new_n112), .out0(new_n121));
  inv040aa1d32x5               g026(.a(\a[6] ), .o1(new_n122));
  inv020aa1n16x5               g027(.a(\b[5] ), .o1(new_n123));
  norp02aa1n03x5               g028(.a(\b[4] ), .b(\a[5] ), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(new_n122), .b(new_n123), .c(new_n124), .o1(new_n125));
  inv030aa1n02x5               g030(.a(new_n114), .o1(new_n126));
  tech160nm_fioaoi03aa1n02p5x5 g031(.a(\a[8] ), .b(\b[7] ), .c(new_n126), .o1(new_n127));
  oab012aa1n12x5               g032(.a(new_n127), .b(new_n121), .c(new_n125), .out0(new_n128));
  oai012aa1d24x5               g033(.a(new_n128), .b(new_n110), .c(new_n120), .o1(new_n129));
  nor042aa1d18x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nand22aa1n12x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(new_n129), .b(new_n133), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nand02aa1d28x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n134), .c(new_n97), .out0(\s[10] ));
  nona23aa1n09x5               g043(.a(new_n136), .b(new_n131), .c(new_n130), .d(new_n135), .out0(new_n139));
  nanb02aa1n06x5               g044(.a(new_n139), .b(new_n129), .out0(new_n140));
  aoi012aa1n06x5               g045(.a(new_n135), .b(new_n130), .c(new_n136), .o1(new_n141));
  nor002aa1d32x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand02aa1d06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  inv000aa1d42x5               g049(.a(new_n144), .o1(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n140), .c(new_n141), .out0(\s[11] ));
  aob012aa1n02x5               g051(.a(new_n145), .b(new_n140), .c(new_n141), .out0(new_n147));
  nor002aa1d32x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nand02aa1n06x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  inv000aa1d42x5               g055(.a(\a[11] ), .o1(new_n151));
  inv000aa1d42x5               g056(.a(\b[10] ), .o1(new_n152));
  aboi22aa1n03x5               g057(.a(new_n148), .b(new_n149), .c(new_n151), .d(new_n152), .out0(new_n153));
  inv040aa1n08x5               g058(.a(new_n142), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n144), .c(new_n140), .d(new_n141), .o1(new_n155));
  aoi022aa1n03x5               g060(.a(new_n155), .b(new_n150), .c(new_n147), .d(new_n153), .o1(\s[12] ));
  nona23aa1n09x5               g061(.a(new_n149), .b(new_n143), .c(new_n142), .d(new_n148), .out0(new_n157));
  nor042aa1n04x5               g062(.a(new_n157), .b(new_n139), .o1(new_n158));
  oaoi03aa1n12x5               g063(.a(\a[12] ), .b(\b[11] ), .c(new_n154), .o1(new_n159));
  inv040aa1n02x5               g064(.a(new_n159), .o1(new_n160));
  tech160nm_fioai012aa1n03p5x5 g065(.a(new_n160), .b(new_n157), .c(new_n141), .o1(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[12] ), .b(\a[13] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n161), .c(new_n129), .d(new_n158), .o1(new_n164));
  aoi112aa1n02x5               g069(.a(new_n163), .b(new_n161), .c(new_n129), .d(new_n158), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(\s[13] ));
  xnrc02aa1n12x5               g071(.a(\b[13] ), .b(\a[14] ), .out0(new_n167));
  nor002aa1n03x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  oai012aa1n02x5               g074(.a(new_n164), .b(\b[12] ), .c(\a[13] ), .o1(new_n170));
  aboi22aa1n03x5               g075(.a(new_n167), .b(new_n170), .c(new_n164), .d(new_n169), .out0(\s[14] ));
  nor042aa1n06x5               g076(.a(new_n167), .b(new_n162), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n161), .c(new_n129), .d(new_n158), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nanp02aa1n02x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  aoi012aa1n02x7               g080(.a(new_n174), .b(new_n168), .c(new_n175), .o1(new_n176));
  nor002aa1d32x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanp02aa1n04x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  norb02aa1n09x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n173), .c(new_n176), .out0(\s[15] ));
  aob012aa1n03x5               g085(.a(new_n179), .b(new_n173), .c(new_n176), .out0(new_n181));
  nor022aa1n12x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nanp02aa1n04x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  aoib12aa1n02x5               g089(.a(new_n177), .b(new_n183), .c(new_n182), .out0(new_n185));
  inv000aa1d42x5               g090(.a(new_n177), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n179), .o1(new_n187));
  aoai13aa1n02x7               g092(.a(new_n186), .b(new_n187), .c(new_n173), .d(new_n176), .o1(new_n188));
  aoi022aa1n03x5               g093(.a(new_n188), .b(new_n184), .c(new_n181), .d(new_n185), .o1(\s[16] ));
  nona23aa1d18x5               g094(.a(new_n183), .b(new_n178), .c(new_n177), .d(new_n182), .out0(new_n190));
  nona32aa1n09x5               g095(.a(new_n158), .b(new_n190), .c(new_n167), .d(new_n162), .out0(new_n191));
  inv030aa1n02x5               g096(.a(new_n191), .o1(new_n192));
  nanp02aa1n09x5               g097(.a(new_n129), .b(new_n192), .o1(new_n193));
  aobi12aa1n06x5               g098(.a(new_n176), .b(new_n161), .c(new_n172), .out0(new_n194));
  oai012aa1n02x5               g099(.a(new_n183), .b(new_n182), .c(new_n177), .o1(new_n195));
  oai112aa1n06x5               g100(.a(new_n193), .b(new_n195), .c(new_n194), .d(new_n190), .o1(new_n196));
  xorb03aa1n03x5               g101(.a(new_n196), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g102(.a(\a[17] ), .o1(new_n198));
  inv040aa1d28x5               g103(.a(\b[16] ), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(new_n199), .b(new_n198), .o1(new_n200));
  oaoi13aa1n12x5               g105(.a(new_n191), .b(new_n128), .c(new_n110), .d(new_n120), .o1(new_n201));
  inv000aa1n02x5               g106(.a(new_n141), .o1(new_n202));
  nano23aa1n03x7               g107(.a(new_n142), .b(new_n148), .c(new_n149), .d(new_n143), .out0(new_n203));
  aoai13aa1n09x5               g108(.a(new_n172), .b(new_n159), .c(new_n203), .d(new_n202), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n195), .b(new_n190), .c(new_n204), .d(new_n176), .o1(new_n205));
  xorc02aa1n06x5               g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  oaih12aa1n02x5               g111(.a(new_n206), .b(new_n205), .c(new_n201), .o1(new_n207));
  nor022aa1n08x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand42aa1n16x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  norb02aa1n06x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  xnbna2aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n200), .out0(\s[18] ));
  and002aa1n02x5               g116(.a(new_n206), .b(new_n210), .o(new_n212));
  oaih12aa1n02x5               g117(.a(new_n212), .b(new_n205), .c(new_n201), .o1(new_n213));
  aoi013aa1n09x5               g118(.a(new_n208), .b(new_n209), .c(new_n198), .d(new_n199), .o1(new_n214));
  nor002aa1d32x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand42aa1n20x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n213), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fioaoi03aa1n02p5x5 g124(.a(\a[18] ), .b(\b[17] ), .c(new_n200), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n217), .b(new_n220), .c(new_n196), .d(new_n212), .o1(new_n221));
  nor002aa1d32x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand02aa1n06x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  inv000aa1d42x5               g129(.a(\a[19] ), .o1(new_n225));
  inv000aa1d42x5               g130(.a(\b[18] ), .o1(new_n226));
  aboi22aa1n03x5               g131(.a(new_n222), .b(new_n223), .c(new_n225), .d(new_n226), .out0(new_n227));
  inv040aa1n08x5               g132(.a(new_n215), .o1(new_n228));
  inv000aa1n02x5               g133(.a(new_n217), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n228), .b(new_n229), .c(new_n213), .d(new_n214), .o1(new_n230));
  aoi022aa1n03x5               g135(.a(new_n230), .b(new_n224), .c(new_n221), .d(new_n227), .o1(\s[20] ));
  nona23aa1d24x5               g136(.a(new_n223), .b(new_n216), .c(new_n215), .d(new_n222), .out0(new_n232));
  nano22aa1n12x5               g137(.a(new_n232), .b(new_n206), .c(new_n210), .out0(new_n233));
  oaih12aa1n02x5               g138(.a(new_n233), .b(new_n205), .c(new_n201), .o1(new_n234));
  oaoi03aa1n09x5               g139(.a(\a[20] ), .b(\b[19] ), .c(new_n228), .o1(new_n235));
  inv040aa1n02x5               g140(.a(new_n235), .o1(new_n236));
  oai012aa1d24x5               g141(.a(new_n236), .b(new_n232), .c(new_n214), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[20] ), .b(\a[21] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  xnbna2aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n238), .out0(\s[21] ));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n237), .c(new_n196), .d(new_n233), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  nor042aa1n06x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n243), .b(new_n245), .out0(new_n246));
  inv000aa1n09x5               g151(.a(new_n245), .o1(new_n247));
  aoai13aa1n02x5               g152(.a(new_n247), .b(new_n239), .c(new_n234), .d(new_n238), .o1(new_n248));
  aoi022aa1n03x5               g153(.a(new_n248), .b(new_n244), .c(new_n242), .d(new_n246), .o1(\s[22] ));
  nor042aa1n06x5               g154(.a(new_n243), .b(new_n239), .o1(new_n250));
  nano32aa1n02x4               g155(.a(new_n232), .b(new_n250), .c(new_n206), .d(new_n210), .out0(new_n251));
  oaih12aa1n02x5               g156(.a(new_n251), .b(new_n205), .c(new_n201), .o1(new_n252));
  oaoi03aa1n03x5               g157(.a(\a[22] ), .b(\b[21] ), .c(new_n247), .o1(new_n253));
  aoi012aa1n02x5               g158(.a(new_n253), .b(new_n237), .c(new_n250), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  xnbna2aa1n03x5               g160(.a(new_n255), .b(new_n252), .c(new_n254), .out0(\s[23] ));
  inv000aa1n02x5               g161(.a(new_n254), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n255), .b(new_n257), .c(new_n196), .d(new_n251), .o1(new_n258));
  tech160nm_fixorc02aa1n02p5x5 g163(.a(\a[24] ), .b(\b[23] ), .out0(new_n259));
  nor042aa1n09x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  norp02aa1n02x5               g165(.a(new_n259), .b(new_n260), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n260), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n255), .o1(new_n263));
  aoai13aa1n02x5               g168(.a(new_n262), .b(new_n263), .c(new_n252), .d(new_n254), .o1(new_n264));
  aoi022aa1n03x5               g169(.a(new_n264), .b(new_n259), .c(new_n258), .d(new_n261), .o1(\s[24] ));
  inv000aa1d42x5               g170(.a(new_n233), .o1(new_n266));
  and002aa1n06x5               g171(.a(new_n259), .b(new_n255), .o(new_n267));
  nano22aa1n02x4               g172(.a(new_n266), .b(new_n267), .c(new_n250), .out0(new_n268));
  oaih12aa1n02x5               g173(.a(new_n268), .b(new_n205), .c(new_n201), .o1(new_n269));
  nano23aa1n03x7               g174(.a(new_n215), .b(new_n222), .c(new_n223), .d(new_n216), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n250), .b(new_n235), .c(new_n270), .d(new_n220), .o1(new_n271));
  inv000aa1n02x5               g176(.a(new_n253), .o1(new_n272));
  inv000aa1n06x5               g177(.a(new_n267), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[24] ), .b(\b[23] ), .c(new_n262), .carry(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n271), .d(new_n272), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n269), .c(new_n276), .out0(\s[25] ));
  aoai13aa1n03x5               g183(.a(new_n277), .b(new_n275), .c(new_n196), .d(new_n268), .o1(new_n279));
  xorc02aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .out0(new_n280));
  norp02aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .o1(new_n281));
  norp02aa1n02x5               g186(.a(new_n280), .b(new_n281), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n281), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n277), .o1(new_n284));
  aoai13aa1n02x5               g189(.a(new_n283), .b(new_n284), .c(new_n269), .d(new_n276), .o1(new_n285));
  aoi022aa1n03x5               g190(.a(new_n285), .b(new_n280), .c(new_n279), .d(new_n282), .o1(\s[26] ));
  and002aa1n06x5               g191(.a(new_n280), .b(new_n277), .o(new_n287));
  inv000aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nano32aa1n03x7               g193(.a(new_n288), .b(new_n233), .c(new_n267), .d(new_n250), .out0(new_n289));
  oai012aa1n06x5               g194(.a(new_n289), .b(new_n205), .c(new_n201), .o1(new_n290));
  nanp02aa1n02x5               g195(.a(\b[25] ), .b(\a[26] ), .o1(new_n291));
  oai022aa1n02x5               g196(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n292));
  aoi022aa1n06x5               g197(.a(new_n275), .b(new_n287), .c(new_n291), .d(new_n292), .o1(new_n293));
  nand42aa1n02x5               g198(.a(new_n290), .b(new_n293), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoi122aa1n02x7               g200(.a(new_n295), .b(new_n291), .c(new_n292), .d(new_n275), .e(new_n287), .o1(new_n296));
  aoi022aa1n02x7               g201(.a(new_n294), .b(new_n295), .c(new_n296), .d(new_n290), .o1(\s[27] ));
  aoai13aa1n02x5               g202(.a(new_n267), .b(new_n253), .c(new_n237), .d(new_n250), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n292), .b(new_n291), .o1(new_n299));
  aoai13aa1n04x5               g204(.a(new_n299), .b(new_n288), .c(new_n298), .d(new_n274), .o1(new_n300));
  aoai13aa1n02x7               g205(.a(new_n295), .b(new_n300), .c(new_n196), .d(new_n289), .o1(new_n301));
  tech160nm_fixorc02aa1n03p5x5 g206(.a(\a[28] ), .b(\b[27] ), .out0(new_n302));
  norp02aa1n02x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  norp02aa1n02x5               g208(.a(new_n302), .b(new_n303), .o1(new_n304));
  inv000aa1n03x5               g209(.a(new_n303), .o1(new_n305));
  inv020aa1n02x5               g210(.a(new_n295), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n305), .b(new_n306), .c(new_n290), .d(new_n293), .o1(new_n307));
  aoi022aa1n03x5               g212(.a(new_n307), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[28] ));
  and002aa1n02x5               g213(.a(new_n302), .b(new_n295), .o(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n300), .c(new_n196), .d(new_n289), .o1(new_n310));
  tech160nm_fixorc02aa1n03p5x5 g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  oao003aa1n02x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n305), .carry(new_n312));
  norb02aa1n02x5               g217(.a(new_n312), .b(new_n311), .out0(new_n313));
  inv000aa1d42x5               g218(.a(new_n309), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n312), .b(new_n314), .c(new_n290), .d(new_n293), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n310), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g221(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g222(.a(new_n306), .b(new_n302), .c(new_n311), .out0(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n300), .c(new_n196), .d(new_n289), .o1(new_n319));
  tech160nm_fixorc02aa1n05x5   g224(.a(\a[30] ), .b(\b[29] ), .out0(new_n320));
  and002aa1n02x5               g225(.a(\b[28] ), .b(\a[29] ), .o(new_n321));
  oabi12aa1n02x5               g226(.a(new_n320), .b(\a[29] ), .c(\b[28] ), .out0(new_n322));
  oab012aa1n02x4               g227(.a(new_n322), .b(new_n312), .c(new_n321), .out0(new_n323));
  inv000aa1d42x5               g228(.a(new_n318), .o1(new_n324));
  oaoi03aa1n02x5               g229(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .o1(new_n325));
  inv000aa1n03x5               g230(.a(new_n325), .o1(new_n326));
  aoai13aa1n02x7               g231(.a(new_n326), .b(new_n324), .c(new_n290), .d(new_n293), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n320), .c(new_n319), .d(new_n323), .o1(\s[30] ));
  nano32aa1n02x5               g233(.a(new_n306), .b(new_n320), .c(new_n302), .d(new_n311), .out0(new_n329));
  aoai13aa1n02x7               g234(.a(new_n329), .b(new_n300), .c(new_n196), .d(new_n289), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  oao003aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n332));
  norb02aa1n02x5               g237(.a(new_n332), .b(new_n331), .out0(new_n333));
  inv000aa1n02x5               g238(.a(new_n329), .o1(new_n334));
  aoai13aa1n03x5               g239(.a(new_n332), .b(new_n334), .c(new_n290), .d(new_n293), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n335), .b(new_n331), .c(new_n330), .d(new_n333), .o1(\s[31] ));
  aoi022aa1n02x5               g241(.a(new_n99), .b(new_n98), .c(\a[1] ), .d(\b[0] ), .o1(new_n337));
  oaib12aa1n02x5               g242(.a(new_n337), .b(new_n99), .c(\a[2] ), .out0(new_n338));
  norb02aa1n02x5               g243(.a(new_n105), .b(new_n104), .out0(new_n339));
  aboi22aa1n03x5               g244(.a(new_n104), .b(new_n105), .c(new_n98), .d(new_n99), .out0(new_n340));
  aoi022aa1n02x5               g245(.a(new_n101), .b(new_n339), .c(new_n338), .d(new_n340), .o1(\s[3] ));
  obai22aa1n02x7               g246(.a(new_n103), .b(new_n102), .c(\a[3] ), .d(\b[2] ), .out0(new_n342));
  aoi012aa1n02x5               g247(.a(new_n342), .b(new_n101), .c(new_n339), .o1(new_n343));
  oab012aa1n02x4               g248(.a(new_n343), .b(new_n110), .c(new_n102), .out0(\s[4] ));
  nanp02aa1n02x5               g249(.a(new_n106), .b(new_n101), .o1(new_n345));
  xnbna2aa1n03x5               g250(.a(new_n119), .b(new_n345), .c(new_n109), .out0(\s[5] ));
  oaoi03aa1n02x5               g251(.a(\a[5] ), .b(\b[4] ), .c(new_n110), .o1(new_n347));
  norp02aa1n02x5               g252(.a(new_n117), .b(new_n124), .o1(new_n348));
  oaib12aa1n06x5               g253(.a(new_n348), .b(new_n110), .c(new_n119), .out0(new_n349));
  aob012aa1n02x5               g254(.a(new_n349), .b(new_n347), .c(new_n117), .out0(\s[6] ));
  inv000aa1d42x5               g255(.a(new_n116), .o1(new_n351));
  oaoi13aa1n02x5               g256(.a(new_n351), .b(new_n349), .c(new_n122), .d(new_n123), .o1(new_n352));
  oai112aa1n02x5               g257(.a(new_n349), .b(new_n351), .c(new_n123), .d(new_n122), .o1(new_n353));
  norb02aa1n02x5               g258(.a(new_n353), .b(new_n352), .out0(\s[7] ));
  xobna2aa1n03x5               g259(.a(new_n113), .b(new_n353), .c(new_n126), .out0(\s[8] ));
  oai112aa1n02x5               g260(.a(new_n128), .b(new_n132), .c(new_n110), .d(new_n120), .o1(new_n356));
  aobi12aa1n02x5               g261(.a(new_n356), .b(new_n133), .c(new_n129), .out0(\s[9] ));
endmodule


