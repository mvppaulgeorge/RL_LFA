// Benchmark "adder" written by ABC on Thu Jul 18 01:13:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n323, new_n324,
    new_n327, new_n328, new_n329, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  norp02aa1n09x5               g004(.a(\b[5] ), .b(\a[6] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[4] ), .b(\a[5] ), .o1(new_n102));
  nand42aa1n06x5               g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  nano23aa1n06x5               g008(.a(new_n100), .b(new_n102), .c(new_n103), .d(new_n101), .out0(new_n104));
  nor002aa1d32x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nand02aa1d08x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nor042aa1n06x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand02aa1n06x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nona23aa1n09x5               g013(.a(new_n108), .b(new_n106), .c(new_n105), .d(new_n107), .out0(new_n109));
  norb02aa1n06x5               g014(.a(new_n104), .b(new_n109), .out0(new_n110));
  nor042aa1n04x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  nand42aa1n06x5               g016(.a(\b[0] ), .b(\a[1] ), .o1(new_n112));
  nanp02aa1n12x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  aoi012aa1d18x5               g018(.a(new_n111), .b(new_n112), .c(new_n113), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  nand02aa1n08x5               g020(.a(\b[3] ), .b(\a[4] ), .o1(new_n116));
  nor022aa1n16x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  nanp02aa1n04x5               g022(.a(\b[2] ), .b(\a[3] ), .o1(new_n118));
  nona23aa1n09x5               g023(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n119));
  aoi012aa1n09x5               g024(.a(new_n115), .b(new_n117), .c(new_n116), .o1(new_n120));
  oaih12aa1n12x5               g025(.a(new_n120), .b(new_n119), .c(new_n114), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n105), .o1(new_n122));
  nand42aa1n03x5               g027(.a(new_n107), .b(new_n106), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\a[5] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[4] ), .o1(new_n125));
  aoai13aa1n04x5               g030(.a(new_n101), .b(new_n100), .c(new_n124), .d(new_n125), .o1(new_n126));
  oai112aa1n06x5               g031(.a(new_n122), .b(new_n123), .c(new_n109), .d(new_n126), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n127), .c(new_n110), .d(new_n121), .o1(new_n129));
  nor002aa1d32x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand02aa1d16x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n15x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g038(.a(new_n130), .o1(new_n134));
  inv000aa1d42x5               g039(.a(new_n132), .o1(new_n135));
  aoai13aa1n04x5               g040(.a(new_n134), .b(new_n135), .c(new_n129), .d(new_n99), .o1(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand42aa1d28x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  nor002aa1d32x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1d28x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  aoi112aa1n02x5               g048(.a(new_n143), .b(new_n138), .c(new_n136), .d(new_n140), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n143), .b(new_n138), .c(new_n136), .d(new_n139), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(\s[12] ));
  nanb02aa1n02x5               g051(.a(new_n105), .b(new_n106), .out0(new_n147));
  nanb02aa1n02x5               g052(.a(new_n107), .b(new_n108), .out0(new_n148));
  nona22aa1n02x4               g053(.a(new_n104), .b(new_n147), .c(new_n148), .out0(new_n149));
  inv000aa1n06x5               g054(.a(new_n114), .o1(new_n150));
  nano23aa1n02x5               g055(.a(new_n115), .b(new_n117), .c(new_n118), .d(new_n116), .out0(new_n151));
  aobi12aa1n03x5               g056(.a(new_n120), .b(new_n151), .c(new_n150), .out0(new_n152));
  norp03aa1n02x5               g057(.a(new_n126), .b(new_n148), .c(new_n147), .o1(new_n153));
  nano22aa1n03x5               g058(.a(new_n153), .b(new_n122), .c(new_n123), .out0(new_n154));
  tech160nm_fioai012aa1n05x5   g059(.a(new_n154), .b(new_n152), .c(new_n149), .o1(new_n155));
  nano23aa1d15x5               g060(.a(new_n138), .b(new_n141), .c(new_n142), .d(new_n139), .out0(new_n156));
  nand23aa1d12x5               g061(.a(new_n156), .b(new_n128), .c(new_n132), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nona23aa1n12x5               g063(.a(new_n142), .b(new_n139), .c(new_n138), .d(new_n141), .out0(new_n159));
  tech160nm_fioai012aa1n03p5x5 g064(.a(new_n142), .b(new_n141), .c(new_n138), .o1(new_n160));
  aoai13aa1n12x5               g065(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n161));
  oai012aa1d24x5               g066(.a(new_n160), .b(new_n159), .c(new_n161), .o1(new_n162));
  tech160nm_fiaoi012aa1n05x5   g067(.a(new_n162), .b(new_n155), .c(new_n158), .o1(new_n163));
  xnrb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n02x5               g069(.a(\a[13] ), .b(\b[12] ), .c(new_n163), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  aoai13aa1n03x5               g071(.a(new_n158), .b(new_n127), .c(new_n110), .d(new_n121), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n162), .o1(new_n168));
  norp02aa1n09x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  tech160nm_finand02aa1n03p5x5 g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  nor002aa1n12x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nanp02aa1n04x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nona23aa1n03x5               g077(.a(new_n172), .b(new_n170), .c(new_n169), .d(new_n171), .out0(new_n173));
  oai012aa1n06x5               g078(.a(new_n172), .b(new_n171), .c(new_n169), .o1(new_n174));
  aoai13aa1n03x5               g079(.a(new_n174), .b(new_n173), .c(new_n167), .d(new_n168), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  tech160nm_fixorc02aa1n03p5x5 g082(.a(\a[15] ), .b(\b[14] ), .out0(new_n178));
  xnrc02aa1n12x5               g083(.a(\b[15] ), .b(\a[16] ), .out0(new_n179));
  inv040aa1n02x5               g084(.a(new_n179), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n177), .b(new_n180), .c(new_n175), .d(new_n178), .o1(new_n181));
  aoai13aa1n03x5               g086(.a(new_n180), .b(new_n177), .c(new_n175), .d(new_n178), .o1(new_n182));
  norb02aa1n02x7               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano23aa1n06x5               g088(.a(new_n169), .b(new_n171), .c(new_n172), .d(new_n170), .out0(new_n184));
  nano32aa1d12x5               g089(.a(new_n157), .b(new_n180), .c(new_n184), .d(new_n178), .out0(new_n185));
  aoai13aa1n12x5               g090(.a(new_n185), .b(new_n127), .c(new_n110), .d(new_n121), .o1(new_n186));
  tech160nm_fixnrc02aa1n03p5x5 g091(.a(\b[14] ), .b(\a[15] ), .out0(new_n187));
  nor003aa1n03x5               g092(.a(new_n173), .b(new_n187), .c(new_n179), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n189));
  nor002aa1n04x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n190), .o1(new_n191));
  oai013aa1n03x5               g096(.a(new_n191), .b(new_n187), .c(new_n179), .d(new_n174), .o1(new_n192));
  aoi112aa1n09x5               g097(.a(new_n192), .b(new_n189), .c(new_n162), .d(new_n188), .o1(new_n193));
  xorc02aa1n02x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n186), .c(new_n193), .out0(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[17] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[16] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(new_n162), .b(new_n188), .o1(new_n199));
  nona22aa1n03x5               g104(.a(new_n199), .b(new_n192), .c(new_n189), .out0(new_n200));
  aoai13aa1n02x5               g105(.a(new_n194), .b(new_n200), .c(new_n155), .d(new_n185), .o1(new_n201));
  nor042aa1n06x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nanp02aa1n06x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nanb02aa1n12x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  xobna2aa1n03x5               g109(.a(new_n204), .b(new_n201), .c(new_n198), .out0(\s[18] ));
  nanp02aa1n02x5               g110(.a(\b[16] ), .b(\a[17] ), .o1(new_n206));
  nano22aa1d15x5               g111(.a(new_n204), .b(new_n198), .c(new_n206), .out0(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  aoai13aa1n04x5               g113(.a(new_n203), .b(new_n202), .c(new_n196), .d(new_n197), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n208), .c(new_n186), .d(new_n193), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand42aa1n08x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  inv000aa1d42x5               g119(.a(\b[19] ), .o1(new_n215));
  nanb02aa1n06x5               g120(.a(\a[20] ), .b(new_n215), .out0(new_n216));
  nand42aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  aoi122aa1n03x5               g122(.a(new_n213), .b(new_n216), .c(new_n217), .d(new_n210), .e(new_n214), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n213), .o1(new_n219));
  nanb02aa1n12x5               g124(.a(new_n213), .b(new_n214), .out0(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  nand02aa1n02x5               g126(.a(new_n210), .b(new_n221), .o1(new_n222));
  nand02aa1n03x5               g127(.a(new_n216), .b(new_n217), .o1(new_n223));
  tech160nm_fiaoi012aa1n02p5x5 g128(.a(new_n223), .b(new_n222), .c(new_n219), .o1(new_n224));
  norp02aa1n03x5               g129(.a(new_n224), .b(new_n218), .o1(\s[20] ));
  nona22aa1n02x4               g130(.a(new_n207), .b(new_n220), .c(new_n223), .out0(new_n226));
  nand42aa1n02x5               g131(.a(new_n213), .b(new_n217), .o1(new_n227));
  nor043aa1n03x5               g132(.a(new_n209), .b(new_n220), .c(new_n223), .o1(new_n228));
  nano22aa1n03x7               g133(.a(new_n228), .b(new_n216), .c(new_n227), .out0(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n226), .c(new_n186), .d(new_n193), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[20] ), .b(\a[21] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[21] ), .b(\a[22] ), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi112aa1n03x4               g141(.a(new_n232), .b(new_n236), .c(new_n230), .d(new_n234), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n232), .c(new_n230), .d(new_n234), .o1(new_n238));
  norb02aa1n02x7               g143(.a(new_n238), .b(new_n237), .out0(\s[22] ));
  nor022aa1n04x5               g144(.a(\b[19] ), .b(\a[20] ), .o1(new_n240));
  nona23aa1n09x5               g145(.a(new_n217), .b(new_n214), .c(new_n213), .d(new_n240), .out0(new_n241));
  nor042aa1n06x5               g146(.a(new_n235), .b(new_n233), .o1(new_n242));
  nanb03aa1d18x5               g147(.a(new_n241), .b(new_n242), .c(new_n207), .out0(new_n243));
  oai112aa1n04x5               g148(.a(new_n227), .b(new_n216), .c(new_n241), .d(new_n209), .o1(new_n244));
  oai022aa1n02x5               g149(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n245));
  aob012aa1n02x5               g150(.a(new_n245), .b(\b[21] ), .c(\a[22] ), .out0(new_n246));
  aobi12aa1n02x5               g151(.a(new_n246), .b(new_n244), .c(new_n242), .out0(new_n247));
  aoai13aa1n04x5               g152(.a(new_n247), .b(new_n243), .c(new_n186), .d(new_n193), .o1(new_n248));
  xorb03aa1n02x5               g153(.a(new_n248), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  tech160nm_fixorc02aa1n05x5   g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  tech160nm_fixorc02aa1n05x5   g156(.a(\a[24] ), .b(\b[23] ), .out0(new_n252));
  aoi112aa1n02x5               g157(.a(new_n250), .b(new_n252), .c(new_n248), .d(new_n251), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n252), .b(new_n250), .c(new_n248), .d(new_n251), .o1(new_n254));
  norb02aa1n02x7               g159(.a(new_n254), .b(new_n253), .out0(\s[24] ));
  nanp02aa1n03x5               g160(.a(new_n252), .b(new_n251), .o1(new_n256));
  nona23aa1n02x4               g161(.a(new_n242), .b(new_n207), .c(new_n256), .d(new_n241), .out0(new_n257));
  inv000aa1d42x5               g162(.a(\a[23] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(\a[24] ), .o1(new_n259));
  xroi22aa1d04x5               g164(.a(new_n258), .b(\b[22] ), .c(new_n259), .d(\b[23] ), .out0(new_n260));
  inv000aa1d42x5               g165(.a(\b[23] ), .o1(new_n261));
  oaoi03aa1n02x5               g166(.a(new_n259), .b(new_n261), .c(new_n250), .o1(new_n262));
  tech160nm_fioai012aa1n05x5   g167(.a(new_n262), .b(new_n256), .c(new_n246), .o1(new_n263));
  aoi013aa1n06x4               g168(.a(new_n263), .b(new_n244), .c(new_n242), .d(new_n260), .o1(new_n264));
  aoai13aa1n04x5               g169(.a(new_n264), .b(new_n257), .c(new_n186), .d(new_n193), .o1(new_n265));
  xorb03aa1n02x5               g170(.a(new_n265), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor002aa1n03x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  xorc02aa1n12x5               g172(.a(\a[25] ), .b(\b[24] ), .out0(new_n268));
  xorc02aa1n12x5               g173(.a(\a[26] ), .b(\b[25] ), .out0(new_n269));
  aoi112aa1n03x4               g174(.a(new_n267), .b(new_n269), .c(new_n265), .d(new_n268), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n269), .b(new_n267), .c(new_n265), .d(new_n268), .o1(new_n271));
  norb02aa1n02x7               g176(.a(new_n271), .b(new_n270), .out0(\s[26] ));
  and002aa1n06x5               g177(.a(new_n269), .b(new_n268), .o(new_n273));
  nano22aa1n12x5               g178(.a(new_n243), .b(new_n273), .c(new_n260), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n200), .c(new_n155), .d(new_n185), .o1(new_n275));
  nano22aa1n03x5               g180(.a(new_n229), .b(new_n242), .c(new_n260), .out0(new_n276));
  inv000aa1d42x5               g181(.a(\a[26] ), .o1(new_n277));
  inv000aa1d42x5               g182(.a(\b[25] ), .o1(new_n278));
  tech160nm_fioaoi03aa1n03p5x5 g183(.a(new_n277), .b(new_n278), .c(new_n267), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  oaoi13aa1n09x5               g185(.a(new_n280), .b(new_n273), .c(new_n276), .d(new_n263), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n275), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  aobi12aa1n02x7               g190(.a(new_n282), .b(new_n281), .c(new_n275), .out0(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[27] ), .b(\a[28] ), .out0(new_n287));
  nano22aa1n03x5               g192(.a(new_n286), .b(new_n285), .c(new_n287), .out0(new_n288));
  nanp02aa1n06x5               g193(.a(new_n186), .b(new_n193), .o1(new_n289));
  nona32aa1n02x5               g194(.a(new_n244), .b(new_n256), .c(new_n235), .d(new_n233), .out0(new_n290));
  inv040aa1n02x5               g195(.a(new_n263), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n273), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n279), .b(new_n292), .c(new_n290), .d(new_n291), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n282), .b(new_n293), .c(new_n289), .d(new_n274), .o1(new_n294));
  tech160nm_fiaoi012aa1n02p5x5 g199(.a(new_n287), .b(new_n294), .c(new_n285), .o1(new_n295));
  norp02aa1n03x5               g200(.a(new_n295), .b(new_n288), .o1(\s[28] ));
  norb02aa1n02x5               g201(.a(new_n282), .b(new_n287), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n293), .c(new_n289), .d(new_n274), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[28] ), .b(\a[29] ), .out0(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n298), .c(new_n299), .o1(new_n301));
  aobi12aa1n02x7               g206(.a(new_n297), .b(new_n281), .c(new_n275), .out0(new_n302));
  nano22aa1n02x4               g207(.a(new_n302), .b(new_n299), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n112), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g210(.a(new_n282), .b(new_n300), .c(new_n287), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n293), .c(new_n289), .d(new_n274), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n299), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[29] ), .b(\a[30] ), .out0(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  aobi12aa1n02x7               g215(.a(new_n306), .b(new_n281), .c(new_n275), .out0(new_n311));
  nano22aa1n02x4               g216(.a(new_n311), .b(new_n308), .c(new_n309), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n310), .b(new_n312), .o1(\s[30] ));
  xnrc02aa1n02x5               g218(.a(\b[30] ), .b(\a[31] ), .out0(new_n314));
  norb02aa1n02x7               g219(.a(new_n306), .b(new_n309), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n293), .c(new_n289), .d(new_n274), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n317));
  tech160nm_fiaoi012aa1n02p5x5 g222(.a(new_n314), .b(new_n316), .c(new_n317), .o1(new_n318));
  aobi12aa1n02x7               g223(.a(new_n315), .b(new_n281), .c(new_n275), .out0(new_n319));
  nano22aa1n02x4               g224(.a(new_n319), .b(new_n314), .c(new_n317), .out0(new_n320));
  norp02aa1n03x5               g225(.a(new_n318), .b(new_n320), .o1(\s[31] ));
  xnrb03aa1n02x5               g226(.a(new_n114), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g227(.a(new_n115), .o1(new_n323));
  aoi122aa1n02x5               g228(.a(new_n117), .b(new_n323), .c(new_n116), .d(new_n150), .e(new_n118), .o1(new_n324));
  aoi012aa1n02x5               g229(.a(new_n324), .b(new_n323), .c(new_n121), .o1(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  orn002aa1n02x5               g231(.a(\a[6] ), .b(\b[5] ), .o(new_n327));
  oaib12aa1n02x5               g232(.a(new_n126), .b(new_n152), .c(new_n104), .out0(new_n328));
  aoi122aa1n02x5               g233(.a(new_n102), .b(new_n101), .c(new_n327), .d(new_n121), .e(new_n103), .o1(new_n329));
  aoi012aa1n02x5               g234(.a(new_n329), .b(new_n328), .c(new_n327), .o1(\s[6] ));
  xorb03aa1n02x5               g235(.a(new_n328), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g236(.a(new_n107), .b(new_n328), .c(new_n108), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n122), .c(new_n106), .out0(\s[8] ));
  xorb03aa1n02x5               g238(.a(new_n155), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


