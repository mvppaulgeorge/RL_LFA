// Benchmark "adder" written by ABC on Thu Jul 18 03:29:46 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n326, new_n328, new_n329, new_n332, new_n334,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n09x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand22aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n06x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(new_n102), .o1(new_n103));
  nand02aa1d24x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nand02aa1d06x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  norb03aa1n02x7               g011(.a(new_n105), .b(new_n104), .c(new_n106), .out0(new_n107));
  nor002aa1n16x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  tech160nm_finand02aa1n03p5x5 g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanb03aa1n02x5               g014(.a(new_n108), .b(new_n109), .c(new_n105), .out0(new_n110));
  oab012aa1n09x5               g015(.a(new_n108), .b(\a[4] ), .c(\b[3] ), .out0(new_n111));
  oaoi13aa1n04x5               g016(.a(new_n103), .b(new_n111), .c(new_n107), .d(new_n110), .o1(new_n112));
  nor042aa1n06x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1d28x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor042aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n08x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .out0(new_n118));
  tech160nm_fixnrc02aa1n02p5x5 g023(.a(\b[4] ), .b(\a[5] ), .out0(new_n119));
  nor043aa1n02x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  nano23aa1n09x5               g025(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n121));
  oa0012aa1n02x5               g026(.a(new_n114), .b(new_n115), .c(new_n113), .o(new_n122));
  inv000aa1d42x5               g027(.a(\a[5] ), .o1(new_n123));
  nanb02aa1n12x5               g028(.a(\b[4] ), .b(new_n123), .out0(new_n124));
  oaoi03aa1n06x5               g029(.a(\a[6] ), .b(\b[5] ), .c(new_n124), .o1(new_n125));
  aoi012aa1n12x5               g030(.a(new_n122), .b(new_n121), .c(new_n125), .o1(new_n126));
  inv000aa1d42x5               g031(.a(new_n126), .o1(new_n127));
  nand02aa1d06x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n06x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n127), .c(new_n112), .d(new_n120), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  nona22aa1n03x5               g036(.a(new_n105), .b(new_n106), .c(new_n104), .out0(new_n132));
  nano22aa1n03x7               g037(.a(new_n108), .b(new_n105), .c(new_n109), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n111), .o1(new_n134));
  aoai13aa1n09x5               g039(.a(new_n102), .b(new_n134), .c(new_n133), .d(new_n132), .o1(new_n135));
  nona22aa1n03x5               g040(.a(new_n121), .b(new_n118), .c(new_n119), .out0(new_n136));
  oai012aa1n02x5               g041(.a(new_n126), .b(new_n135), .c(new_n136), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n99), .b(new_n100), .c(new_n137), .d(new_n128), .o1(new_n138));
  tech160nm_fioai012aa1n03p5x5 g043(.a(new_n98), .b(new_n100), .c(new_n97), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nand02aa1n04x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n139), .out0(\s[11] ));
  inv000aa1d42x5               g048(.a(new_n140), .o1(new_n144));
  nanp02aa1n03x5               g049(.a(new_n130), .b(new_n101), .o1(new_n145));
  inv040aa1n06x5               g050(.a(new_n139), .o1(new_n146));
  aoai13aa1n02x5               g051(.a(new_n142), .b(new_n146), .c(new_n145), .d(new_n99), .o1(new_n147));
  nor022aa1n12x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nanp02aa1n04x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  aobi12aa1n06x5               g055(.a(new_n150), .b(new_n147), .c(new_n144), .out0(new_n151));
  nona22aa1n02x4               g056(.a(new_n147), .b(new_n150), .c(new_n140), .out0(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(\s[12] ));
  nona23aa1d18x5               g058(.a(new_n149), .b(new_n141), .c(new_n140), .d(new_n148), .out0(new_n154));
  nano22aa1n03x7               g059(.a(new_n154), .b(new_n99), .c(new_n129), .out0(new_n155));
  aoai13aa1n02x5               g060(.a(new_n155), .b(new_n127), .c(new_n112), .d(new_n120), .o1(new_n156));
  oaoi03aa1n12x5               g061(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n157));
  oabi12aa1n12x5               g062(.a(new_n157), .b(new_n154), .c(new_n139), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  norp02aa1n09x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand42aa1n03x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nanb02aa1n03x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  xobna2aa1n03x5               g067(.a(new_n162), .b(new_n156), .c(new_n159), .out0(\s[13] ));
  oai012aa1n02x5               g068(.a(new_n111), .b(new_n107), .c(new_n110), .o1(new_n164));
  nanp03aa1n02x5               g069(.a(new_n120), .b(new_n164), .c(new_n102), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n140), .b(new_n148), .c(new_n149), .d(new_n141), .out0(new_n166));
  nanp03aa1n02x5               g071(.a(new_n166), .b(new_n99), .c(new_n129), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n159), .b(new_n167), .c(new_n165), .d(new_n126), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n160), .b(new_n168), .c(new_n161), .o1(new_n169));
  xnrb03aa1n02x5               g074(.a(new_n169), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1n02x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nano23aa1n06x5               g077(.a(new_n160), .b(new_n171), .c(new_n172), .d(new_n161), .out0(new_n173));
  oai012aa1n09x5               g078(.a(new_n172), .b(new_n171), .c(new_n160), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  nor022aa1n12x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  tech160nm_finand02aa1n03p5x5 g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n175), .c(new_n168), .d(new_n173), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n175), .c(new_n168), .d(new_n173), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(\s[15] ));
  nor022aa1n16x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nand42aa1n04x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n183), .b(new_n184), .out0(new_n185));
  oaoi13aa1n02x5               g090(.a(new_n185), .b(new_n180), .c(\a[15] ), .d(\b[14] ), .o1(new_n186));
  oai112aa1n02x5               g091(.a(new_n180), .b(new_n185), .c(\b[14] ), .d(\a[15] ), .o1(new_n187));
  norb02aa1n02x7               g092(.a(new_n187), .b(new_n186), .out0(\s[16] ));
  nanb02aa1n03x5               g093(.a(new_n171), .b(new_n172), .out0(new_n189));
  nona23aa1d16x5               g094(.a(new_n184), .b(new_n177), .c(new_n176), .d(new_n183), .out0(new_n190));
  nona32aa1n09x5               g095(.a(new_n155), .b(new_n190), .c(new_n189), .d(new_n162), .out0(new_n191));
  oaoi13aa1n12x5               g096(.a(new_n191), .b(new_n126), .c(new_n135), .d(new_n136), .o1(new_n192));
  aoai13aa1n12x5               g097(.a(new_n173), .b(new_n157), .c(new_n166), .d(new_n146), .o1(new_n193));
  tech160nm_fiaoi012aa1n03p5x5 g098(.a(new_n183), .b(new_n176), .c(new_n184), .o1(new_n194));
  aoai13aa1n12x5               g099(.a(new_n194), .b(new_n190), .c(new_n193), .d(new_n174), .o1(new_n195));
  nor042aa1n06x5               g100(.a(new_n195), .b(new_n192), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\a[17] ), .o1(new_n197));
  inv000aa1d42x5               g102(.a(\b[16] ), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(new_n198), .b(new_n197), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n196), .b(new_n200), .c(new_n199), .out0(\s[17] ));
  nor002aa1d32x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nanp02aa1n24x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nanb02aa1n06x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  tech160nm_fioaoi03aa1n03p5x5 g109(.a(\a[17] ), .b(\b[16] ), .c(new_n196), .o1(new_n205));
  xnrc02aa1n02x5               g110(.a(new_n205), .b(new_n204), .out0(\s[18] ));
  nano22aa1n03x7               g111(.a(new_n204), .b(new_n199), .c(new_n200), .out0(new_n207));
  oai012aa1n06x5               g112(.a(new_n207), .b(new_n195), .c(new_n192), .o1(new_n208));
  aoai13aa1n12x5               g113(.a(new_n203), .b(new_n202), .c(new_n197), .d(new_n198), .o1(new_n209));
  nor042aa1n09x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nand42aa1n02x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  xobna2aa1n03x5               g117(.a(new_n212), .b(new_n208), .c(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv020aa1n06x5               g119(.a(new_n209), .o1(new_n215));
  oaoi13aa1n06x5               g120(.a(new_n215), .b(new_n207), .c(new_n195), .d(new_n192), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n210), .o1(new_n217));
  nor042aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand02aa1n04x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nanb02aa1n02x5               g124(.a(new_n218), .b(new_n219), .out0(new_n220));
  oaoi13aa1n02x7               g125(.a(new_n220), .b(new_n217), .c(new_n216), .d(new_n212), .o1(new_n221));
  tech160nm_fiaoi012aa1n02p5x5 g126(.a(new_n212), .b(new_n208), .c(new_n209), .o1(new_n222));
  nano22aa1n03x5               g127(.a(new_n222), .b(new_n217), .c(new_n220), .out0(new_n223));
  norp02aa1n03x5               g128(.a(new_n221), .b(new_n223), .o1(\s[20] ));
  nano23aa1n06x5               g129(.a(new_n210), .b(new_n218), .c(new_n219), .d(new_n211), .out0(new_n225));
  nand02aa1d04x5               g130(.a(new_n207), .b(new_n225), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nona23aa1n09x5               g132(.a(new_n219), .b(new_n211), .c(new_n210), .d(new_n218), .out0(new_n228));
  tech160nm_fiaoi012aa1n05x5   g133(.a(new_n218), .b(new_n210), .c(new_n219), .o1(new_n229));
  oai012aa1n18x5               g134(.a(new_n229), .b(new_n228), .c(new_n209), .o1(new_n230));
  oaoi13aa1n06x5               g135(.a(new_n230), .b(new_n227), .c(new_n195), .d(new_n192), .o1(new_n231));
  xnrb03aa1n03x5               g136(.a(new_n231), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n03x5               g139(.a(\b[20] ), .b(\a[21] ), .out0(new_n235));
  xnrc02aa1n03x5               g140(.a(\b[21] ), .b(\a[22] ), .out0(new_n236));
  oaoi13aa1n02x7               g141(.a(new_n236), .b(new_n234), .c(new_n231), .d(new_n235), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n230), .o1(new_n238));
  oaoi13aa1n02x7               g143(.a(new_n235), .b(new_n238), .c(new_n196), .d(new_n226), .o1(new_n239));
  nano22aa1n03x5               g144(.a(new_n239), .b(new_n234), .c(new_n236), .out0(new_n240));
  norp02aa1n03x5               g145(.a(new_n237), .b(new_n240), .o1(\s[22] ));
  norp02aa1n06x5               g146(.a(new_n236), .b(new_n235), .o1(new_n242));
  norb02aa1n09x5               g147(.a(new_n242), .b(new_n226), .out0(new_n243));
  oao003aa1n06x5               g148(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .carry(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  aoi012aa1n02x5               g150(.a(new_n245), .b(new_n230), .c(new_n242), .o1(new_n246));
  inv040aa1n03x5               g151(.a(new_n246), .o1(new_n247));
  oaoi13aa1n06x5               g152(.a(new_n247), .b(new_n243), .c(new_n195), .d(new_n192), .o1(new_n248));
  xnrb03aa1n03x5               g153(.a(new_n248), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  tech160nm_fixnrc02aa1n04x5   g156(.a(\b[22] ), .b(\a[23] ), .out0(new_n252));
  tech160nm_fixnrc02aa1n04x5   g157(.a(\b[23] ), .b(\a[24] ), .out0(new_n253));
  oaoi13aa1n02x7               g158(.a(new_n253), .b(new_n251), .c(new_n248), .d(new_n252), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n243), .o1(new_n255));
  oaoi13aa1n04x5               g160(.a(new_n252), .b(new_n246), .c(new_n196), .d(new_n255), .o1(new_n256));
  nano22aa1n03x5               g161(.a(new_n256), .b(new_n251), .c(new_n253), .out0(new_n257));
  norp02aa1n03x5               g162(.a(new_n254), .b(new_n257), .o1(\s[24] ));
  norp02aa1n02x5               g163(.a(new_n253), .b(new_n252), .o1(new_n259));
  nano22aa1n02x4               g164(.a(new_n226), .b(new_n242), .c(new_n259), .out0(new_n260));
  oaih12aa1n02x5               g165(.a(new_n260), .b(new_n195), .c(new_n192), .o1(new_n261));
  inv000aa1n04x5               g166(.a(new_n229), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n242), .b(new_n262), .c(new_n225), .d(new_n215), .o1(new_n263));
  inv020aa1n02x5               g168(.a(new_n259), .o1(new_n264));
  oao003aa1n02x5               g169(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .carry(new_n265));
  aoai13aa1n12x5               g170(.a(new_n265), .b(new_n264), .c(new_n263), .d(new_n244), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnrc02aa1n12x5               g172(.a(\b[24] ), .b(\a[25] ), .out0(new_n268));
  xobna2aa1n03x5               g173(.a(new_n268), .b(new_n261), .c(new_n267), .out0(\s[25] ));
  oaoi13aa1n03x5               g174(.a(new_n266), .b(new_n260), .c(new_n195), .d(new_n192), .o1(new_n270));
  nor042aa1n03x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  tech160nm_fixnrc02aa1n04x5   g177(.a(\b[25] ), .b(\a[26] ), .out0(new_n273));
  oaoi13aa1n03x5               g178(.a(new_n273), .b(new_n272), .c(new_n270), .d(new_n268), .o1(new_n274));
  aoi012aa1n03x5               g179(.a(new_n268), .b(new_n261), .c(new_n267), .o1(new_n275));
  nano22aa1n03x5               g180(.a(new_n275), .b(new_n272), .c(new_n273), .out0(new_n276));
  norp02aa1n03x5               g181(.a(new_n274), .b(new_n276), .o1(\s[26] ));
  nor002aa1n03x5               g182(.a(new_n273), .b(new_n268), .o1(new_n278));
  nano32aa1n03x7               g183(.a(new_n226), .b(new_n278), .c(new_n242), .d(new_n259), .out0(new_n279));
  oai012aa1n12x5               g184(.a(new_n279), .b(new_n195), .c(new_n192), .o1(new_n280));
  oao003aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .c(new_n272), .carry(new_n281));
  aobi12aa1n12x5               g186(.a(new_n281), .b(new_n266), .c(new_n278), .out0(new_n282));
  xorc02aa1n02x5               g187(.a(\a[27] ), .b(\b[26] ), .out0(new_n283));
  xnbna2aa1n03x5               g188(.a(new_n283), .b(new_n282), .c(new_n280), .out0(\s[27] ));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  inv040aa1n03x5               g190(.a(new_n285), .o1(new_n286));
  nano23aa1n02x4               g191(.a(new_n176), .b(new_n183), .c(new_n184), .d(new_n177), .out0(new_n287));
  nano22aa1n02x4               g192(.a(new_n167), .b(new_n173), .c(new_n287), .out0(new_n288));
  aoai13aa1n02x5               g193(.a(new_n288), .b(new_n127), .c(new_n112), .d(new_n120), .o1(new_n289));
  aoai13aa1n02x7               g194(.a(new_n287), .b(new_n175), .c(new_n158), .d(new_n173), .o1(new_n290));
  nanp03aa1n03x5               g195(.a(new_n289), .b(new_n290), .c(new_n194), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n259), .b(new_n245), .c(new_n230), .d(new_n242), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n278), .o1(new_n293));
  aoai13aa1n04x5               g198(.a(new_n281), .b(new_n293), .c(new_n292), .d(new_n265), .o1(new_n294));
  aoai13aa1n06x5               g199(.a(new_n283), .b(new_n294), .c(new_n291), .d(new_n279), .o1(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  tech160nm_fiaoi012aa1n02p5x5 g201(.a(new_n296), .b(new_n295), .c(new_n286), .o1(new_n297));
  aobi12aa1n06x5               g202(.a(new_n283), .b(new_n282), .c(new_n280), .out0(new_n298));
  nano22aa1n03x7               g203(.a(new_n298), .b(new_n286), .c(new_n296), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[28] ));
  norb02aa1n02x5               g205(.a(new_n283), .b(new_n296), .out0(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n294), .c(new_n291), .d(new_n279), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n286), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  aoi012aa1n03x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  aobi12aa1n06x5               g210(.a(new_n301), .b(new_n282), .c(new_n280), .out0(new_n306));
  nano22aa1n03x7               g211(.a(new_n306), .b(new_n303), .c(new_n304), .out0(new_n307));
  norp02aa1n03x5               g212(.a(new_n305), .b(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g214(.a(new_n283), .b(new_n304), .c(new_n296), .out0(new_n310));
  aoai13aa1n06x5               g215(.a(new_n310), .b(new_n294), .c(new_n291), .d(new_n279), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[29] ), .b(\a[30] ), .out0(new_n313));
  aoi012aa1n02x5               g218(.a(new_n313), .b(new_n311), .c(new_n312), .o1(new_n314));
  aobi12aa1n06x5               g219(.a(new_n310), .b(new_n282), .c(new_n280), .out0(new_n315));
  nano22aa1n03x7               g220(.a(new_n315), .b(new_n312), .c(new_n313), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n314), .b(new_n316), .o1(\s[30] ));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n310), .b(new_n313), .out0(new_n319));
  aoai13aa1n02x5               g224(.a(new_n319), .b(new_n294), .c(new_n291), .d(new_n279), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n321));
  aoi012aa1n03x5               g226(.a(new_n318), .b(new_n320), .c(new_n321), .o1(new_n322));
  aobi12aa1n06x5               g227(.a(new_n319), .b(new_n282), .c(new_n280), .out0(new_n323));
  nano22aa1n03x7               g228(.a(new_n323), .b(new_n318), .c(new_n321), .out0(new_n324));
  norp02aa1n03x5               g229(.a(new_n322), .b(new_n324), .o1(\s[31] ));
  nanb02aa1n02x5               g230(.a(new_n108), .b(new_n109), .out0(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n326), .b(new_n132), .c(new_n105), .out0(\s[3] ));
  xorc02aa1n02x5               g232(.a(\a[4] ), .b(\b[3] ), .out0(new_n328));
  aoi112aa1n02x5               g233(.a(new_n328), .b(new_n108), .c(new_n133), .d(new_n132), .o1(new_n329));
  oaoi13aa1n02x5               g234(.a(new_n329), .b(new_n112), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g235(.a(new_n135), .b(\b[4] ), .c(new_n123), .out0(\s[5] ));
  oao003aa1n02x5               g236(.a(\a[5] ), .b(\b[4] ), .c(new_n135), .carry(new_n332));
  xnrb03aa1n02x5               g237(.a(new_n332), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g238(.a(\a[6] ), .b(\b[5] ), .c(new_n332), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g240(.a(new_n115), .b(new_n334), .c(new_n116), .o1(new_n336));
  xnrb03aa1n02x5               g241(.a(new_n336), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g242(.a(new_n129), .b(new_n165), .c(new_n126), .out0(\s[9] ));
endmodule


