// Benchmark "adder" written by ABC on Thu Jul 18 10:46:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n333, new_n334, new_n335, new_n336, new_n338,
    new_n339, new_n341, new_n342, new_n343, new_n345, new_n346, new_n348,
    new_n349, new_n350, new_n353;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1n08x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oao003aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .carry(new_n102));
  nor042aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor042aa1d18x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano23aa1n06x5               g011(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n107));
  inv000aa1n02x5               g012(.a(new_n105), .o1(new_n108));
  oaoi03aa1n12x5               g013(.a(\a[4] ), .b(\b[3] ), .c(new_n108), .o1(new_n109));
  inv040aa1d30x5               g014(.a(\a[6] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[5] ), .o1(new_n111));
  aoi022aa1n02x7               g016(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n112));
  oai122aa1n03x5               g017(.a(new_n112), .b(\a[7] ), .c(\b[6] ), .d(new_n110), .e(new_n111), .o1(new_n113));
  inv000aa1n15x5               g018(.a(\a[5] ), .o1(new_n114));
  inv020aa1n20x5               g019(.a(\b[4] ), .o1(new_n115));
  aboi22aa1d24x5               g020(.a(\b[5] ), .b(new_n110), .c(new_n114), .d(new_n115), .out0(new_n116));
  nor042aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand42aa1n06x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  norb02aa1n06x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  nano22aa1n03x7               g024(.a(new_n113), .b(new_n119), .c(new_n116), .out0(new_n120));
  aoai13aa1n06x5               g025(.a(new_n120), .b(new_n109), .c(new_n102), .d(new_n107), .o1(new_n121));
  inv000aa1d42x5               g026(.a(new_n116), .o1(new_n122));
  oai022aa1n02x5               g027(.a(new_n110), .b(new_n111), .c(\b[6] ), .d(\a[7] ), .o1(new_n123));
  nanp02aa1n03x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  norb02aa1n03x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  orn002aa1n02x5               g030(.a(\a[7] ), .b(\b[6] ), .o(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[8] ), .b(\b[7] ), .c(new_n126), .o1(new_n127));
  aoi013aa1n06x4               g032(.a(new_n127), .b(new_n125), .c(new_n119), .d(new_n122), .o1(new_n128));
  nand22aa1n06x5               g033(.a(new_n121), .b(new_n128), .o1(new_n129));
  tech160nm_finand02aa1n03p5x5 g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nanb02aa1n02x5               g035(.a(new_n97), .b(new_n130), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(new_n129), .b(new_n132), .o1(new_n133));
  nor022aa1n08x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nand42aa1n03x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n136), .b(new_n133), .c(new_n98), .out0(\s[10] ));
  nona22aa1n02x4               g042(.a(new_n129), .b(new_n131), .c(new_n136), .out0(new_n138));
  oaoi03aa1n12x5               g043(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nor042aa1n04x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nanp02aa1n04x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  norb02aa1n06x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  xnbna2aa1n03x5               g048(.a(new_n143), .b(new_n138), .c(new_n140), .out0(\s[11] ));
  aob012aa1n02x5               g049(.a(new_n143), .b(new_n138), .c(new_n140), .out0(new_n145));
  oai012aa1n02x5               g050(.a(new_n145), .b(\b[10] ), .c(\a[11] ), .o1(new_n146));
  nor042aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n03x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  aoib12aa1n02x5               g054(.a(new_n141), .b(new_n148), .c(new_n147), .out0(new_n150));
  aoi022aa1n02x5               g055(.a(new_n146), .b(new_n149), .c(new_n145), .d(new_n150), .o1(\s[12] ));
  nona23aa1n09x5               g056(.a(new_n135), .b(new_n130), .c(new_n97), .d(new_n134), .out0(new_n152));
  nano22aa1n12x5               g057(.a(new_n152), .b(new_n143), .c(new_n149), .out0(new_n153));
  nano23aa1n03x7               g058(.a(new_n141), .b(new_n147), .c(new_n148), .d(new_n142), .out0(new_n154));
  tech160nm_fiao0012aa1n02p5x5 g059(.a(new_n147), .b(new_n141), .c(new_n148), .o(new_n155));
  tech160nm_fiao0012aa1n02p5x5 g060(.a(new_n155), .b(new_n154), .c(new_n139), .o(new_n156));
  xnrc02aa1n12x5               g061(.a(\b[12] ), .b(\a[13] ), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n156), .c(new_n129), .d(new_n153), .o1(new_n159));
  aoi112aa1n02x5               g064(.a(new_n155), .b(new_n158), .c(new_n154), .d(new_n139), .o1(new_n160));
  aobi12aa1n02x5               g065(.a(new_n160), .b(new_n129), .c(new_n153), .out0(new_n161));
  norb02aa1n02x5               g066(.a(new_n159), .b(new_n161), .out0(\s[13] ));
  orn002aa1n02x5               g067(.a(\a[13] ), .b(\b[12] ), .o(new_n163));
  tech160nm_fixnrc02aa1n03p5x5 g068(.a(\b[13] ), .b(\a[14] ), .out0(new_n164));
  xobna2aa1n03x5               g069(.a(new_n164), .b(new_n159), .c(new_n163), .out0(\s[14] ));
  inv000aa1d42x5               g070(.a(new_n153), .o1(new_n166));
  nona32aa1n02x4               g071(.a(new_n129), .b(new_n164), .c(new_n157), .d(new_n166), .out0(new_n167));
  nor042aa1n06x5               g072(.a(new_n164), .b(new_n157), .o1(new_n168));
  aoai13aa1n12x5               g073(.a(new_n168), .b(new_n155), .c(new_n154), .d(new_n139), .o1(new_n169));
  oao003aa1n02x5               g074(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .carry(new_n170));
  and002aa1n02x5               g075(.a(new_n169), .b(new_n170), .o(new_n171));
  xorc02aa1n02x5               g076(.a(\a[15] ), .b(\b[14] ), .out0(new_n172));
  aob012aa1n06x5               g077(.a(new_n172), .b(new_n167), .c(new_n171), .out0(new_n173));
  nano22aa1n02x4               g078(.a(new_n172), .b(new_n169), .c(new_n170), .out0(new_n174));
  aobi12aa1n02x5               g079(.a(new_n173), .b(new_n174), .c(new_n167), .out0(\s[15] ));
  inv000aa1d42x5               g080(.a(\a[15] ), .o1(new_n176));
  oaib12aa1n02x5               g081(.a(new_n173), .b(\b[14] ), .c(new_n176), .out0(new_n177));
  xorc02aa1n02x5               g082(.a(\a[16] ), .b(\b[15] ), .out0(new_n178));
  aoib12aa1n02x5               g083(.a(new_n178), .b(new_n176), .c(\b[14] ), .out0(new_n179));
  aoi022aa1n02x5               g084(.a(new_n177), .b(new_n178), .c(new_n173), .d(new_n179), .o1(\s[16] ));
  inv040aa1d32x5               g085(.a(\a[16] ), .o1(new_n181));
  xroi22aa1d06x4               g086(.a(new_n176), .b(\b[14] ), .c(new_n181), .d(\b[15] ), .out0(new_n182));
  nand23aa1n03x5               g087(.a(new_n153), .b(new_n168), .c(new_n182), .o1(new_n183));
  inv020aa1n02x5               g088(.a(new_n183), .o1(new_n184));
  nand42aa1n06x5               g089(.a(new_n129), .b(new_n184), .o1(new_n185));
  aob012aa1n03x5               g090(.a(new_n182), .b(new_n169), .c(new_n170), .out0(new_n186));
  aoi112aa1n02x5               g091(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n187));
  aoib12aa1n09x5               g092(.a(new_n187), .b(new_n181), .c(\b[15] ), .out0(new_n188));
  nanp03aa1n06x5               g093(.a(new_n185), .b(new_n186), .c(new_n188), .o1(new_n189));
  tech160nm_fixorc02aa1n03p5x5 g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  nano22aa1n02x4               g095(.a(new_n190), .b(new_n186), .c(new_n188), .out0(new_n191));
  aoi022aa1n02x5               g096(.a(new_n191), .b(new_n185), .c(new_n189), .d(new_n190), .o1(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[17] ), .o1(new_n193));
  nanb02aa1n06x5               g098(.a(\b[16] ), .b(new_n193), .out0(new_n194));
  aoi012aa1n12x5               g099(.a(new_n183), .b(new_n121), .c(new_n128), .o1(new_n195));
  inv000aa1n02x5               g100(.a(new_n182), .o1(new_n196));
  aoai13aa1n12x5               g101(.a(new_n188), .b(new_n196), .c(new_n169), .d(new_n170), .o1(new_n197));
  tech160nm_fioai012aa1n05x5   g102(.a(new_n190), .b(new_n197), .c(new_n195), .o1(new_n198));
  xorc02aa1n02x5               g103(.a(\a[18] ), .b(\b[17] ), .out0(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n198), .c(new_n194), .out0(\s[18] ));
  inv000aa1d42x5               g105(.a(\a[18] ), .o1(new_n201));
  xroi22aa1d04x5               g106(.a(new_n193), .b(\b[16] ), .c(new_n201), .d(\b[17] ), .out0(new_n202));
  oai012aa1n03x5               g107(.a(new_n202), .b(new_n197), .c(new_n195), .o1(new_n203));
  norp02aa1n02x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  aoi112aa1n03x5               g109(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n205));
  nor002aa1n03x5               g110(.a(new_n205), .b(new_n204), .o1(new_n206));
  nor022aa1n16x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand02aa1n06x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n203), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fioaoi03aa1n04x5   g116(.a(\a[18] ), .b(\b[17] ), .c(new_n194), .o1(new_n212));
  aoai13aa1n03x5               g117(.a(new_n209), .b(new_n212), .c(new_n189), .d(new_n202), .o1(new_n213));
  inv040aa1n02x5               g118(.a(new_n207), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n209), .o1(new_n215));
  aoai13aa1n02x7               g120(.a(new_n214), .b(new_n215), .c(new_n203), .d(new_n206), .o1(new_n216));
  nor042aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1n06x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  aoib12aa1n02x5               g124(.a(new_n207), .b(new_n218), .c(new_n217), .out0(new_n220));
  aoi022aa1n02x7               g125(.a(new_n216), .b(new_n219), .c(new_n213), .d(new_n220), .o1(\s[20] ));
  nona23aa1n09x5               g126(.a(new_n218), .b(new_n208), .c(new_n207), .d(new_n217), .out0(new_n222));
  nano22aa1n02x5               g127(.a(new_n222), .b(new_n190), .c(new_n199), .out0(new_n223));
  tech160nm_fioai012aa1n05x5   g128(.a(new_n223), .b(new_n197), .c(new_n195), .o1(new_n224));
  oaoi03aa1n09x5               g129(.a(\a[20] ), .b(\b[19] ), .c(new_n214), .o1(new_n225));
  oabi12aa1n18x5               g130(.a(new_n225), .b(new_n222), .c(new_n206), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nand42aa1n04x5               g132(.a(new_n224), .b(new_n227), .o1(new_n228));
  xorc02aa1n02x5               g133(.a(\a[21] ), .b(\b[20] ), .out0(new_n229));
  nano23aa1n09x5               g134(.a(new_n207), .b(new_n217), .c(new_n218), .d(new_n208), .out0(new_n230));
  aoi112aa1n02x5               g135(.a(new_n225), .b(new_n229), .c(new_n230), .d(new_n212), .o1(new_n231));
  aoi022aa1n02x5               g136(.a(new_n228), .b(new_n229), .c(new_n224), .d(new_n231), .o1(\s[21] ));
  nand22aa1n03x5               g137(.a(new_n228), .b(new_n229), .o1(new_n233));
  nor002aa1d32x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n229), .o1(new_n236));
  aoai13aa1n02x5               g141(.a(new_n235), .b(new_n236), .c(new_n224), .d(new_n227), .o1(new_n237));
  xorc02aa1n02x5               g142(.a(\a[22] ), .b(\b[21] ), .out0(new_n238));
  norp02aa1n02x5               g143(.a(new_n238), .b(new_n234), .o1(new_n239));
  aoi022aa1n03x5               g144(.a(new_n237), .b(new_n238), .c(new_n233), .d(new_n239), .o1(\s[22] ));
  nanp02aa1n02x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  xnrc02aa1n02x5               g146(.a(\b[21] ), .b(\a[22] ), .out0(new_n242));
  nano22aa1n03x7               g147(.a(new_n242), .b(new_n235), .c(new_n241), .out0(new_n243));
  and003aa1n02x5               g148(.a(new_n202), .b(new_n243), .c(new_n230), .o(new_n244));
  tech160nm_fioai012aa1n05x5   g149(.a(new_n244), .b(new_n197), .c(new_n195), .o1(new_n245));
  oao003aa1n12x5               g150(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .carry(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aoi012aa1n02x5               g152(.a(new_n247), .b(new_n226), .c(new_n243), .o1(new_n248));
  nanp02aa1n06x5               g153(.a(new_n245), .b(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  aoi112aa1n02x5               g155(.a(new_n250), .b(new_n247), .c(new_n226), .d(new_n243), .o1(new_n251));
  aoi022aa1n02x5               g156(.a(new_n249), .b(new_n250), .c(new_n245), .d(new_n251), .o1(\s[23] ));
  nand22aa1n03x5               g157(.a(new_n249), .b(new_n250), .o1(new_n253));
  nor042aa1n06x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n250), .o1(new_n256));
  aoai13aa1n02x7               g161(.a(new_n255), .b(new_n256), .c(new_n245), .d(new_n248), .o1(new_n257));
  xorc02aa1n02x5               g162(.a(\a[24] ), .b(\b[23] ), .out0(new_n258));
  norp02aa1n02x5               g163(.a(new_n258), .b(new_n254), .o1(new_n259));
  aoi022aa1n03x5               g164(.a(new_n257), .b(new_n258), .c(new_n253), .d(new_n259), .o1(\s[24] ));
  and002aa1n12x5               g165(.a(new_n258), .b(new_n250), .o(new_n261));
  inv000aa1n09x5               g166(.a(new_n261), .o1(new_n262));
  nano32aa1n02x4               g167(.a(new_n262), .b(new_n202), .c(new_n230), .d(new_n243), .out0(new_n263));
  tech160nm_fioai012aa1n05x5   g168(.a(new_n263), .b(new_n197), .c(new_n195), .o1(new_n264));
  aoai13aa1n06x5               g169(.a(new_n243), .b(new_n225), .c(new_n230), .d(new_n212), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n255), .carry(new_n266));
  aoai13aa1n12x5               g171(.a(new_n266), .b(new_n262), .c(new_n265), .d(new_n246), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  nand42aa1n04x5               g173(.a(new_n264), .b(new_n268), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n261), .b(new_n247), .c(new_n226), .d(new_n243), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n270), .o1(new_n272));
  and003aa1n02x5               g177(.a(new_n271), .b(new_n272), .c(new_n266), .o(new_n273));
  aoi022aa1n02x5               g178(.a(new_n269), .b(new_n270), .c(new_n264), .d(new_n273), .o1(\s[25] ));
  nand22aa1n03x5               g179(.a(new_n269), .b(new_n270), .o1(new_n275));
  nor042aa1n03x5               g180(.a(\b[24] ), .b(\a[25] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoai13aa1n02x7               g182(.a(new_n277), .b(new_n272), .c(new_n264), .d(new_n268), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  norp02aa1n02x5               g184(.a(new_n279), .b(new_n276), .o1(new_n280));
  aoi022aa1n03x5               g185(.a(new_n278), .b(new_n279), .c(new_n275), .d(new_n280), .o1(\s[26] ));
  and002aa1n02x7               g186(.a(new_n279), .b(new_n270), .o(new_n282));
  inv000aa1n02x5               g187(.a(new_n282), .o1(new_n283));
  nano32aa1n06x5               g188(.a(new_n283), .b(new_n223), .c(new_n243), .d(new_n261), .out0(new_n284));
  tech160nm_fioai012aa1n05x5   g189(.a(new_n284), .b(new_n197), .c(new_n195), .o1(new_n285));
  oao003aa1n12x5               g190(.a(\a[26] ), .b(\b[25] ), .c(new_n277), .carry(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  aoi012aa1n06x5               g192(.a(new_n287), .b(new_n267), .c(new_n282), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(new_n288), .b(new_n285), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[27] ), .b(\b[26] ), .out0(new_n290));
  aoi112aa1n02x5               g195(.a(new_n290), .b(new_n287), .c(new_n267), .d(new_n282), .o1(new_n291));
  aoi022aa1n02x5               g196(.a(new_n289), .b(new_n290), .c(new_n285), .d(new_n291), .o1(\s[27] ));
  aoai13aa1n04x5               g197(.a(new_n286), .b(new_n283), .c(new_n271), .d(new_n266), .o1(new_n293));
  aoai13aa1n02x5               g198(.a(new_n290), .b(new_n293), .c(new_n189), .d(new_n284), .o1(new_n294));
  nor042aa1d18x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  inv000aa1n06x5               g200(.a(new_n295), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n290), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n296), .b(new_n297), .c(new_n288), .d(new_n285), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  norp02aa1n02x5               g204(.a(new_n299), .b(new_n295), .o1(new_n300));
  aoi022aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n294), .d(new_n300), .o1(\s[28] ));
  and002aa1n02x5               g206(.a(new_n299), .b(new_n290), .o(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n293), .c(new_n189), .d(new_n284), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n302), .o1(new_n304));
  oao003aa1n03x5               g209(.a(\a[28] ), .b(\b[27] ), .c(new_n296), .carry(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n304), .c(new_n288), .d(new_n285), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g215(.a(new_n297), .b(new_n299), .c(new_n307), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n293), .c(new_n189), .d(new_n284), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  tech160nm_fioaoi03aa1n02p5x5 g218(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n288), .d(new_n285), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .out0(new_n317));
  and002aa1n02x5               g222(.a(\b[28] ), .b(\a[29] ), .o(new_n318));
  oabi12aa1n02x5               g223(.a(new_n317), .b(\a[29] ), .c(\b[28] ), .out0(new_n319));
  oab012aa1n02x4               g224(.a(new_n319), .b(new_n305), .c(new_n318), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n316), .b(new_n317), .c(new_n312), .d(new_n320), .o1(\s[30] ));
  nano32aa1n06x5               g226(.a(new_n297), .b(new_n317), .c(new_n299), .d(new_n307), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n293), .c(new_n189), .d(new_n284), .o1(new_n323));
  inv000aa1d42x5               g228(.a(new_n322), .o1(new_n324));
  inv000aa1d42x5               g229(.a(\a[30] ), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[29] ), .o1(new_n326));
  oaoi03aa1n02x5               g231(.a(new_n325), .b(new_n326), .c(new_n314), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n324), .c(new_n288), .d(new_n285), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  oabi12aa1n02x5               g234(.a(new_n329), .b(\a[30] ), .c(\b[29] ), .out0(new_n330));
  oaoi13aa1n03x5               g235(.a(new_n330), .b(new_n314), .c(new_n325), .d(new_n326), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n328), .b(new_n329), .c(new_n323), .d(new_n331), .o1(\s[31] ));
  aoi022aa1n02x5               g237(.a(new_n100), .b(new_n99), .c(\a[1] ), .d(\b[0] ), .o1(new_n333));
  oaib12aa1n02x5               g238(.a(new_n333), .b(new_n100), .c(\a[2] ), .out0(new_n334));
  norb02aa1n02x5               g239(.a(new_n106), .b(new_n105), .out0(new_n335));
  aboi22aa1n03x5               g240(.a(new_n105), .b(new_n106), .c(new_n99), .d(new_n100), .out0(new_n336));
  aoi022aa1n02x5               g241(.a(new_n102), .b(new_n335), .c(new_n334), .d(new_n336), .o1(\s[3] ));
  norb02aa1n02x5               g242(.a(new_n104), .b(new_n103), .out0(new_n338));
  nanp02aa1n02x5               g243(.a(new_n102), .b(new_n335), .o1(new_n339));
  xnbna2aa1n03x5               g244(.a(new_n338), .b(new_n339), .c(new_n108), .out0(\s[4] ));
  xorc02aa1n02x5               g245(.a(\a[5] ), .b(\b[4] ), .out0(new_n341));
  aoai13aa1n02x5               g246(.a(new_n341), .b(new_n109), .c(new_n107), .d(new_n102), .o1(new_n342));
  aoi112aa1n02x5               g247(.a(new_n109), .b(new_n341), .c(new_n107), .d(new_n102), .o1(new_n343));
  norb02aa1n02x5               g248(.a(new_n342), .b(new_n343), .out0(\s[5] ));
  nanp02aa1n02x5               g249(.a(new_n115), .b(new_n114), .o1(new_n345));
  xorc02aa1n02x5               g250(.a(\a[6] ), .b(\b[5] ), .out0(new_n346));
  xnbna2aa1n03x5               g251(.a(new_n346), .b(new_n342), .c(new_n345), .out0(\s[6] ));
  aobi12aa1n02x5               g252(.a(new_n346), .b(new_n342), .c(new_n345), .out0(new_n348));
  aob012aa1n02x5               g253(.a(new_n125), .b(new_n342), .c(new_n116), .out0(new_n349));
  ao0022aa1n03x5               g254(.a(new_n126), .b(new_n124), .c(new_n110), .d(new_n111), .o(new_n350));
  oa0012aa1n02x5               g255(.a(new_n349), .b(new_n348), .c(new_n350), .o(\s[7] ));
  xnbna2aa1n03x5               g256(.a(new_n119), .b(new_n349), .c(new_n126), .out0(\s[8] ));
  aoi113aa1n02x5               g257(.a(new_n132), .b(new_n127), .c(new_n125), .d(new_n119), .e(new_n122), .o1(new_n353));
  aoi022aa1n02x5               g258(.a(new_n129), .b(new_n132), .c(new_n121), .d(new_n353), .o1(\s[9] ));
endmodule


