// Benchmark "adder" written by ABC on Thu Jul 18 08:58:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n185, new_n186, new_n187, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n310,
    new_n312, new_n314, new_n316, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nand42aa1n03x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1n03x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nanp02aa1n09x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor042aa1n03x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nand42aa1n04x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nano23aa1n03x5               g007(.a(new_n99), .b(new_n101), .c(new_n102), .d(new_n100), .out0(new_n103));
  nand42aa1n02x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  norp02aa1n04x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nor022aa1n06x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  oa0012aa1n03x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o(new_n107));
  oa0012aa1n02x5               g012(.a(new_n100), .b(new_n101), .c(new_n99), .o(new_n108));
  aoi012aa1n06x5               g013(.a(new_n108), .b(new_n103), .c(new_n107), .o1(new_n109));
  nor042aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  norb02aa1n06x4               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  nor042aa1n03x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  norb02aa1n02x7               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  and002aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o(new_n116));
  nor042aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  nand22aa1n09x5               g022(.a(\b[0] ), .b(\a[1] ), .o1(new_n118));
  oab012aa1n03x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .out0(new_n119));
  nand23aa1n04x5               g024(.a(new_n119), .b(new_n112), .c(new_n115), .o1(new_n120));
  tech160nm_fioai012aa1n03p5x5 g025(.a(new_n111), .b(new_n113), .c(new_n110), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  nano23aa1n02x5               g027(.a(new_n106), .b(new_n105), .c(new_n122), .d(new_n104), .out0(new_n123));
  nand02aa1n02x5               g028(.a(new_n123), .b(new_n103), .o1(new_n124));
  aoai13aa1n12x5               g029(.a(new_n109), .b(new_n124), .c(new_n120), .d(new_n121), .o1(new_n125));
  oa0012aa1n02x5               g030(.a(new_n97), .b(new_n125), .c(new_n98), .o(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand02aa1n03x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nor042aa1n03x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  nor002aa1n03x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  oaoi13aa1n04x5               g037(.a(new_n132), .b(new_n97), .c(new_n125), .d(new_n98), .o1(new_n133));
  nano22aa1n03x5               g038(.a(new_n133), .b(new_n128), .c(new_n131), .out0(new_n134));
  aoib12aa1n02x5               g039(.a(new_n131), .b(new_n128), .c(new_n133), .out0(new_n135));
  norp02aa1n02x5               g040(.a(new_n135), .b(new_n134), .o1(\s[11] ));
  nor042aa1n02x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand42aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(new_n139));
  oai012aa1n02x5               g044(.a(new_n139), .b(new_n134), .c(new_n129), .o1(new_n140));
  orn003aa1n03x7               g045(.a(new_n134), .b(new_n129), .c(new_n139), .o(new_n141));
  nanp02aa1n03x5               g046(.a(new_n141), .b(new_n140), .o1(\s[12] ));
  nano23aa1n06x5               g047(.a(new_n129), .b(new_n137), .c(new_n138), .d(new_n130), .out0(new_n143));
  oa0012aa1n06x5               g048(.a(new_n128), .b(new_n98), .c(new_n132), .o(new_n144));
  oa0012aa1n02x5               g049(.a(new_n138), .b(new_n137), .c(new_n129), .o(new_n145));
  aoi012aa1n12x5               g050(.a(new_n145), .b(new_n143), .c(new_n144), .o1(new_n146));
  nano23aa1n03x7               g051(.a(new_n98), .b(new_n132), .c(new_n128), .d(new_n97), .out0(new_n147));
  nanp02aa1n02x5               g052(.a(new_n147), .b(new_n143), .o1(new_n148));
  nanb02aa1n06x5               g053(.a(new_n148), .b(new_n125), .out0(new_n149));
  xorc02aa1n12x5               g054(.a(\a[13] ), .b(\b[12] ), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n149), .c(new_n146), .out0(\s[13] ));
  inv000aa1d42x5               g056(.a(\a[14] ), .o1(new_n152));
  nanp02aa1n03x5               g057(.a(new_n149), .b(new_n146), .o1(new_n153));
  nor042aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  tech160nm_fiaoi012aa1n05x5   g059(.a(new_n154), .b(new_n153), .c(new_n150), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(new_n152), .out0(\s[14] ));
  xnrc02aa1n02x5               g061(.a(\b[13] ), .b(\a[14] ), .out0(new_n157));
  nanb02aa1n02x5               g062(.a(new_n157), .b(new_n150), .out0(new_n158));
  inv000aa1d42x5               g063(.a(\b[13] ), .o1(new_n159));
  oaoi03aa1n02x5               g064(.a(new_n152), .b(new_n159), .c(new_n154), .o1(new_n160));
  aoai13aa1n04x5               g065(.a(new_n160), .b(new_n158), .c(new_n149), .d(new_n146), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  nor042aa1n02x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n163), .c(new_n161), .d(new_n165), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(new_n161), .b(new_n165), .o1(new_n170));
  nona22aa1n02x4               g075(.a(new_n170), .b(new_n168), .c(new_n163), .out0(new_n171));
  nanp02aa1n03x5               g076(.a(new_n171), .b(new_n169), .o1(\s[16] ));
  nano23aa1n06x5               g077(.a(new_n163), .b(new_n166), .c(new_n167), .d(new_n164), .out0(new_n173));
  oao003aa1n02x5               g078(.a(new_n152), .b(new_n159), .c(new_n154), .carry(new_n174));
  oai012aa1n02x5               g079(.a(new_n167), .b(new_n166), .c(new_n163), .o1(new_n175));
  aobi12aa1n06x5               g080(.a(new_n175), .b(new_n173), .c(new_n174), .out0(new_n176));
  inv000aa1n02x5               g081(.a(new_n176), .o1(new_n177));
  nanb03aa1n06x5               g082(.a(new_n157), .b(new_n173), .c(new_n150), .out0(new_n178));
  oab012aa1n12x5               g083(.a(new_n177), .b(new_n146), .c(new_n178), .out0(new_n179));
  nano32aa1n03x7               g084(.a(new_n158), .b(new_n173), .c(new_n143), .d(new_n147), .out0(new_n180));
  nand02aa1d10x5               g085(.a(new_n125), .b(new_n180), .o1(new_n181));
  xorc02aa1n02x5               g086(.a(\a[17] ), .b(\b[16] ), .out0(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n181), .c(new_n179), .out0(\s[17] ));
  inv000aa1d42x5               g088(.a(\a[18] ), .o1(new_n184));
  nanp02aa1n06x5               g089(.a(new_n181), .b(new_n179), .o1(new_n185));
  norp02aa1n04x5               g090(.a(\b[16] ), .b(\a[17] ), .o1(new_n186));
  tech160nm_fiaoi012aa1n05x5   g091(.a(new_n186), .b(new_n185), .c(new_n182), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[17] ), .c(new_n184), .out0(\s[18] ));
  oai012aa1n04x7               g093(.a(new_n176), .b(new_n146), .c(new_n178), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  xroi22aa1d04x5               g095(.a(new_n190), .b(\b[16] ), .c(new_n184), .d(\b[17] ), .out0(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n189), .c(new_n125), .d(new_n180), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[17] ), .o1(new_n193));
  oaoi03aa1n09x5               g098(.a(new_n184), .b(new_n193), .c(new_n186), .o1(new_n194));
  nor022aa1n08x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand22aa1n03x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nanb02aa1n02x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  xnbna2aa1n03x5               g103(.a(new_n198), .b(new_n192), .c(new_n194), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g105(.a(new_n192), .b(new_n194), .o1(new_n201));
  nor022aa1n06x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nanp02aa1n03x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  nanb02aa1n02x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  aoai13aa1n02x5               g109(.a(new_n204), .b(new_n195), .c(new_n201), .d(new_n198), .o1(new_n205));
  nanp02aa1n02x5               g110(.a(new_n201), .b(new_n198), .o1(new_n206));
  nona22aa1n02x4               g111(.a(new_n206), .b(new_n204), .c(new_n195), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n205), .o1(\s[20] ));
  nona23aa1n09x5               g113(.a(new_n203), .b(new_n196), .c(new_n195), .d(new_n202), .out0(new_n209));
  oa0012aa1n06x5               g114(.a(new_n203), .b(new_n202), .c(new_n195), .o(new_n210));
  inv030aa1n03x5               g115(.a(new_n210), .o1(new_n211));
  oai012aa1d24x5               g116(.a(new_n211), .b(new_n209), .c(new_n194), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  nano23aa1n06x5               g118(.a(new_n195), .b(new_n202), .c(new_n203), .d(new_n196), .out0(new_n214));
  nanp02aa1n02x5               g119(.a(new_n191), .b(new_n214), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n213), .b(new_n215), .c(new_n181), .d(new_n179), .o1(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  xorc02aa1n02x5               g123(.a(\a[21] ), .b(\b[20] ), .out0(new_n219));
  xorc02aa1n02x5               g124(.a(\a[22] ), .b(\b[21] ), .out0(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n218), .c(new_n216), .d(new_n219), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(new_n216), .b(new_n219), .o1(new_n223));
  nona22aa1n02x4               g128(.a(new_n223), .b(new_n221), .c(new_n218), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n224), .b(new_n222), .o1(\s[22] ));
  inv000aa1d42x5               g130(.a(\a[21] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d04x5               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(\b[21] ), .o1(new_n229));
  oao003aa1n02x5               g134(.a(new_n227), .b(new_n229), .c(new_n218), .carry(new_n230));
  aoi012aa1n02x5               g135(.a(new_n230), .b(new_n212), .c(new_n228), .o1(new_n231));
  nand03aa1n02x5               g136(.a(new_n228), .b(new_n191), .c(new_n214), .o1(new_n232));
  aoai13aa1n04x5               g137(.a(new_n231), .b(new_n232), .c(new_n181), .d(new_n179), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  xorc02aa1n12x5               g140(.a(\a[23] ), .b(\b[22] ), .out0(new_n236));
  xnrc02aa1n02x5               g141(.a(\b[23] ), .b(\a[24] ), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n235), .c(new_n233), .d(new_n236), .o1(new_n238));
  nanp02aa1n02x5               g143(.a(new_n233), .b(new_n236), .o1(new_n239));
  nona22aa1n02x4               g144(.a(new_n239), .b(new_n237), .c(new_n235), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[24] ));
  norb02aa1n02x5               g146(.a(new_n236), .b(new_n237), .out0(new_n242));
  nano22aa1n02x4               g147(.a(new_n215), .b(new_n242), .c(new_n228), .out0(new_n243));
  aoai13aa1n02x5               g148(.a(new_n243), .b(new_n189), .c(new_n125), .d(new_n180), .o1(new_n244));
  oao003aa1n02x5               g149(.a(new_n184), .b(new_n193), .c(new_n186), .carry(new_n245));
  aoai13aa1n06x5               g150(.a(new_n228), .b(new_n210), .c(new_n214), .d(new_n245), .o1(new_n246));
  inv000aa1n02x5               g151(.a(new_n230), .o1(new_n247));
  inv020aa1n02x5               g152(.a(new_n242), .o1(new_n248));
  orn002aa1n03x5               g153(.a(\a[23] ), .b(\b[22] ), .o(new_n249));
  oaoi03aa1n06x5               g154(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n02x5               g156(.a(new_n251), .b(new_n248), .c(new_n246), .d(new_n247), .o1(new_n252));
  nanb02aa1n03x5               g157(.a(new_n252), .b(new_n244), .out0(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g159(.a(\b[24] ), .b(\a[25] ), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[25] ), .b(\b[24] ), .out0(new_n256));
  nor002aa1n02x5               g161(.a(\b[25] ), .b(\a[26] ), .o1(new_n257));
  nand42aa1n06x5               g162(.a(\b[25] ), .b(\a[26] ), .o1(new_n258));
  norb02aa1n03x5               g163(.a(new_n258), .b(new_n257), .out0(new_n259));
  inv040aa1n03x5               g164(.a(new_n259), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n255), .c(new_n253), .d(new_n256), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n256), .b(new_n252), .c(new_n185), .d(new_n243), .o1(new_n262));
  nona22aa1n03x5               g167(.a(new_n262), .b(new_n260), .c(new_n255), .out0(new_n263));
  nanp02aa1n02x5               g168(.a(new_n261), .b(new_n263), .o1(\s[26] ));
  norb02aa1n09x5               g169(.a(new_n256), .b(new_n260), .out0(new_n265));
  nanp02aa1n02x5               g170(.a(new_n252), .b(new_n265), .o1(new_n266));
  oai012aa1n02x5               g171(.a(new_n258), .b(new_n257), .c(new_n255), .o1(new_n267));
  nano22aa1n03x5               g172(.a(new_n232), .b(new_n242), .c(new_n265), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n189), .c(new_n125), .d(new_n180), .o1(new_n269));
  nanp03aa1n06x5               g174(.a(new_n266), .b(new_n269), .c(new_n267), .o1(new_n270));
  xorb03aa1n02x5               g175(.a(new_n270), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[27] ), .b(\b[26] ), .out0(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[27] ), .b(\a[28] ), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n242), .b(new_n230), .c(new_n212), .d(new_n228), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n265), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n267), .b(new_n277), .c(new_n276), .d(new_n251), .o1(new_n278));
  aobi12aa1n12x5               g183(.a(new_n268), .b(new_n181), .c(new_n179), .out0(new_n279));
  oaih12aa1n02x5               g184(.a(new_n273), .b(new_n278), .c(new_n279), .o1(new_n280));
  nona22aa1n03x5               g185(.a(new_n280), .b(new_n274), .c(new_n272), .out0(new_n281));
  nanp02aa1n03x5               g186(.a(new_n275), .b(new_n281), .o1(\s[28] ));
  norb02aa1n02x5               g187(.a(new_n273), .b(new_n274), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n283), .b(new_n278), .c(new_n279), .o1(new_n284));
  inv000aa1n03x5               g189(.a(new_n272), .o1(new_n285));
  oaoi03aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .o1(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[28] ), .b(\a[29] ), .out0(new_n287));
  nona22aa1n03x5               g192(.a(new_n284), .b(new_n286), .c(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n287), .b(new_n286), .c(new_n270), .d(new_n283), .o1(new_n289));
  nanp02aa1n03x5               g194(.a(new_n289), .b(new_n288), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n118), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g196(.a(new_n273), .b(new_n287), .c(new_n274), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n293));
  oaoi03aa1n02x5               g198(.a(\a[29] ), .b(\b[28] ), .c(new_n293), .o1(new_n294));
  tech160nm_fixorc02aa1n03p5x5 g199(.a(\a[30] ), .b(\b[29] ), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n294), .c(new_n270), .d(new_n292), .o1(new_n297));
  oaih12aa1n02x5               g202(.a(new_n292), .b(new_n278), .c(new_n279), .o1(new_n298));
  nona22aa1n03x5               g203(.a(new_n298), .b(new_n294), .c(new_n296), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[30] ));
  nanp02aa1n02x5               g205(.a(new_n294), .b(new_n295), .o1(new_n301));
  oai012aa1n02x5               g206(.a(new_n301), .b(\b[29] ), .c(\a[30] ), .o1(new_n302));
  nano23aa1n02x4               g207(.a(new_n287), .b(new_n274), .c(new_n295), .d(new_n273), .out0(new_n303));
  oaih12aa1n02x5               g208(.a(new_n303), .b(new_n278), .c(new_n279), .o1(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[30] ), .b(\a[31] ), .out0(new_n305));
  nona22aa1n03x5               g210(.a(new_n304), .b(new_n305), .c(new_n302), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n305), .b(new_n302), .c(new_n270), .d(new_n303), .o1(new_n307));
  nanp02aa1n03x5               g212(.a(new_n307), .b(new_n306), .o1(\s[31] ));
  xorb03aa1n02x5               g213(.a(new_n119), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi012aa1n02x5               g214(.a(new_n113), .b(new_n119), .c(new_n115), .o1(new_n310));
  xnrc02aa1n02x5               g215(.a(new_n310), .b(new_n112), .out0(\s[4] ));
  nanp02aa1n02x5               g216(.a(new_n120), .b(new_n121), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g218(.a(new_n106), .b(new_n312), .c(new_n122), .o1(new_n314));
  xnrb03aa1n02x5               g219(.a(new_n314), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g220(.a(new_n107), .b(new_n312), .c(new_n123), .o(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g222(.a(new_n101), .b(new_n316), .c(new_n102), .o1(new_n318));
  xnrb03aa1n02x5               g223(.a(new_n318), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g224(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


