// Benchmark "adder" written by ABC on Thu Jul 18 04:18:56 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n346, new_n347, new_n348, new_n350, new_n351, new_n353,
    new_n355, new_n356, new_n357, new_n359, new_n360, new_n361, new_n362,
    new_n364, new_n366, new_n367, new_n368;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n04x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nona22aa1n09x5               g004(.a(new_n98), .b(new_n97), .c(new_n99), .out0(new_n100));
  inv000aa1d42x5               g005(.a(\a[4] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[3] ), .o1(new_n102));
  aoi022aa1n02x7               g007(.a(new_n102), .b(new_n101), .c(\a[2] ), .d(\b[1] ), .o1(new_n103));
  and002aa1n12x5               g008(.a(\b[2] ), .b(\a[3] ), .o(new_n104));
  nor042aa1d18x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  aoi112aa1n06x5               g010(.a(new_n104), .b(new_n105), .c(\a[4] ), .d(\b[3] ), .o1(new_n106));
  nand23aa1n04x5               g011(.a(new_n106), .b(new_n100), .c(new_n103), .o1(new_n107));
  tech160nm_fioaoi03aa1n03p5x5 g012(.a(new_n101), .b(new_n102), .c(new_n105), .o1(new_n108));
  nor002aa1d24x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1n06x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor002aa1d32x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nano23aa1n03x7               g017(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n113));
  nor002aa1n06x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  and002aa1n12x5               g019(.a(\b[5] ), .b(\a[6] ), .o(new_n115));
  nor042aa1n02x5               g020(.a(new_n115), .b(new_n114), .o1(new_n116));
  nand02aa1d04x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor042aa1n04x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  norb02aa1n03x5               g023(.a(new_n117), .b(new_n118), .out0(new_n119));
  nand23aa1n03x5               g024(.a(new_n113), .b(new_n116), .c(new_n119), .o1(new_n120));
  norb03aa1n03x4               g025(.a(new_n110), .b(new_n109), .c(new_n118), .out0(new_n121));
  aob012aa1n03x5               g026(.a(new_n117), .b(\b[5] ), .c(\a[6] ), .out0(new_n122));
  oab012aa1n02x5               g027(.a(new_n122), .b(new_n111), .c(new_n114), .out0(new_n123));
  aoi012aa1n02x7               g028(.a(new_n118), .b(new_n109), .c(new_n117), .o1(new_n124));
  aobi12aa1n06x5               g029(.a(new_n124), .b(new_n123), .c(new_n121), .out0(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n120), .c(new_n107), .d(new_n108), .o1(new_n126));
  nor022aa1n08x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  xnrc02aa1n12x5               g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .out0(new_n130));
  aoi112aa1n02x5               g035(.a(new_n127), .b(new_n130), .c(new_n126), .d(new_n129), .o1(new_n131));
  aoai13aa1n06x5               g036(.a(new_n130), .b(new_n127), .c(new_n126), .d(new_n129), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(\s[10] ));
  norp02aa1n02x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  oai012aa1n02x5               g040(.a(new_n135), .b(new_n134), .c(new_n127), .o1(new_n136));
  xorc02aa1n12x5               g041(.a(\a[11] ), .b(\b[10] ), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n132), .c(new_n136), .out0(\s[11] ));
  aob012aa1n03x5               g043(.a(new_n137), .b(new_n132), .c(new_n136), .out0(new_n139));
  tech160nm_fixnrc02aa1n04x5   g044(.a(\b[11] ), .b(\a[12] ), .out0(new_n140));
  nor002aa1n03x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norp02aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  and002aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o(new_n143));
  oab012aa1n02x4               g048(.a(new_n141), .b(new_n143), .c(new_n142), .out0(new_n144));
  inv000aa1n02x5               g049(.a(new_n141), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n137), .o1(new_n146));
  aoai13aa1n02x5               g051(.a(new_n145), .b(new_n146), .c(new_n132), .d(new_n136), .o1(new_n147));
  aboi22aa1n03x5               g052(.a(new_n140), .b(new_n147), .c(new_n139), .d(new_n144), .out0(\s[12] ));
  nona23aa1d24x5               g053(.a(new_n137), .b(new_n130), .c(new_n140), .d(new_n128), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoi112aa1n03x5               g055(.a(new_n143), .b(new_n142), .c(\a[11] ), .d(\b[10] ), .o1(new_n151));
  aoi012aa1n02x7               g056(.a(new_n141), .b(\a[10] ), .c(\b[9] ), .o1(new_n152));
  oai112aa1n04x5               g057(.a(new_n151), .b(new_n152), .c(new_n134), .d(new_n127), .o1(new_n153));
  oab012aa1n02x5               g058(.a(new_n142), .b(new_n145), .c(new_n143), .out0(new_n154));
  nand42aa1n02x5               g059(.a(new_n153), .b(new_n154), .o1(new_n155));
  tech160nm_fixnrc02aa1n04x5   g060(.a(\b[12] ), .b(\a[13] ), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n03x5               g062(.a(new_n157), .b(new_n155), .c(new_n126), .d(new_n150), .o1(new_n158));
  and003aa1n02x5               g063(.a(new_n153), .b(new_n156), .c(new_n154), .o(new_n159));
  aobi12aa1n02x5               g064(.a(new_n159), .b(new_n126), .c(new_n150), .out0(new_n160));
  norb02aa1n03x4               g065(.a(new_n158), .b(new_n160), .out0(\s[13] ));
  inv000aa1d42x5               g066(.a(\a[13] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(\b[12] ), .b(new_n162), .out0(new_n163));
  xorc02aa1n02x5               g068(.a(\a[14] ), .b(\b[13] ), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n158), .c(new_n163), .out0(\s[14] ));
  inv000aa1d42x5               g070(.a(\a[14] ), .o1(new_n166));
  xroi22aa1d06x4               g071(.a(new_n162), .b(\b[12] ), .c(new_n166), .d(\b[13] ), .out0(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n155), .c(new_n126), .d(new_n150), .o1(new_n168));
  oaoi03aa1n02x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  nor042aa1n12x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norb02aa1n06x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n168), .c(new_n170), .out0(\s[15] ));
  aob012aa1n03x5               g079(.a(new_n173), .b(new_n168), .c(new_n170), .out0(new_n175));
  xorc02aa1n02x5               g080(.a(\a[16] ), .b(\b[15] ), .out0(new_n176));
  inv040aa1d30x5               g081(.a(\a[16] ), .o1(new_n177));
  inv000aa1d42x5               g082(.a(\b[15] ), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(new_n178), .b(new_n177), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  aoi012aa1n02x5               g085(.a(new_n171), .b(new_n179), .c(new_n180), .o1(new_n181));
  inv030aa1n02x5               g086(.a(new_n171), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n173), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n168), .d(new_n170), .o1(new_n184));
  aoi022aa1n03x5               g089(.a(new_n184), .b(new_n176), .c(new_n175), .d(new_n181), .o1(\s[16] ));
  nano32aa1n03x7               g090(.a(new_n171), .b(new_n180), .c(new_n172), .d(new_n179), .out0(new_n186));
  nano22aa1d24x5               g091(.a(new_n149), .b(new_n167), .c(new_n186), .out0(new_n187));
  nand22aa1n12x5               g092(.a(new_n126), .b(new_n187), .o1(new_n188));
  nand22aa1n02x5               g093(.a(new_n167), .b(new_n186), .o1(new_n189));
  inv000aa1n02x5               g094(.a(new_n189), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(\b[13] ), .b(\a[14] ), .o1(new_n191));
  oai022aa1n02x5               g096(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n192));
  nand03aa1n02x5               g097(.a(new_n179), .b(new_n172), .c(new_n180), .o1(new_n193));
  nano32aa1n02x4               g098(.a(new_n193), .b(new_n192), .c(new_n182), .d(new_n191), .out0(new_n194));
  oaoi03aa1n02x5               g099(.a(new_n177), .b(new_n178), .c(new_n171), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aobi12aa1n12x5               g101(.a(new_n196), .b(new_n190), .c(new_n155), .out0(new_n197));
  nand02aa1d16x5               g102(.a(new_n197), .b(new_n188), .o1(new_n198));
  xorc02aa1n12x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  nona22aa1n02x4               g104(.a(new_n195), .b(new_n194), .c(new_n199), .out0(new_n200));
  aoi013aa1n02x4               g105(.a(new_n200), .b(new_n155), .c(new_n167), .d(new_n186), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n198), .b(new_n199), .c(new_n188), .d(new_n201), .o1(\s[17] ));
  nor002aa1d32x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n04x5               g109(.a(new_n196), .b(new_n189), .c(new_n153), .d(new_n154), .o1(new_n205));
  aoai13aa1n03x5               g110(.a(new_n199), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n206));
  nor042aa1n06x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nand02aa1d08x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  norb02aa1n06x4               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n206), .c(new_n204), .out0(\s[18] ));
  and002aa1n02x5               g115(.a(new_n199), .b(new_n209), .o(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n212));
  oaoi03aa1n02x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nor042aa1d18x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand02aa1n06x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n12x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n06x5               g124(.a(new_n217), .b(new_n213), .c(new_n198), .d(new_n211), .o1(new_n220));
  nor042aa1n09x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1d28x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  inv000aa1d42x5               g128(.a(\a[19] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\b[18] ), .o1(new_n225));
  aboi22aa1n03x5               g130(.a(new_n221), .b(new_n222), .c(new_n224), .d(new_n225), .out0(new_n226));
  inv040aa1n02x5               g131(.a(new_n215), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n217), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n227), .b(new_n228), .c(new_n212), .d(new_n214), .o1(new_n229));
  aoi022aa1n03x5               g134(.a(new_n229), .b(new_n223), .c(new_n220), .d(new_n226), .o1(\s[20] ));
  nano32aa1n03x7               g135(.a(new_n228), .b(new_n199), .c(new_n223), .d(new_n209), .out0(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n232));
  nanb03aa1n12x5               g137(.a(new_n221), .b(new_n222), .c(new_n216), .out0(new_n233));
  oai112aa1n06x5               g138(.a(new_n227), .b(new_n208), .c(new_n207), .d(new_n203), .o1(new_n234));
  aoi012aa1n12x5               g139(.a(new_n221), .b(new_n215), .c(new_n222), .o1(new_n235));
  oai012aa1d24x5               g140(.a(new_n235), .b(new_n234), .c(new_n233), .o1(new_n236));
  nor042aa1d18x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  nand02aa1n04x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  norb02aa1d27x5               g143(.a(new_n238), .b(new_n237), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n236), .c(new_n198), .d(new_n231), .o1(new_n240));
  nano22aa1n03x5               g145(.a(new_n221), .b(new_n216), .c(new_n222), .out0(new_n241));
  oai012aa1n02x5               g146(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .o1(new_n242));
  oab012aa1n03x5               g147(.a(new_n242), .b(new_n203), .c(new_n207), .out0(new_n243));
  inv020aa1n02x5               g148(.a(new_n235), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(new_n244), .b(new_n239), .c(new_n243), .d(new_n241), .o1(new_n245));
  aobi12aa1n02x7               g150(.a(new_n240), .b(new_n245), .c(new_n232), .out0(\s[21] ));
  nor042aa1n06x5               g151(.a(\b[21] ), .b(\a[22] ), .o1(new_n247));
  nand02aa1n08x5               g152(.a(\b[21] ), .b(\a[22] ), .o1(new_n248));
  norb02aa1n02x5               g153(.a(new_n248), .b(new_n247), .out0(new_n249));
  aoib12aa1n02x5               g154(.a(new_n237), .b(new_n248), .c(new_n247), .out0(new_n250));
  inv000aa1d42x5               g155(.a(new_n236), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n237), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n239), .o1(new_n253));
  aoai13aa1n02x7               g158(.a(new_n252), .b(new_n253), .c(new_n232), .d(new_n251), .o1(new_n254));
  aoi022aa1n03x5               g159(.a(new_n254), .b(new_n249), .c(new_n240), .d(new_n250), .o1(\s[22] ));
  inv020aa1n02x5               g160(.a(new_n231), .o1(new_n256));
  nano22aa1n06x5               g161(.a(new_n256), .b(new_n239), .c(new_n249), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n258));
  nano23aa1d15x5               g163(.a(new_n237), .b(new_n247), .c(new_n248), .d(new_n238), .out0(new_n259));
  aoi012aa1d24x5               g164(.a(new_n247), .b(new_n237), .c(new_n248), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  tech160nm_fiaoi012aa1n03p5x5 g166(.a(new_n261), .b(new_n236), .c(new_n259), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n263), .c(new_n198), .d(new_n257), .o1(new_n265));
  aoi112aa1n02x5               g170(.a(new_n264), .b(new_n261), .c(new_n236), .d(new_n259), .o1(new_n266));
  aobi12aa1n02x7               g171(.a(new_n265), .b(new_n266), .c(new_n258), .out0(\s[23] ));
  xorc02aa1n02x5               g172(.a(\a[24] ), .b(\b[23] ), .out0(new_n268));
  nor042aa1n06x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  norp02aa1n02x5               g174(.a(new_n268), .b(new_n269), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n269), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n264), .o1(new_n272));
  aoai13aa1n02x7               g177(.a(new_n271), .b(new_n272), .c(new_n258), .d(new_n262), .o1(new_n273));
  aoi022aa1n03x5               g178(.a(new_n273), .b(new_n268), .c(new_n265), .d(new_n270), .o1(\s[24] ));
  and002aa1n06x5               g179(.a(new_n268), .b(new_n264), .o(new_n275));
  nano22aa1n02x5               g180(.a(new_n256), .b(new_n275), .c(new_n259), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n259), .b(new_n244), .c(new_n243), .d(new_n241), .o1(new_n278));
  inv000aa1n06x5               g183(.a(new_n275), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[24] ), .b(\b[23] ), .c(new_n271), .carry(new_n280));
  aoai13aa1n12x5               g185(.a(new_n280), .b(new_n279), .c(new_n278), .d(new_n260), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n281), .c(new_n198), .d(new_n276), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n275), .b(new_n261), .c(new_n236), .d(new_n259), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n282), .o1(new_n285));
  and003aa1n02x5               g190(.a(new_n284), .b(new_n285), .c(new_n280), .o(new_n286));
  aobi12aa1n03x7               g191(.a(new_n283), .b(new_n286), .c(new_n277), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g192(.a(\a[26] ), .b(\b[25] ), .out0(new_n288));
  nor042aa1n03x5               g193(.a(\b[24] ), .b(\a[25] ), .o1(new_n289));
  norp02aa1n02x5               g194(.a(new_n288), .b(new_n289), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n281), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n289), .o1(new_n292));
  aoai13aa1n02x5               g197(.a(new_n292), .b(new_n285), .c(new_n277), .d(new_n291), .o1(new_n293));
  aoi022aa1n03x5               g198(.a(new_n293), .b(new_n288), .c(new_n283), .d(new_n290), .o1(\s[26] ));
  and002aa1n12x5               g199(.a(new_n288), .b(new_n282), .o(new_n295));
  nano32aa1n03x7               g200(.a(new_n256), .b(new_n295), .c(new_n259), .d(new_n275), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n205), .c(new_n126), .d(new_n187), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n295), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[26] ), .b(\b[25] ), .c(new_n292), .carry(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n298), .c(new_n284), .d(new_n280), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n300), .c(new_n198), .d(new_n296), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n299), .o1(new_n303));
  aoi112aa1n02x5               g208(.a(new_n301), .b(new_n303), .c(new_n281), .d(new_n295), .o1(new_n304));
  aobi12aa1n03x7               g209(.a(new_n302), .b(new_n304), .c(new_n297), .out0(\s[27] ));
  tech160nm_fixorc02aa1n02p5x5 g210(.a(\a[28] ), .b(\b[27] ), .out0(new_n306));
  norp02aa1n02x5               g211(.a(\b[26] ), .b(\a[27] ), .o1(new_n307));
  norp02aa1n02x5               g212(.a(new_n306), .b(new_n307), .o1(new_n308));
  tech160nm_fiaoi012aa1n05x5   g213(.a(new_n303), .b(new_n281), .c(new_n295), .o1(new_n309));
  inv000aa1n03x5               g214(.a(new_n307), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n301), .o1(new_n311));
  aoai13aa1n02x7               g216(.a(new_n310), .b(new_n311), .c(new_n309), .d(new_n297), .o1(new_n312));
  aoi022aa1n02x7               g217(.a(new_n312), .b(new_n306), .c(new_n302), .d(new_n308), .o1(\s[28] ));
  and002aa1n06x5               g218(.a(new_n306), .b(new_n301), .o(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n300), .c(new_n198), .d(new_n296), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n314), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[28] ), .b(\b[27] ), .c(new_n310), .carry(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n316), .c(new_n309), .d(new_n297), .o1(new_n318));
  xorc02aa1n03x5               g223(.a(\a[29] ), .b(\b[28] ), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n317), .b(new_n319), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n315), .d(new_n320), .o1(\s[29] ));
  xorb03aa1n02x5               g226(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d33x5               g227(.a(new_n311), .b(new_n306), .c(new_n319), .out0(new_n323));
  aoai13aa1n03x5               g228(.a(new_n323), .b(new_n300), .c(new_n198), .d(new_n296), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[28] ), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\a[29] ), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n317), .b(\b[28] ), .c(new_n327), .out0(new_n328));
  oaib12aa1n02x5               g233(.a(new_n328), .b(new_n326), .c(\a[29] ), .out0(new_n329));
  aoai13aa1n02x7               g234(.a(new_n329), .b(new_n325), .c(new_n309), .d(new_n297), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .out0(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n331), .b(new_n328), .c(new_n327), .d(new_n326), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n324), .d(new_n332), .o1(\s[30] ));
  nano32aa1n06x5               g238(.a(new_n311), .b(new_n331), .c(new_n306), .d(new_n319), .out0(new_n334));
  aoai13aa1n03x5               g239(.a(new_n334), .b(new_n300), .c(new_n198), .d(new_n296), .o1(new_n335));
  aoi022aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n336));
  norb02aa1n02x5               g241(.a(\b[30] ), .b(\a[31] ), .out0(new_n337));
  obai22aa1n02x7               g242(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n338));
  aoi112aa1n02x5               g243(.a(new_n338), .b(new_n337), .c(new_n328), .d(new_n336), .o1(new_n339));
  inv000aa1n02x5               g244(.a(new_n334), .o1(new_n340));
  norp02aa1n02x5               g245(.a(\b[29] ), .b(\a[30] ), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n341), .b(new_n328), .c(new_n336), .o1(new_n342));
  aoai13aa1n02x7               g247(.a(new_n342), .b(new_n340), .c(new_n309), .d(new_n297), .o1(new_n343));
  xorc02aa1n02x5               g248(.a(\a[31] ), .b(\b[30] ), .out0(new_n344));
  aoi022aa1n03x5               g249(.a(new_n343), .b(new_n344), .c(new_n335), .d(new_n339), .o1(\s[31] ));
  inv000aa1d42x5               g250(.a(new_n105), .o1(new_n346));
  nano32aa1n02x4               g251(.a(new_n104), .b(new_n100), .c(new_n98), .d(new_n346), .out0(new_n347));
  oai012aa1n02x5               g252(.a(new_n98), .b(new_n97), .c(new_n99), .o1(new_n348));
  oaoi13aa1n02x5               g253(.a(new_n347), .b(new_n348), .c(new_n104), .d(new_n105), .o1(\s[3] ));
  inv000aa1n03x5               g254(.a(new_n347), .o1(new_n350));
  xorc02aa1n02x5               g255(.a(\a[4] ), .b(\b[3] ), .out0(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n351), .b(new_n350), .c(new_n346), .out0(\s[4] ));
  norb02aa1n02x5               g257(.a(new_n112), .b(new_n111), .out0(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n353), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  inv000aa1d42x5               g259(.a(new_n111), .o1(new_n355));
  nanp02aa1n02x5               g260(.a(new_n107), .b(new_n108), .o1(new_n356));
  nanp02aa1n03x5               g261(.a(new_n356), .b(new_n353), .o1(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n116), .b(new_n357), .c(new_n355), .out0(\s[6] ));
  nona32aa1n02x4               g263(.a(new_n357), .b(new_n115), .c(new_n114), .d(new_n111), .out0(new_n359));
  nona23aa1n03x5               g264(.a(new_n359), .b(new_n110), .c(new_n109), .d(new_n115), .out0(new_n360));
  norb02aa1n02x5               g265(.a(new_n110), .b(new_n109), .out0(new_n361));
  aoib12aa1n02x5               g266(.a(new_n361), .b(new_n359), .c(new_n115), .out0(new_n362));
  norb02aa1n02x5               g267(.a(new_n360), .b(new_n362), .out0(\s[7] ));
  inv000aa1d42x5               g268(.a(new_n109), .o1(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n119), .b(new_n360), .c(new_n364), .out0(\s[8] ));
  nanb02aa1n02x5               g270(.a(new_n120), .b(new_n356), .out0(new_n366));
  nanp02aa1n02x5               g271(.a(new_n128), .b(new_n124), .o1(new_n367));
  aoi012aa1n02x5               g272(.a(new_n367), .b(new_n123), .c(new_n121), .o1(new_n368));
  aoi022aa1n02x5               g273(.a(new_n368), .b(new_n366), .c(new_n126), .d(new_n129), .o1(\s[9] ));
endmodule


