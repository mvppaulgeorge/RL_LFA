// Benchmark "adder" written by ABC on Thu Jul 18 01:00:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n335, new_n337, new_n338,
    new_n341, new_n342, new_n343, new_n345, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1n04x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  inv030aa1n02x5               g003(.a(new_n98), .o1(new_n99));
  nand22aa1n04x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n09x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n03x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  norp02aa1n24x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  tech160nm_finand02aa1n03p5x5 g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n02x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor042aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n06x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n03x4               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nand23aa1n03x5               g013(.a(new_n102), .b(new_n105), .c(new_n108), .o1(new_n109));
  inv040aa1d32x5               g014(.a(\a[3] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[2] ), .o1(new_n111));
  nanp02aa1n06x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  oaoi03aa1n03x5               g017(.a(\a[4] ), .b(\b[3] ), .c(new_n112), .o1(new_n113));
  inv000aa1n02x5               g018(.a(new_n113), .o1(new_n114));
  norp02aa1n12x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand22aa1n12x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  norb02aa1n02x7               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nor002aa1d32x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nand22aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  norb02aa1n03x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  nor042aa1n04x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nand42aa1n08x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  nor002aa1d32x5               g027(.a(\b[6] ), .b(\a[7] ), .o1(new_n123));
  nanp02aa1n12x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nano23aa1d15x5               g029(.a(new_n121), .b(new_n123), .c(new_n124), .d(new_n122), .out0(new_n125));
  nand23aa1n03x5               g030(.a(new_n125), .b(new_n117), .c(new_n120), .o1(new_n126));
  ao0012aa1n12x5               g031(.a(new_n115), .b(new_n118), .c(new_n116), .o(new_n127));
  inv000aa1n02x5               g032(.a(new_n123), .o1(new_n128));
  oaoi03aa1n12x5               g033(.a(\a[8] ), .b(\b[7] ), .c(new_n128), .o1(new_n129));
  aoi012aa1d24x5               g034(.a(new_n129), .b(new_n125), .c(new_n127), .o1(new_n130));
  aoai13aa1n12x5               g035(.a(new_n130), .b(new_n126), .c(new_n109), .d(new_n114), .o1(new_n131));
  nand42aa1n03x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  aoi012aa1n03x5               g037(.a(new_n97), .b(new_n131), .c(new_n132), .o1(new_n133));
  xnrb03aa1n03x5               g038(.a(new_n133), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n12x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nand02aa1d28x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  nano23aa1n06x5               g041(.a(new_n97), .b(new_n135), .c(new_n136), .d(new_n132), .out0(new_n137));
  aoi012aa1d24x5               g042(.a(new_n135), .b(new_n97), .c(new_n136), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nanp02aa1n09x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n139), .c(new_n131), .d(new_n137), .o1(new_n143));
  aoi112aa1n02x5               g048(.a(new_n142), .b(new_n139), .c(new_n131), .d(new_n137), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(\s[11] ));
  inv000aa1d42x5               g050(.a(new_n140), .o1(new_n146));
  nor002aa1d32x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand02aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  xnbna2aa1n03x5               g054(.a(new_n149), .b(new_n143), .c(new_n146), .out0(\s[12] ));
  nona23aa1d18x5               g055(.a(new_n148), .b(new_n141), .c(new_n140), .d(new_n147), .out0(new_n151));
  norb02aa1n02x5               g056(.a(new_n137), .b(new_n151), .out0(new_n152));
  tech160nm_fioai012aa1n03p5x5 g057(.a(new_n148), .b(new_n147), .c(new_n140), .o1(new_n153));
  oai012aa1n12x5               g058(.a(new_n153), .b(new_n151), .c(new_n138), .o1(new_n154));
  ao0012aa1n03x7               g059(.a(new_n154), .b(new_n131), .c(new_n152), .o(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  xnrc02aa1n12x5               g061(.a(\b[12] ), .b(\a[13] ), .out0(new_n157));
  nanb02aa1n06x5               g062(.a(new_n157), .b(new_n155), .out0(new_n158));
  oai012aa1n06x5               g063(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .o1(new_n159));
  tech160nm_fixnrc02aa1n05x5   g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  nor002aa1n04x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  aboi22aa1n03x5               g067(.a(new_n160), .b(new_n159), .c(new_n162), .d(new_n158), .out0(\s[14] ));
  nor042aa1n02x5               g068(.a(new_n160), .b(new_n157), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n154), .c(new_n131), .d(new_n152), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\a[14] ), .o1(new_n166));
  inv000aa1d42x5               g071(.a(\b[13] ), .o1(new_n167));
  tech160nm_fioaoi03aa1n03p5x5 g072(.a(new_n166), .b(new_n167), .c(new_n161), .o1(new_n168));
  nor002aa1d32x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nanp02aa1n04x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nanb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n165), .c(new_n168), .out0(\s[15] ));
  aob012aa1n03x5               g078(.a(new_n172), .b(new_n165), .c(new_n168), .out0(new_n174));
  inv000aa1d42x5               g079(.a(new_n169), .o1(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n171), .c(new_n165), .d(new_n168), .o1(new_n176));
  nor002aa1d32x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand02aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  aoib12aa1n02x5               g084(.a(new_n169), .b(new_n178), .c(new_n177), .out0(new_n180));
  aboi22aa1n03x5               g085(.a(new_n179), .b(new_n176), .c(new_n174), .d(new_n180), .out0(\s[16] ));
  tech160nm_fiaoi012aa1n05x5   g086(.a(new_n98), .b(new_n100), .c(new_n101), .o1(new_n182));
  nanb02aa1n03x5               g087(.a(new_n103), .b(new_n104), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n112), .b(new_n107), .o1(new_n184));
  norp03aa1n02x5               g089(.a(new_n182), .b(new_n183), .c(new_n184), .o1(new_n185));
  nona23aa1n03x5               g090(.a(new_n119), .b(new_n116), .c(new_n115), .d(new_n118), .out0(new_n186));
  norb02aa1n06x4               g091(.a(new_n122), .b(new_n121), .out0(new_n187));
  norb02aa1n06x5               g092(.a(new_n124), .b(new_n123), .out0(new_n188));
  nano22aa1n03x7               g093(.a(new_n186), .b(new_n187), .c(new_n188), .out0(new_n189));
  tech160nm_fioai012aa1n05x5   g094(.a(new_n189), .b(new_n185), .c(new_n113), .o1(new_n190));
  nona23aa1n09x5               g095(.a(new_n178), .b(new_n170), .c(new_n169), .d(new_n177), .out0(new_n191));
  nona23aa1n09x5               g096(.a(new_n164), .b(new_n137), .c(new_n191), .d(new_n151), .out0(new_n192));
  nor003aa1n02x5               g097(.a(new_n191), .b(new_n160), .c(new_n157), .o1(new_n193));
  oai012aa1n02x5               g098(.a(new_n178), .b(new_n177), .c(new_n169), .o1(new_n194));
  oai012aa1n02x5               g099(.a(new_n194), .b(new_n191), .c(new_n168), .o1(new_n195));
  aoi012aa1n06x5               g100(.a(new_n195), .b(new_n154), .c(new_n193), .o1(new_n196));
  aoai13aa1n12x5               g101(.a(new_n196), .b(new_n192), .c(new_n190), .d(new_n130), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g103(.a(\a[17] ), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\b[16] ), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(new_n200), .b(new_n199), .o1(new_n201));
  nano23aa1n02x4               g106(.a(new_n140), .b(new_n147), .c(new_n148), .d(new_n141), .out0(new_n202));
  nano23aa1n06x5               g107(.a(new_n169), .b(new_n177), .c(new_n178), .d(new_n170), .out0(new_n203));
  nona22aa1n02x4               g108(.a(new_n203), .b(new_n160), .c(new_n157), .out0(new_n204));
  nano22aa1n03x7               g109(.a(new_n204), .b(new_n137), .c(new_n202), .out0(new_n205));
  nand02aa1n02x5               g110(.a(new_n202), .b(new_n139), .o1(new_n206));
  oao003aa1n02x5               g111(.a(new_n166), .b(new_n167), .c(new_n161), .carry(new_n207));
  aobi12aa1n02x5               g112(.a(new_n194), .b(new_n203), .c(new_n207), .out0(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n204), .c(new_n206), .d(new_n153), .o1(new_n209));
  tech160nm_fixorc02aa1n03p5x5 g114(.a(\a[17] ), .b(\b[16] ), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n209), .c(new_n131), .d(new_n205), .o1(new_n211));
  nor002aa1n03x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nand42aa1n08x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  norb02aa1n06x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  xnbna2aa1n03x5               g119(.a(new_n214), .b(new_n211), .c(new_n201), .out0(\s[18] ));
  and002aa1n02x5               g120(.a(new_n210), .b(new_n214), .o(new_n216));
  oaoi03aa1n02x5               g121(.a(\a[18] ), .b(\b[17] ), .c(new_n201), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[19] ), .b(\b[18] ), .out0(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n217), .c(new_n197), .d(new_n216), .o1(new_n219));
  aoi112aa1n02x5               g124(.a(new_n218), .b(new_n217), .c(new_n197), .d(new_n216), .o1(new_n220));
  norb02aa1n03x4               g125(.a(new_n219), .b(new_n220), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  orn002aa1n24x5               g127(.a(\a[19] ), .b(\b[18] ), .o(new_n223));
  nanp02aa1n03x5               g128(.a(new_n219), .b(new_n223), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[20] ), .b(\b[19] ), .out0(new_n225));
  norb02aa1n02x5               g130(.a(new_n223), .b(new_n225), .out0(new_n226));
  aoi022aa1n02x7               g131(.a(new_n224), .b(new_n225), .c(new_n219), .d(new_n226), .o1(\s[20] ));
  xnrc02aa1n03x5               g132(.a(\b[19] ), .b(\a[20] ), .out0(new_n228));
  nano32aa1n02x4               g133(.a(new_n228), .b(new_n218), .c(new_n210), .d(new_n214), .out0(new_n229));
  aoi013aa1n02x4               g134(.a(new_n212), .b(new_n213), .c(new_n199), .d(new_n200), .o1(new_n230));
  tech160nm_fixnrc02aa1n02p5x5 g135(.a(\b[18] ), .b(\a[19] ), .out0(new_n231));
  oaoi03aa1n12x5               g136(.a(\a[20] ), .b(\b[19] ), .c(new_n223), .o1(new_n232));
  inv040aa1n03x5               g137(.a(new_n232), .o1(new_n233));
  oai013aa1n02x4               g138(.a(new_n233), .b(new_n230), .c(new_n231), .d(new_n228), .o1(new_n234));
  nor002aa1n16x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nand42aa1n08x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nanb02aa1n12x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n234), .c(new_n197), .d(new_n229), .o1(new_n239));
  nand03aa1n02x5               g144(.a(new_n217), .b(new_n218), .c(new_n225), .o1(new_n240));
  nona22aa1n02x4               g145(.a(new_n240), .b(new_n232), .c(new_n238), .out0(new_n241));
  aoi012aa1n02x5               g146(.a(new_n241), .b(new_n197), .c(new_n229), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n239), .b(new_n242), .out0(\s[21] ));
  tech160nm_fioai012aa1n04x5   g148(.a(new_n239), .b(\b[20] ), .c(\a[21] ), .o1(new_n244));
  nor022aa1n16x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  nand02aa1n08x5               g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  nanb02aa1n12x5               g151(.a(new_n245), .b(new_n246), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  aoib12aa1n02x5               g153(.a(new_n235), .b(new_n246), .c(new_n245), .out0(new_n249));
  aoi022aa1n02x7               g154(.a(new_n244), .b(new_n248), .c(new_n239), .d(new_n249), .o1(\s[22] ));
  nor002aa1n02x5               g155(.a(new_n228), .b(new_n231), .o1(new_n251));
  nona23aa1d18x5               g156(.a(new_n246), .b(new_n236), .c(new_n235), .d(new_n245), .out0(new_n252));
  nano32aa1n02x4               g157(.a(new_n252), .b(new_n251), .c(new_n214), .d(new_n210), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n209), .c(new_n131), .d(new_n205), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n252), .o1(new_n255));
  ao0012aa1n12x5               g160(.a(new_n245), .b(new_n235), .c(new_n246), .o(new_n256));
  aoi012aa1n02x5               g161(.a(new_n256), .b(new_n234), .c(new_n255), .o1(new_n257));
  xnrc02aa1n12x5               g162(.a(\b[22] ), .b(\a[23] ), .out0(new_n258));
  inv040aa1n02x5               g163(.a(new_n258), .o1(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n254), .c(new_n257), .out0(\s[23] ));
  aob012aa1n03x5               g165(.a(new_n259), .b(new_n254), .c(new_n257), .out0(new_n261));
  nor042aa1n06x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n03x5               g168(.a(new_n263), .b(new_n258), .c(new_n254), .d(new_n257), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[24] ), .b(\b[23] ), .out0(new_n265));
  norp02aa1n02x5               g170(.a(new_n265), .b(new_n262), .o1(new_n266));
  aoi022aa1n03x5               g171(.a(new_n264), .b(new_n265), .c(new_n261), .d(new_n266), .o1(\s[24] ));
  nona23aa1n09x5               g172(.a(new_n259), .b(new_n265), .c(new_n247), .d(new_n237), .out0(new_n268));
  nano32aa1n02x5               g173(.a(new_n268), .b(new_n251), .c(new_n214), .d(new_n210), .out0(new_n269));
  oaoi03aa1n02x5               g174(.a(\a[24] ), .b(\b[23] ), .c(new_n263), .o1(new_n270));
  aoi013aa1n06x4               g175(.a(new_n270), .b(new_n259), .c(new_n256), .d(new_n265), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n268), .c(new_n240), .d(new_n233), .o1(new_n272));
  xorc02aa1n12x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n272), .c(new_n197), .d(new_n269), .o1(new_n274));
  aoai13aa1n02x7               g179(.a(new_n269), .b(new_n209), .c(new_n131), .d(new_n205), .o1(new_n275));
  nor003aa1n02x5               g180(.a(new_n230), .b(new_n231), .c(new_n228), .o1(new_n276));
  norb03aa1n06x5               g181(.a(new_n265), .b(new_n252), .c(new_n258), .out0(new_n277));
  tech160nm_fioai012aa1n04x5   g182(.a(new_n277), .b(new_n276), .c(new_n232), .o1(new_n278));
  aoi113aa1n02x5               g183(.a(new_n273), .b(new_n270), .c(new_n259), .d(new_n256), .e(new_n265), .o1(new_n279));
  and003aa1n03x7               g184(.a(new_n275), .b(new_n279), .c(new_n278), .o(new_n280));
  norb02aa1n03x4               g185(.a(new_n274), .b(new_n280), .out0(\s[25] ));
  inv000aa1d42x5               g186(.a(\a[25] ), .o1(new_n282));
  oaib12aa1n03x5               g187(.a(new_n274), .b(\b[24] ), .c(new_n282), .out0(new_n283));
  tech160nm_fixorc02aa1n03p5x5 g188(.a(\a[26] ), .b(\b[25] ), .out0(new_n284));
  aoib12aa1n02x5               g189(.a(new_n284), .b(new_n282), .c(\b[24] ), .out0(new_n285));
  aoi022aa1n02x7               g190(.a(new_n283), .b(new_n284), .c(new_n274), .d(new_n285), .o1(\s[26] ));
  and002aa1n09x5               g191(.a(new_n284), .b(new_n273), .o(new_n287));
  nano32aa1n03x7               g192(.a(new_n268), .b(new_n287), .c(new_n216), .d(new_n251), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n209), .c(new_n131), .d(new_n205), .o1(new_n289));
  nanp02aa1n02x5               g194(.a(\b[25] ), .b(\a[26] ), .o1(new_n290));
  oai022aa1n02x5               g195(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n291));
  aoi022aa1n03x5               g196(.a(new_n272), .b(new_n287), .c(new_n290), .d(new_n291), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  xnbna2aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n292), .out0(\s[27] ));
  inv000aa1d42x5               g199(.a(new_n287), .o1(new_n295));
  nanp02aa1n02x5               g200(.a(new_n291), .b(new_n290), .o1(new_n296));
  aoai13aa1n12x5               g201(.a(new_n296), .b(new_n295), .c(new_n278), .d(new_n271), .o1(new_n297));
  aoai13aa1n06x5               g202(.a(new_n293), .b(new_n297), .c(new_n197), .d(new_n288), .o1(new_n298));
  inv000aa1d42x5               g203(.a(\a[27] ), .o1(new_n299));
  oaib12aa1n06x5               g204(.a(new_n298), .b(\b[26] ), .c(new_n299), .out0(new_n300));
  xorc02aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .out0(new_n301));
  norp02aa1n02x5               g206(.a(\b[26] ), .b(\a[27] ), .o1(new_n302));
  norp02aa1n02x5               g207(.a(new_n301), .b(new_n302), .o1(new_n303));
  aoi022aa1n03x5               g208(.a(new_n300), .b(new_n301), .c(new_n298), .d(new_n303), .o1(\s[28] ));
  inv000aa1d42x5               g209(.a(\a[28] ), .o1(new_n305));
  xroi22aa1d04x5               g210(.a(new_n299), .b(\b[26] ), .c(new_n305), .d(\b[27] ), .out0(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n297), .c(new_n197), .d(new_n288), .o1(new_n307));
  inv000aa1d42x5               g212(.a(\b[27] ), .o1(new_n308));
  oao003aa1n09x5               g213(.a(new_n305), .b(new_n308), .c(new_n302), .carry(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  nanp02aa1n03x5               g215(.a(new_n307), .b(new_n310), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norp02aa1n02x5               g217(.a(new_n309), .b(new_n312), .o1(new_n313));
  aoi022aa1n02x7               g218(.a(new_n311), .b(new_n312), .c(new_n307), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g220(.a(new_n293), .b(new_n312), .c(new_n301), .o(new_n316));
  aoai13aa1n06x5               g221(.a(new_n316), .b(new_n297), .c(new_n197), .d(new_n288), .o1(new_n317));
  inv000aa1d42x5               g222(.a(\a[29] ), .o1(new_n318));
  inv000aa1d42x5               g223(.a(\b[28] ), .o1(new_n319));
  oaoi03aa1n02x5               g224(.a(new_n318), .b(new_n319), .c(new_n309), .o1(new_n320));
  nanp02aa1n03x5               g225(.a(new_n317), .b(new_n320), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  oabi12aa1n02x5               g227(.a(new_n322), .b(\a[29] ), .c(\b[28] ), .out0(new_n323));
  oaoi13aa1n02x5               g228(.a(new_n323), .b(new_n309), .c(new_n318), .d(new_n319), .o1(new_n324));
  aoi022aa1n02x7               g229(.a(new_n321), .b(new_n322), .c(new_n317), .d(new_n324), .o1(\s[30] ));
  and003aa1n02x5               g230(.a(new_n306), .b(new_n322), .c(new_n312), .o(new_n326));
  aoai13aa1n02x7               g231(.a(new_n326), .b(new_n297), .c(new_n197), .d(new_n288), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n320), .carry(new_n328));
  nanb02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  nanb02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  aoi022aa1n03x5               g235(.a(new_n327), .b(new_n328), .c(new_n330), .d(new_n329), .o1(new_n331));
  aobi12aa1n03x5               g236(.a(new_n326), .b(new_n289), .c(new_n292), .out0(new_n332));
  nano32aa1n03x7               g237(.a(new_n332), .b(new_n330), .c(new_n328), .d(new_n329), .out0(new_n333));
  nor002aa1n02x5               g238(.a(new_n331), .b(new_n333), .o1(\s[31] ));
  aoi112aa1n02x5               g239(.a(new_n108), .b(new_n98), .c(new_n100), .d(new_n101), .o1(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n102), .c(new_n108), .o1(\s[3] ));
  oai013aa1n02x4               g241(.a(new_n114), .b(new_n182), .c(new_n183), .d(new_n184), .o1(new_n337));
  aoi112aa1n02x5               g242(.a(new_n106), .b(new_n105), .c(new_n102), .d(new_n107), .o1(new_n338));
  aoib12aa1n02x5               g243(.a(new_n338), .b(new_n337), .c(new_n103), .out0(\s[4] ));
  xnbna2aa1n03x5               g244(.a(new_n120), .b(new_n109), .c(new_n114), .out0(\s[5] ));
  aoi112aa1n02x5               g245(.a(new_n118), .b(new_n117), .c(new_n337), .d(new_n120), .o1(new_n341));
  inv000aa1d42x5               g246(.a(new_n127), .o1(new_n342));
  aoai13aa1n02x5               g247(.a(new_n342), .b(new_n186), .c(new_n109), .d(new_n114), .o1(new_n343));
  aoib12aa1n02x5               g248(.a(new_n341), .b(new_n343), .c(new_n115), .out0(\s[6] ));
  aoi113aa1n02x5               g249(.a(new_n188), .b(new_n127), .c(new_n337), .d(new_n117), .e(new_n120), .o1(new_n345));
  aoi012aa1n02x5               g250(.a(new_n345), .b(new_n188), .c(new_n343), .o1(\s[7] ));
  nanp02aa1n02x5               g251(.a(new_n343), .b(new_n188), .o1(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n187), .b(new_n347), .c(new_n128), .out0(\s[8] ));
  xorb03aa1n02x5               g253(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


