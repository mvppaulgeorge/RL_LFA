// Benchmark "adder" written by ABC on Wed Jul 17 13:53:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n337, new_n338,
    new_n339, new_n341, new_n342, new_n343, new_n344, new_n346, new_n347,
    new_n348, new_n350, new_n351, new_n353, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n08x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  orn002aa1n24x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nanp02aa1n06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n12x5               g005(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(new_n101));
  inv040aa1d32x5               g006(.a(\a[3] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[2] ), .o1(new_n103));
  nand22aa1n04x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand22aa1n04x5               g010(.a(new_n104), .b(new_n105), .o1(new_n106));
  aoi012aa1n02x5               g011(.a(new_n106), .b(new_n101), .c(new_n99), .o1(new_n107));
  oai022aa1n02x5               g012(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n108));
  norp02aa1n03x5               g013(.a(new_n107), .b(new_n108), .o1(new_n109));
  and002aa1n02x5               g014(.a(\b[4] ), .b(\a[5] ), .o(new_n110));
  oai022aa1d18x5               g015(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n111));
  nor042aa1n02x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[4] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[3] ), .o1(new_n114));
  oai022aa1n02x5               g019(.a(new_n113), .b(new_n114), .c(\b[7] ), .d(\a[8] ), .o1(new_n115));
  nand42aa1n03x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  tech160nm_fioai012aa1n04x5   g021(.a(new_n116), .b(\b[6] ), .c(\a[7] ), .o1(new_n117));
  aoi022aa1d24x5               g022(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n118));
  nona23aa1n02x4               g023(.a(new_n112), .b(new_n118), .c(new_n115), .d(new_n117), .out0(new_n119));
  norp02aa1n12x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  and002aa1n03x5               g025(.a(\b[6] ), .b(\a[7] ), .o(new_n121));
  aoi112aa1n03x5               g026(.a(new_n121), .b(new_n120), .c(\a[6] ), .d(\b[5] ), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .out0(new_n123));
  inv000aa1n02x5               g028(.a(new_n120), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n122), .c(new_n123), .d(new_n111), .o1(new_n126));
  oai012aa1n06x5               g031(.a(new_n126), .b(new_n109), .c(new_n119), .o1(new_n127));
  xnrc02aa1n12x5               g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(new_n127), .b(new_n129), .o1(new_n130));
  xnrc02aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  aoai13aa1n03x5               g038(.a(new_n132), .b(new_n97), .c(new_n127), .d(new_n129), .o1(new_n134));
  nand02aa1n04x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  oai022aa1d18x5               g040(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  nor002aa1d32x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nanp02aa1n12x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n06x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n134), .c(new_n137), .out0(\s[11] ));
  aob012aa1n03x5               g046(.a(new_n140), .b(new_n134), .c(new_n137), .out0(new_n142));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1d10x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  norp02aa1n02x5               g050(.a(new_n145), .b(new_n138), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n138), .o1(new_n147));
  inv000aa1d42x5               g052(.a(new_n140), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n147), .b(new_n148), .c(new_n134), .d(new_n137), .o1(new_n149));
  aoi022aa1n03x5               g054(.a(new_n149), .b(new_n145), .c(new_n142), .d(new_n146), .o1(\s[12] ));
  nona23aa1n02x4               g055(.a(new_n144), .b(new_n139), .c(new_n138), .d(new_n143), .out0(new_n151));
  nona32aa1n02x4               g056(.a(new_n127), .b(new_n151), .c(new_n131), .d(new_n128), .out0(new_n152));
  aboi22aa1n03x5               g057(.a(\b[3] ), .b(new_n113), .c(new_n102), .d(new_n103), .out0(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n106), .c(new_n101), .d(new_n99), .o1(new_n154));
  norb03aa1n03x4               g059(.a(new_n118), .b(new_n115), .c(new_n117), .out0(new_n155));
  nand23aa1n06x5               g060(.a(new_n154), .b(new_n112), .c(new_n155), .o1(new_n156));
  nano23aa1n02x4               g061(.a(new_n138), .b(new_n143), .c(new_n144), .d(new_n139), .out0(new_n157));
  nona22aa1n02x4               g062(.a(new_n157), .b(new_n131), .c(new_n128), .out0(new_n158));
  nanb03aa1n09x5               g063(.a(new_n143), .b(new_n144), .c(new_n139), .out0(new_n159));
  oai112aa1n06x5               g064(.a(new_n136), .b(new_n135), .c(\b[10] ), .d(\a[11] ), .o1(new_n160));
  aoi012aa1n12x5               g065(.a(new_n143), .b(new_n138), .c(new_n144), .o1(new_n161));
  oai012aa1d24x5               g066(.a(new_n161), .b(new_n160), .c(new_n159), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoai13aa1n04x5               g068(.a(new_n163), .b(new_n158), .c(new_n156), .d(new_n126), .o1(new_n164));
  nor022aa1n12x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand42aa1n06x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  oaib12aa1n02x5               g072(.a(new_n161), .b(new_n165), .c(new_n166), .out0(new_n168));
  oab012aa1n02x4               g073(.a(new_n168), .b(new_n160), .c(new_n159), .out0(new_n169));
  aoi022aa1n02x5               g074(.a(new_n164), .b(new_n167), .c(new_n152), .d(new_n169), .o1(\s[13] ));
  nor002aa1n06x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1n04x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(new_n165), .b(new_n173), .c(new_n164), .d(new_n167), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n173), .b(new_n165), .c(new_n164), .d(new_n166), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[14] ));
  nano23aa1n03x5               g081(.a(new_n165), .b(new_n171), .c(new_n172), .d(new_n166), .out0(new_n177));
  oa0012aa1n02x5               g082(.a(new_n172), .b(new_n171), .c(new_n165), .o(new_n178));
  nor042aa1n04x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nanp02aa1n02x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n178), .c(new_n164), .d(new_n177), .o1(new_n182));
  aoi112aa1n02x5               g087(.a(new_n181), .b(new_n178), .c(new_n164), .d(new_n177), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n182), .b(new_n183), .out0(\s[15] ));
  nor042aa1n04x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nand22aa1n02x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  norb02aa1n02x5               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  norp02aa1n02x5               g092(.a(new_n187), .b(new_n179), .o1(new_n188));
  tech160nm_fioai012aa1n03p5x5 g093(.a(new_n182), .b(\b[14] ), .c(\a[15] ), .o1(new_n189));
  aoi022aa1n02x5               g094(.a(new_n189), .b(new_n187), .c(new_n182), .d(new_n188), .o1(\s[16] ));
  nano32aa1n03x7               g095(.a(new_n158), .b(new_n187), .c(new_n177), .d(new_n181), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(new_n127), .b(new_n191), .o1(new_n192));
  nona23aa1n03x5               g097(.a(new_n172), .b(new_n166), .c(new_n165), .d(new_n171), .out0(new_n193));
  nona23aa1n03x5               g098(.a(new_n186), .b(new_n180), .c(new_n179), .d(new_n185), .out0(new_n194));
  nor042aa1n03x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  nona32aa1n03x5               g100(.a(new_n195), .b(new_n151), .c(new_n131), .d(new_n128), .out0(new_n196));
  nanb03aa1n02x5               g101(.a(new_n185), .b(new_n186), .c(new_n180), .out0(new_n197));
  oai122aa1n02x5               g102(.a(new_n172), .b(new_n171), .c(new_n165), .d(\b[14] ), .e(\a[15] ), .o1(new_n198));
  aoi012aa1n02x7               g103(.a(new_n185), .b(new_n179), .c(new_n186), .o1(new_n199));
  tech160nm_fioai012aa1n04x5   g104(.a(new_n199), .b(new_n198), .c(new_n197), .o1(new_n200));
  aoi012aa1n12x5               g105(.a(new_n200), .b(new_n162), .c(new_n195), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n201), .b(new_n196), .c(new_n156), .d(new_n126), .o1(new_n202));
  xorc02aa1n12x5               g107(.a(\a[17] ), .b(\b[16] ), .out0(new_n203));
  norp02aa1n02x5               g108(.a(new_n198), .b(new_n197), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n203), .b(new_n199), .out0(new_n205));
  aoi112aa1n02x5               g110(.a(new_n205), .b(new_n204), .c(new_n162), .d(new_n195), .o1(new_n206));
  aoi022aa1n02x5               g111(.a(new_n202), .b(new_n203), .c(new_n192), .d(new_n206), .o1(\s[17] ));
  nor022aa1n06x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  xorc02aa1n12x5               g113(.a(\a[18] ), .b(\b[17] ), .out0(new_n209));
  aoi112aa1n02x5               g114(.a(new_n208), .b(new_n209), .c(new_n202), .d(new_n203), .o1(new_n210));
  aoai13aa1n02x5               g115(.a(new_n209), .b(new_n208), .c(new_n202), .d(new_n203), .o1(new_n211));
  norb02aa1n02x5               g116(.a(new_n211), .b(new_n210), .out0(\s[18] ));
  inv000aa1n02x5               g117(.a(new_n200), .o1(new_n213));
  aob012aa1n03x5               g118(.a(new_n213), .b(new_n162), .c(new_n195), .out0(new_n214));
  and002aa1n12x5               g119(.a(new_n209), .b(new_n203), .o(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n214), .c(new_n127), .d(new_n191), .o1(new_n216));
  inv000aa1d42x5               g121(.a(\a[18] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[17] ), .o1(new_n218));
  oaoi03aa1n02x5               g123(.a(new_n217), .b(new_n218), .c(new_n208), .o1(new_n219));
  tech160nm_fixorc02aa1n04x5   g124(.a(\a[19] ), .b(\b[18] ), .out0(new_n220));
  xnbna2aa1n03x5               g125(.a(new_n220), .b(new_n216), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g127(.a(new_n220), .b(new_n216), .c(new_n219), .out0(new_n223));
  nor042aa1n03x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  and002aa1n12x5               g129(.a(\b[19] ), .b(\a[20] ), .o(new_n225));
  nor002aa1n03x5               g130(.a(new_n225), .b(new_n224), .o1(new_n226));
  norp02aa1n02x5               g131(.a(\b[18] ), .b(\a[19] ), .o1(new_n227));
  oab012aa1n02x4               g132(.a(new_n227), .b(new_n225), .c(new_n224), .out0(new_n228));
  aobi12aa1n03x5               g133(.a(new_n219), .b(new_n202), .c(new_n215), .out0(new_n229));
  oaoi03aa1n03x5               g134(.a(\a[19] ), .b(\b[18] ), .c(new_n229), .o1(new_n230));
  aoi022aa1n03x5               g135(.a(new_n230), .b(new_n226), .c(new_n223), .d(new_n228), .o1(\s[20] ));
  nanp03aa1d12x5               g136(.a(new_n215), .b(new_n220), .c(new_n226), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoi012aa1n02x5               g138(.a(new_n208), .b(new_n217), .c(new_n218), .o1(new_n234));
  aoi112aa1n03x4               g139(.a(new_n225), .b(new_n224), .c(\a[19] ), .d(\b[18] ), .o1(new_n235));
  oai022aa1n02x5               g140(.a(new_n217), .b(new_n218), .c(\b[18] ), .d(\a[19] ), .o1(new_n236));
  nona22aa1n03x5               g141(.a(new_n235), .b(new_n236), .c(new_n234), .out0(new_n237));
  aoib12aa1n06x5               g142(.a(new_n224), .b(new_n227), .c(new_n225), .out0(new_n238));
  nanp02aa1n02x5               g143(.a(new_n237), .b(new_n238), .o1(new_n239));
  xorc02aa1n12x5               g144(.a(\a[21] ), .b(\b[20] ), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n239), .c(new_n202), .d(new_n233), .o1(new_n241));
  nano22aa1n02x4               g146(.a(new_n240), .b(new_n237), .c(new_n238), .out0(new_n242));
  aobi12aa1n02x5               g147(.a(new_n242), .b(new_n202), .c(new_n233), .out0(new_n243));
  norb02aa1n02x5               g148(.a(new_n241), .b(new_n243), .out0(\s[21] ));
  xorc02aa1n12x5               g149(.a(\a[22] ), .b(\b[21] ), .out0(new_n245));
  nor042aa1n06x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  norp02aa1n02x5               g151(.a(new_n245), .b(new_n246), .o1(new_n247));
  inv000aa1d42x5               g152(.a(\a[21] ), .o1(new_n248));
  oaib12aa1n06x5               g153(.a(new_n241), .b(\b[20] ), .c(new_n248), .out0(new_n249));
  aoi022aa1n02x7               g154(.a(new_n249), .b(new_n245), .c(new_n241), .d(new_n247), .o1(\s[22] ));
  nand02aa1d12x5               g155(.a(new_n245), .b(new_n240), .o1(new_n251));
  nano32aa1n02x4               g156(.a(new_n251), .b(new_n215), .c(new_n220), .d(new_n226), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n246), .o1(new_n253));
  oao003aa1n02x5               g158(.a(\a[22] ), .b(\b[21] ), .c(new_n253), .carry(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n251), .c(new_n237), .d(new_n238), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n255), .c(new_n202), .d(new_n252), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n251), .o1(new_n258));
  nanb02aa1n02x5               g163(.a(new_n256), .b(new_n254), .out0(new_n259));
  aoi012aa1n02x5               g164(.a(new_n259), .b(new_n239), .c(new_n258), .o1(new_n260));
  aobi12aa1n02x5               g165(.a(new_n260), .b(new_n202), .c(new_n252), .out0(new_n261));
  norb02aa1n02x5               g166(.a(new_n257), .b(new_n261), .out0(\s[23] ));
  tech160nm_fixorc02aa1n03p5x5 g167(.a(\a[24] ), .b(\b[23] ), .out0(new_n263));
  norp02aa1n02x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  norp02aa1n02x5               g169(.a(new_n263), .b(new_n264), .o1(new_n265));
  tech160nm_fioai012aa1n03p5x5 g170(.a(new_n257), .b(\b[22] ), .c(\a[23] ), .o1(new_n266));
  aoi022aa1n02x7               g171(.a(new_n266), .b(new_n263), .c(new_n257), .d(new_n265), .o1(\s[24] ));
  and002aa1n02x7               g172(.a(new_n263), .b(new_n256), .o(new_n268));
  nona23aa1n06x5               g173(.a(new_n202), .b(new_n268), .c(new_n251), .d(new_n232), .out0(new_n269));
  aob012aa1n02x5               g174(.a(new_n264), .b(\b[23] ), .c(\a[24] ), .out0(new_n270));
  oai012aa1n02x5               g175(.a(new_n270), .b(\b[23] ), .c(\a[24] ), .o1(new_n271));
  aoi012aa1n02x5               g176(.a(new_n271), .b(new_n255), .c(new_n268), .o1(new_n272));
  tech160nm_fiaoi012aa1n02p5x5 g177(.a(new_n214), .b(new_n127), .c(new_n191), .o1(new_n273));
  nano32aa1n03x7               g178(.a(new_n273), .b(new_n268), .c(new_n233), .d(new_n258), .out0(new_n274));
  xorc02aa1n12x5               g179(.a(\a[25] ), .b(\b[24] ), .out0(new_n275));
  oaib12aa1n06x5               g180(.a(new_n275), .b(new_n274), .c(new_n272), .out0(new_n276));
  aoi112aa1n02x5               g181(.a(new_n275), .b(new_n271), .c(new_n255), .d(new_n268), .o1(new_n277));
  aobi12aa1n02x7               g182(.a(new_n276), .b(new_n277), .c(new_n269), .out0(\s[25] ));
  xorc02aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  nor042aa1n03x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n280), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n275), .o1(new_n283));
  aoai13aa1n04x5               g188(.a(new_n282), .b(new_n283), .c(new_n269), .d(new_n272), .o1(new_n284));
  aoi022aa1n03x5               g189(.a(new_n284), .b(new_n279), .c(new_n276), .d(new_n281), .o1(\s[26] ));
  and002aa1n02x5               g190(.a(new_n279), .b(new_n275), .o(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n271), .c(new_n255), .d(new_n268), .o1(new_n287));
  nano32aa1n03x7               g192(.a(new_n232), .b(new_n286), .c(new_n258), .d(new_n268), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n214), .c(new_n127), .d(new_n191), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[26] ), .b(\b[25] ), .c(new_n282), .carry(new_n290));
  nanp03aa1n06x5               g195(.a(new_n289), .b(new_n287), .c(new_n290), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n290), .o1(new_n293));
  aoi112aa1n02x5               g198(.a(new_n292), .b(new_n293), .c(new_n202), .d(new_n288), .o1(new_n294));
  aoi022aa1n02x5               g199(.a(new_n291), .b(new_n292), .c(new_n294), .d(new_n287), .o1(\s[27] ));
  nanp02aa1n03x5               g200(.a(new_n291), .b(new_n292), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .out0(new_n297));
  norp02aa1n02x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  norp02aa1n02x5               g203(.a(new_n297), .b(new_n298), .o1(new_n299));
  tech160nm_fiaoi012aa1n05x5   g204(.a(new_n293), .b(new_n202), .c(new_n288), .o1(new_n300));
  inv000aa1n03x5               g205(.a(new_n298), .o1(new_n301));
  inv030aa1n02x5               g206(.a(new_n292), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n301), .b(new_n302), .c(new_n300), .d(new_n287), .o1(new_n303));
  aoi022aa1n03x5               g208(.a(new_n303), .b(new_n297), .c(new_n296), .d(new_n299), .o1(\s[28] ));
  and002aa1n02x5               g209(.a(new_n297), .b(new_n292), .o(new_n305));
  nanp02aa1n03x5               g210(.a(new_n291), .b(new_n305), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  oao003aa1n02x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n301), .carry(new_n308));
  norb02aa1n02x5               g213(.a(new_n308), .b(new_n307), .out0(new_n309));
  inv000aa1d42x5               g214(.a(new_n305), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n308), .b(new_n310), .c(new_n300), .d(new_n287), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n311), .b(new_n307), .c(new_n306), .d(new_n309), .o1(\s[29] ));
  xorb03aa1n02x5               g217(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g218(.a(new_n297), .b(new_n292), .c(new_n307), .o1(new_n314));
  nanb02aa1n03x5               g219(.a(new_n314), .b(new_n291), .out0(new_n315));
  xorc02aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .out0(new_n316));
  inv000aa1d42x5               g221(.a(\a[29] ), .o1(new_n317));
  inv000aa1d42x5               g222(.a(\b[28] ), .o1(new_n318));
  oaib12aa1n02x5               g223(.a(new_n308), .b(\b[28] ), .c(new_n317), .out0(new_n319));
  oaoi13aa1n02x5               g224(.a(new_n316), .b(new_n319), .c(new_n317), .d(new_n318), .o1(new_n320));
  oaib12aa1n02x5               g225(.a(new_n319), .b(new_n318), .c(\a[29] ), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n314), .c(new_n300), .d(new_n287), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n322), .b(new_n316), .c(new_n315), .d(new_n320), .o1(\s[30] ));
  nano32aa1n02x4               g228(.a(new_n302), .b(new_n316), .c(new_n297), .d(new_n307), .out0(new_n324));
  nanp02aa1n03x5               g229(.a(new_n291), .b(new_n324), .o1(new_n325));
  aoi022aa1n02x5               g230(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n326));
  norb02aa1n02x5               g231(.a(\b[30] ), .b(\a[31] ), .out0(new_n327));
  obai22aa1n02x7               g232(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n328));
  aoi112aa1n02x5               g233(.a(new_n328), .b(new_n327), .c(new_n319), .d(new_n326), .o1(new_n329));
  inv000aa1n02x5               g234(.a(new_n324), .o1(new_n330));
  norp02aa1n02x5               g235(.a(\b[29] ), .b(\a[30] ), .o1(new_n331));
  aoi012aa1n02x5               g236(.a(new_n331), .b(new_n319), .c(new_n326), .o1(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n330), .c(new_n300), .d(new_n287), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  aoi022aa1n03x5               g239(.a(new_n333), .b(new_n334), .c(new_n329), .d(new_n325), .o1(\s[31] ));
  xobna2aa1n03x5               g240(.a(new_n106), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  aoai13aa1n02x5               g241(.a(new_n104), .b(new_n106), .c(new_n101), .d(new_n99), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[4] ), .b(\b[3] ), .out0(new_n338));
  norb02aa1n02x5               g243(.a(new_n104), .b(new_n338), .out0(new_n339));
  aboi22aa1n03x5               g244(.a(new_n107), .b(new_n339), .c(new_n337), .d(new_n338), .out0(\s[4] ));
  norp02aa1n02x5               g245(.a(\b[4] ), .b(\a[5] ), .o1(new_n341));
  aoi112aa1n02x5               g246(.a(new_n110), .b(new_n341), .c(\a[4] ), .d(\b[3] ), .o1(new_n342));
  oaib12aa1n02x5               g247(.a(new_n154), .b(new_n114), .c(\a[4] ), .out0(new_n343));
  xnrc02aa1n02x5               g248(.a(\b[4] ), .b(\a[5] ), .out0(new_n344));
  aoi022aa1n02x5               g249(.a(new_n343), .b(new_n344), .c(new_n342), .d(new_n154), .o1(\s[5] ));
  xorc02aa1n02x5               g250(.a(\a[6] ), .b(\b[5] ), .out0(new_n346));
  aoai13aa1n02x5               g251(.a(new_n346), .b(new_n341), .c(new_n154), .d(new_n342), .o1(new_n347));
  aoi112aa1n02x5               g252(.a(new_n341), .b(new_n346), .c(new_n154), .d(new_n342), .o1(new_n348));
  norb02aa1n02x5               g253(.a(new_n347), .b(new_n348), .out0(\s[6] ));
  orn002aa1n02x5               g254(.a(\a[6] ), .b(\b[5] ), .o(new_n350));
  norp02aa1n02x5               g255(.a(new_n121), .b(new_n120), .o1(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n351), .b(new_n347), .c(new_n350), .out0(\s[7] ));
  aob012aa1n02x5               g257(.a(new_n351), .b(new_n347), .c(new_n350), .out0(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n123), .b(new_n353), .c(new_n124), .out0(\s[8] ));
  aoi113aa1n02x5               g259(.a(new_n129), .b(new_n125), .c(new_n122), .d(new_n123), .e(new_n111), .o1(new_n355));
  aoi022aa1n02x5               g260(.a(new_n127), .b(new_n129), .c(new_n156), .d(new_n355), .o1(\s[9] ));
endmodule


