// Benchmark "adder" written by ABC on Thu Jul 18 01:36:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n323, new_n324,
    new_n327, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor042aa1d18x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  nor042aa1d18x5               g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  norp02aa1n24x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  inv000aa1n03x5               g010(.a(new_n105), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nanp02aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  norb02aa1n06x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nor042aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n09x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  norb02aa1n06x5               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  nona23aa1n03x5               g017(.a(new_n112), .b(new_n109), .c(new_n104), .d(new_n106), .out0(new_n113));
  oai012aa1n02x5               g018(.a(new_n108), .b(new_n110), .c(new_n107), .o1(new_n114));
  nand02aa1d04x5               g019(.a(new_n113), .b(new_n114), .o1(new_n115));
  nor002aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand22aa1n03x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  nand22aa1n02x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  aoi012aa1n06x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .o1(new_n119));
  nor002aa1d32x5               g024(.a(\b[3] ), .b(\a[4] ), .o1(new_n120));
  nanp02aa1n04x5               g025(.a(\b[3] ), .b(\a[4] ), .o1(new_n121));
  nor002aa1n12x5               g026(.a(\b[2] ), .b(\a[3] ), .o1(new_n122));
  nand02aa1n03x5               g027(.a(\b[2] ), .b(\a[3] ), .o1(new_n123));
  nona23aa1n09x5               g028(.a(new_n123), .b(new_n121), .c(new_n120), .d(new_n122), .out0(new_n124));
  tech160nm_fiaoi012aa1n03p5x5 g029(.a(new_n120), .b(new_n122), .c(new_n121), .o1(new_n125));
  oai012aa1n12x5               g030(.a(new_n125), .b(new_n124), .c(new_n119), .o1(new_n126));
  nand42aa1n03x5               g031(.a(\b[4] ), .b(\a[5] ), .o1(new_n127));
  nona23aa1n09x5               g032(.a(new_n105), .b(new_n127), .c(new_n103), .d(new_n102), .out0(new_n128));
  nano22aa1n06x5               g033(.a(new_n128), .b(new_n109), .c(new_n112), .out0(new_n129));
  nand02aa1n16x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n100), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n115), .c(new_n126), .d(new_n129), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n99), .b(new_n132), .c(new_n101), .out0(\s[10] ));
  inv000aa1d42x5               g038(.a(new_n104), .o1(new_n134));
  nano23aa1n02x4               g039(.a(new_n107), .b(new_n110), .c(new_n111), .d(new_n108), .out0(new_n135));
  oa0012aa1n02x5               g040(.a(new_n108), .b(new_n110), .c(new_n107), .o(new_n136));
  aoi013aa1n02x4               g041(.a(new_n136), .b(new_n135), .c(new_n105), .d(new_n134), .o1(new_n137));
  nand42aa1n02x5               g042(.a(new_n126), .b(new_n129), .o1(new_n138));
  nand42aa1n04x5               g043(.a(new_n138), .b(new_n137), .o1(new_n139));
  nanp03aa1n02x5               g044(.a(new_n139), .b(new_n99), .c(new_n131), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n97), .b(new_n100), .c(new_n98), .o1(new_n141));
  nor002aa1d24x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand02aa1d24x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  xobna2aa1n03x5               g049(.a(new_n144), .b(new_n140), .c(new_n141), .out0(\s[11] ));
  inv000aa1d42x5               g050(.a(new_n142), .o1(new_n146));
  aoai13aa1n03x5               g051(.a(new_n146), .b(new_n144), .c(new_n140), .d(new_n141), .o1(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nano23aa1d15x5               g053(.a(new_n97), .b(new_n100), .c(new_n130), .d(new_n98), .out0(new_n149));
  nor042aa1n03x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand42aa1n04x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nano23aa1n06x5               g056(.a(new_n142), .b(new_n150), .c(new_n151), .d(new_n143), .out0(new_n152));
  nand22aa1n12x5               g057(.a(new_n152), .b(new_n149), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n115), .c(new_n126), .d(new_n129), .o1(new_n155));
  aoi112aa1n06x5               g060(.a(new_n142), .b(new_n97), .c(new_n100), .d(new_n98), .o1(new_n156));
  aoi022aa1n06x5               g061(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n157));
  obai22aa1d24x5               g062(.a(new_n157), .b(new_n156), .c(\a[12] ), .d(\b[11] ), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  nor022aa1n08x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand42aa1n03x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  norb02aa1n03x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n155), .c(new_n159), .out0(\s[13] ));
  aoai13aa1n02x5               g068(.a(new_n159), .b(new_n153), .c(new_n138), .d(new_n137), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n160), .b(new_n164), .c(new_n161), .o1(new_n165));
  xnrb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand22aa1n03x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nona23aa1n03x5               g073(.a(new_n168), .b(new_n161), .c(new_n160), .d(new_n167), .out0(new_n169));
  aoi012aa1n02x7               g074(.a(new_n167), .b(new_n160), .c(new_n168), .o1(new_n170));
  aoai13aa1n03x5               g075(.a(new_n170), .b(new_n169), .c(new_n155), .d(new_n159), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n04x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n10x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nor002aa1n12x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand42aa1n03x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  norb02aa1n06x4               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  aoi112aa1n02x5               g082(.a(new_n173), .b(new_n177), .c(new_n171), .d(new_n174), .o1(new_n178));
  aoai13aa1n02x7               g083(.a(new_n177), .b(new_n173), .c(new_n171), .d(new_n174), .o1(new_n179));
  norb02aa1n02x7               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  xnrc02aa1n12x5               g085(.a(\b[16] ), .b(\a[17] ), .out0(new_n181));
  norb02aa1n03x5               g086(.a(new_n168), .b(new_n167), .out0(new_n182));
  nano23aa1n06x5               g087(.a(new_n173), .b(new_n175), .c(new_n176), .d(new_n174), .out0(new_n183));
  nano32aa1d12x5               g088(.a(new_n153), .b(new_n183), .c(new_n162), .d(new_n182), .out0(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n115), .c(new_n126), .d(new_n129), .o1(new_n185));
  inv000aa1n02x5               g090(.a(new_n173), .o1(new_n186));
  nano32aa1n03x7               g091(.a(new_n169), .b(new_n177), .c(new_n186), .d(new_n174), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n175), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(new_n176), .b(new_n174), .o1(new_n189));
  aoai13aa1n06x5               g094(.a(new_n188), .b(new_n189), .c(new_n170), .d(new_n186), .o1(new_n190));
  aoi012aa1d24x5               g095(.a(new_n190), .b(new_n158), .c(new_n187), .o1(new_n191));
  xobna2aa1n03x5               g096(.a(new_n181), .b(new_n185), .c(new_n191), .out0(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[18] ), .o1(new_n193));
  norp02aa1n02x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  nanp02aa1n09x5               g099(.a(new_n185), .b(new_n191), .o1(new_n195));
  aoib12aa1n06x5               g100(.a(new_n194), .b(new_n195), .c(new_n181), .out0(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  xnrc02aa1n02x5               g102(.a(\b[17] ), .b(\a[18] ), .out0(new_n198));
  nor042aa1n06x5               g103(.a(new_n198), .b(new_n181), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n199), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[17] ), .o1(new_n201));
  oao003aa1n02x5               g106(.a(new_n193), .b(new_n201), .c(new_n194), .carry(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  aoai13aa1n04x5               g108(.a(new_n203), .b(new_n200), .c(new_n185), .d(new_n191), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand42aa1n04x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nor042aa1n06x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand22aa1n09x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  aoi112aa1n02x5               g116(.a(new_n207), .b(new_n211), .c(new_n204), .d(new_n208), .o1(new_n212));
  aoai13aa1n03x5               g117(.a(new_n211), .b(new_n207), .c(new_n204), .d(new_n208), .o1(new_n213));
  norb02aa1n02x7               g118(.a(new_n213), .b(new_n212), .out0(\s[20] ));
  nanb03aa1n12x5               g119(.a(new_n209), .b(new_n210), .c(new_n208), .out0(new_n215));
  nona22aa1n02x4               g120(.a(new_n199), .b(new_n207), .c(new_n215), .out0(new_n216));
  oai022aa1d24x5               g121(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[18] ), .o1(new_n218));
  nanb02aa1n06x5               g123(.a(\a[19] ), .b(new_n218), .out0(new_n219));
  oai112aa1n06x5               g124(.a(new_n217), .b(new_n219), .c(new_n201), .d(new_n193), .o1(new_n220));
  aoi012aa1n12x5               g125(.a(new_n209), .b(new_n207), .c(new_n210), .o1(new_n221));
  oai012aa1d24x5               g126(.a(new_n221), .b(new_n220), .c(new_n215), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n04x5               g128(.a(new_n223), .b(new_n216), .c(new_n185), .d(new_n191), .o1(new_n224));
  xorb03aa1n02x5               g129(.a(new_n224), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  xnrc02aa1n12x5               g133(.a(\b[21] ), .b(\a[22] ), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoi112aa1n03x5               g135(.a(new_n226), .b(new_n230), .c(new_n224), .d(new_n228), .o1(new_n231));
  aoai13aa1n03x5               g136(.a(new_n230), .b(new_n226), .c(new_n224), .d(new_n228), .o1(new_n232));
  norb02aa1n02x7               g137(.a(new_n232), .b(new_n231), .out0(\s[22] ));
  nor042aa1n06x5               g138(.a(new_n229), .b(new_n227), .o1(new_n234));
  nona23aa1n09x5               g139(.a(new_n199), .b(new_n234), .c(new_n215), .d(new_n207), .out0(new_n235));
  inv000aa1d42x5               g140(.a(\a[22] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(\b[21] ), .o1(new_n237));
  oaoi03aa1n12x5               g142(.a(new_n236), .b(new_n237), .c(new_n226), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n222), .c(new_n234), .o1(new_n240));
  aoai13aa1n04x5               g145(.a(new_n240), .b(new_n235), .c(new_n185), .d(new_n191), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  tech160nm_fixorc02aa1n05x5   g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  xorc02aa1n02x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoi112aa1n02x7               g150(.a(new_n243), .b(new_n245), .c(new_n241), .d(new_n244), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n247));
  norb02aa1n02x7               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  nano22aa1n02x4               g153(.a(new_n209), .b(new_n208), .c(new_n210), .out0(new_n249));
  oai022aa1n02x5               g154(.a(new_n193), .b(new_n201), .c(\b[18] ), .d(\a[19] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n217), .b(new_n250), .out0(new_n251));
  inv040aa1n03x5               g156(.a(new_n221), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n234), .b(new_n252), .c(new_n251), .d(new_n249), .o1(new_n253));
  and002aa1n02x5               g158(.a(new_n245), .b(new_n244), .o(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  orn002aa1n02x5               g160(.a(\a[23] ), .b(\b[22] ), .o(new_n256));
  oao003aa1n02x5               g161(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .carry(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n255), .c(new_n253), .d(new_n238), .o1(new_n258));
  nano32aa1n02x5               g163(.a(new_n216), .b(new_n245), .c(new_n234), .d(new_n244), .out0(new_n259));
  xorc02aa1n06x5               g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n258), .c(new_n195), .d(new_n259), .o1(new_n261));
  aoi112aa1n02x5               g166(.a(new_n258), .b(new_n260), .c(new_n195), .d(new_n259), .o1(new_n262));
  norb02aa1n02x5               g167(.a(new_n261), .b(new_n262), .out0(\s[25] ));
  nor042aa1n03x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  tech160nm_fixorc02aa1n03p5x5 g169(.a(\a[26] ), .b(\b[25] ), .out0(new_n265));
  nona22aa1n02x5               g170(.a(new_n261), .b(new_n265), .c(new_n264), .out0(new_n266));
  inv040aa1n03x5               g171(.a(new_n264), .o1(new_n267));
  aobi12aa1n06x5               g172(.a(new_n265), .b(new_n261), .c(new_n267), .out0(new_n268));
  norb02aa1n03x4               g173(.a(new_n266), .b(new_n268), .out0(\s[26] ));
  inv000aa1n06x5               g174(.a(new_n191), .o1(new_n270));
  and002aa1n06x5               g175(.a(new_n265), .b(new_n260), .o(new_n271));
  nano22aa1n03x7               g176(.a(new_n235), .b(new_n254), .c(new_n271), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n270), .c(new_n139), .d(new_n184), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .c(new_n267), .carry(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  tech160nm_fiaoi012aa1n05x5   g180(.a(new_n275), .b(new_n258), .c(new_n271), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n276), .c(new_n273), .out0(\s[27] ));
  nor042aa1n03x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n277), .o1(new_n281));
  tech160nm_fiaoi012aa1n05x5   g186(.a(new_n281), .b(new_n276), .c(new_n273), .o1(new_n282));
  xnrc02aa1n12x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  nano22aa1n03x5               g188(.a(new_n282), .b(new_n280), .c(new_n283), .out0(new_n284));
  inv040aa1n03x5               g189(.a(new_n272), .o1(new_n285));
  aoi012aa1n06x5               g190(.a(new_n285), .b(new_n185), .c(new_n191), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n254), .b(new_n239), .c(new_n222), .d(new_n234), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n271), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n274), .b(new_n288), .c(new_n287), .d(new_n257), .o1(new_n289));
  oaih12aa1n02x5               g194(.a(new_n277), .b(new_n289), .c(new_n286), .o1(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n283), .b(new_n290), .c(new_n280), .o1(new_n291));
  norp02aa1n03x5               g196(.a(new_n291), .b(new_n284), .o1(\s[28] ));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  norb02aa1d21x5               g198(.a(new_n277), .b(new_n283), .out0(new_n294));
  oaih12aa1n02x5               g199(.a(new_n294), .b(new_n289), .c(new_n286), .o1(new_n295));
  oao003aa1n03x5               g200(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n296));
  tech160nm_fiaoi012aa1n02p5x5 g201(.a(new_n293), .b(new_n295), .c(new_n296), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n294), .o1(new_n298));
  aoi012aa1n06x5               g203(.a(new_n298), .b(new_n276), .c(new_n273), .o1(new_n299));
  nano22aa1n03x5               g204(.a(new_n299), .b(new_n293), .c(new_n296), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n297), .b(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g206(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g207(.a(\b[29] ), .b(\a[30] ), .out0(new_n303));
  norb03aa1n12x5               g208(.a(new_n277), .b(new_n293), .c(new_n283), .out0(new_n304));
  oaih12aa1n02x5               g209(.a(new_n304), .b(new_n289), .c(new_n286), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n306));
  tech160nm_fiaoi012aa1n05x5   g211(.a(new_n303), .b(new_n305), .c(new_n306), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n304), .o1(new_n308));
  tech160nm_fiaoi012aa1n04x5   g213(.a(new_n308), .b(new_n276), .c(new_n273), .o1(new_n309));
  nano22aa1n03x5               g214(.a(new_n309), .b(new_n303), .c(new_n306), .out0(new_n310));
  norp02aa1n03x5               g215(.a(new_n307), .b(new_n310), .o1(\s[30] ));
  norb02aa1n03x4               g216(.a(new_n304), .b(new_n303), .out0(new_n312));
  oaih12aa1n02x5               g217(.a(new_n312), .b(new_n289), .c(new_n286), .o1(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  tech160nm_fiaoi012aa1n02p5x5 g220(.a(new_n315), .b(new_n313), .c(new_n314), .o1(new_n316));
  inv000aa1n02x5               g221(.a(new_n312), .o1(new_n317));
  tech160nm_fiaoi012aa1n02p5x5 g222(.a(new_n317), .b(new_n276), .c(new_n273), .o1(new_n318));
  nano22aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n315), .out0(new_n319));
  norp02aa1n03x5               g224(.a(new_n316), .b(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g225(.a(new_n119), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g226(.a(new_n120), .o1(new_n322));
  nona22aa1n02x4               g227(.a(new_n123), .b(new_n119), .c(new_n122), .out0(new_n323));
  aoi012aa1n02x5               g228(.a(new_n122), .b(new_n322), .c(new_n121), .o1(new_n324));
  aoi022aa1n02x5               g229(.a(new_n126), .b(new_n322), .c(new_n323), .d(new_n324), .o1(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n126), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fiao0012aa1n02p5x5 g231(.a(new_n103), .b(new_n126), .c(new_n127), .o(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi012aa1n02x5               g233(.a(new_n102), .b(new_n327), .c(new_n105), .o1(new_n329));
  xnrc02aa1n02x5               g234(.a(new_n329), .b(new_n112), .out0(\s[7] ));
  oaoi03aa1n02x5               g235(.a(\a[7] ), .b(\b[6] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g237(.a(new_n131), .b(new_n138), .c(new_n137), .out0(\s[9] ));
endmodule


