// Benchmark "adder" written by ABC on Thu Jul 18 06:52:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n353, new_n354, new_n357, new_n359, new_n360, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[6] ), .b(\a[7] ), .o1(new_n97));
  inv030aa1n04x5               g002(.a(new_n97), .o1(new_n98));
  oaoi03aa1n02x5               g003(.a(\a[8] ), .b(\b[7] ), .c(new_n98), .o1(new_n99));
  nand22aa1n12x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor042aa1d18x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  norb02aa1n06x5               g006(.a(new_n100), .b(new_n101), .out0(new_n102));
  inv040aa1d32x5               g007(.a(\a[5] ), .o1(new_n103));
  inv030aa1d32x5               g008(.a(\b[4] ), .o1(new_n104));
  nand02aa1n04x5               g009(.a(new_n104), .b(new_n103), .o1(new_n105));
  oaoi03aa1n09x5               g010(.a(\a[6] ), .b(\b[5] ), .c(new_n105), .o1(new_n106));
  nand42aa1n16x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  norb02aa1n06x5               g012(.a(new_n107), .b(new_n97), .out0(new_n108));
  nanp03aa1n03x5               g013(.a(new_n106), .b(new_n102), .c(new_n108), .o1(new_n109));
  nanb02aa1n06x5               g014(.a(new_n99), .b(new_n109), .out0(new_n110));
  nor042aa1n04x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  nand22aa1n09x5               g016(.a(\b[0] ), .b(\a[1] ), .o1(new_n112));
  nand22aa1n09x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  aoi012aa1d24x5               g018(.a(new_n111), .b(new_n112), .c(new_n113), .o1(new_n114));
  nand02aa1n06x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  inv040aa1d32x5               g020(.a(\a[4] ), .o1(new_n116));
  inv040aa1d32x5               g021(.a(\b[3] ), .o1(new_n117));
  nand02aa1n08x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  nand02aa1n06x5               g023(.a(new_n118), .b(new_n115), .o1(new_n119));
  inv040aa1d32x5               g024(.a(\a[3] ), .o1(new_n120));
  inv040aa1d28x5               g025(.a(\b[2] ), .o1(new_n121));
  nand22aa1n04x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  nand02aa1d06x5               g027(.a(\b[2] ), .b(\a[3] ), .o1(new_n123));
  nand02aa1n06x5               g028(.a(new_n122), .b(new_n123), .o1(new_n124));
  nor042aa1d18x5               g029(.a(\b[2] ), .b(\a[3] ), .o1(new_n125));
  oaoi03aa1n09x5               g030(.a(new_n116), .b(new_n117), .c(new_n125), .o1(new_n126));
  oai013aa1n09x5               g031(.a(new_n126), .b(new_n114), .c(new_n119), .d(new_n124), .o1(new_n127));
  nanb02aa1n12x5               g032(.a(new_n101), .b(new_n100), .out0(new_n128));
  xnrc02aa1n12x5               g033(.a(\b[4] ), .b(\a[5] ), .out0(new_n129));
  nanp02aa1n06x5               g034(.a(\b[5] ), .b(\a[6] ), .o1(new_n130));
  nor022aa1n16x5               g035(.a(\b[5] ), .b(\a[6] ), .o1(new_n131));
  nona23aa1d18x5               g036(.a(new_n107), .b(new_n130), .c(new_n97), .d(new_n131), .out0(new_n132));
  nor043aa1d12x5               g037(.a(new_n132), .b(new_n129), .c(new_n128), .o1(new_n133));
  xorc02aa1n12x5               g038(.a(\a[9] ), .b(\b[8] ), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n134), .b(new_n110), .c(new_n127), .d(new_n133), .o1(new_n135));
  tech160nm_fioai012aa1n03p5x5 g040(.a(new_n135), .b(\b[8] ), .c(\a[9] ), .o1(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1d28x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  xnrc02aa1n12x5               g043(.a(\b[10] ), .b(\a[11] ), .out0(new_n139));
  oai122aa1n06x5               g044(.a(new_n135), .b(\b[9] ), .c(\a[10] ), .d(\b[8] ), .e(\a[9] ), .o1(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n139), .b(new_n140), .c(new_n138), .out0(\s[11] ));
  nor002aa1d24x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  xorc02aa1n02x5               g048(.a(\a[11] ), .b(\b[10] ), .out0(new_n144));
  nanp03aa1n02x5               g049(.a(new_n140), .b(new_n138), .c(new_n144), .o1(new_n145));
  nor042aa1n04x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nanp02aa1n12x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  aobi12aa1n02x7               g053(.a(new_n148), .b(new_n145), .c(new_n143), .out0(new_n149));
  aoi113aa1n02x5               g054(.a(new_n142), .b(new_n148), .c(new_n140), .d(new_n144), .e(new_n138), .o1(new_n150));
  nor002aa1n02x5               g055(.a(new_n149), .b(new_n150), .o1(\s[12] ));
  aoi013aa1n06x5               g056(.a(new_n99), .b(new_n106), .c(new_n108), .d(new_n102), .o1(new_n152));
  nor043aa1n03x5               g057(.a(new_n114), .b(new_n119), .c(new_n124), .o1(new_n153));
  inv030aa1n02x5               g058(.a(new_n126), .o1(new_n154));
  oai012aa1n06x5               g059(.a(new_n133), .b(new_n153), .c(new_n154), .o1(new_n155));
  nor042aa1n06x5               g060(.a(\b[9] ), .b(\a[10] ), .o1(new_n156));
  nano23aa1n02x5               g061(.a(new_n156), .b(new_n146), .c(new_n147), .d(new_n138), .out0(new_n157));
  nand23aa1n03x5               g062(.a(new_n157), .b(new_n134), .c(new_n144), .o1(new_n158));
  nor042aa1n02x5               g063(.a(new_n146), .b(new_n142), .o1(new_n159));
  oab012aa1n06x5               g064(.a(new_n156), .b(\a[9] ), .c(\b[8] ), .out0(new_n160));
  aob012aa1d18x5               g065(.a(new_n138), .b(\b[10] ), .c(\a[11] ), .out0(new_n161));
  oai012aa1n12x5               g066(.a(new_n159), .b(new_n160), .c(new_n161), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(new_n162), .b(new_n147), .o1(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n158), .c(new_n155), .d(new_n152), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  nand42aa1d28x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n166), .b(new_n164), .c(new_n167), .o1(new_n168));
  xnrb03aa1n03x5               g073(.a(new_n168), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nona23aa1n03x5               g074(.a(new_n147), .b(new_n138), .c(new_n156), .d(new_n146), .out0(new_n170));
  norb03aa1n03x5               g075(.a(new_n134), .b(new_n170), .c(new_n139), .out0(new_n171));
  aoai13aa1n03x5               g076(.a(new_n171), .b(new_n110), .c(new_n127), .d(new_n133), .o1(new_n172));
  nor002aa1d32x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nand42aa1n16x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nona23aa1n03x5               g079(.a(new_n174), .b(new_n167), .c(new_n166), .d(new_n173), .out0(new_n175));
  inv000aa1n02x5               g080(.a(new_n166), .o1(new_n176));
  oaoi03aa1n02x5               g081(.a(\a[14] ), .b(\b[13] ), .c(new_n176), .o1(new_n177));
  inv000aa1n02x5               g082(.a(new_n177), .o1(new_n178));
  aoai13aa1n03x5               g083(.a(new_n178), .b(new_n175), .c(new_n172), .d(new_n163), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n16x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  inv040aa1n02x5               g086(.a(new_n181), .o1(new_n182));
  nano23aa1d15x5               g087(.a(new_n166), .b(new_n173), .c(new_n174), .d(new_n167), .out0(new_n183));
  nand02aa1n08x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norb02aa1n09x5               g089(.a(new_n184), .b(new_n181), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n177), .c(new_n164), .d(new_n183), .o1(new_n186));
  nor042aa1n09x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nand02aa1d24x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  norb02aa1n15x5               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  inv040aa1n03x5               g094(.a(new_n189), .o1(new_n190));
  tech160nm_fiaoi012aa1n02p5x5 g095(.a(new_n190), .b(new_n186), .c(new_n182), .o1(new_n191));
  aoi112aa1n02x5               g096(.a(new_n181), .b(new_n189), .c(new_n179), .d(new_n184), .o1(new_n192));
  nor002aa1n02x5               g097(.a(new_n191), .b(new_n192), .o1(\s[16] ));
  nano32aa1n03x7               g098(.a(new_n190), .b(new_n182), .c(new_n184), .d(new_n147), .out0(new_n194));
  oai112aa1n04x5               g099(.a(new_n174), .b(new_n184), .c(new_n173), .d(new_n166), .o1(new_n195));
  nor042aa1n02x5               g100(.a(new_n187), .b(new_n181), .o1(new_n196));
  aoi022aa1n06x5               g101(.a(new_n195), .b(new_n196), .c(\b[15] ), .d(\a[16] ), .o1(new_n197));
  aoi013aa1n09x5               g102(.a(new_n197), .b(new_n194), .c(new_n162), .d(new_n183), .o1(new_n198));
  nano22aa1n02x4               g103(.a(new_n175), .b(new_n185), .c(new_n189), .out0(new_n199));
  nand02aa1n02x5               g104(.a(new_n171), .b(new_n199), .o1(new_n200));
  aoai13aa1n12x5               g105(.a(new_n198), .b(new_n200), .c(new_n155), .d(new_n152), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  inv000aa1n06x5               g108(.a(new_n203), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n123), .b(new_n125), .out0(new_n205));
  nona22aa1n03x5               g110(.a(new_n205), .b(new_n114), .c(new_n119), .out0(new_n206));
  nano23aa1n02x4               g111(.a(new_n97), .b(new_n131), .c(new_n107), .d(new_n130), .out0(new_n207));
  nona22aa1n02x4               g112(.a(new_n207), .b(new_n129), .c(new_n128), .out0(new_n208));
  aoai13aa1n06x5               g113(.a(new_n152), .b(new_n208), .c(new_n206), .d(new_n126), .o1(new_n209));
  nanp03aa1n02x5               g114(.a(new_n194), .b(new_n162), .c(new_n183), .o1(new_n210));
  nanb02aa1n02x5               g115(.a(new_n197), .b(new_n210), .out0(new_n211));
  nano32aa1n03x7               g116(.a(new_n158), .b(new_n189), .c(new_n183), .d(new_n185), .out0(new_n212));
  xorc02aa1n12x5               g117(.a(\a[17] ), .b(\b[16] ), .out0(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n211), .c(new_n209), .d(new_n212), .o1(new_n214));
  nor042aa1n09x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  nanp02aa1n04x5               g120(.a(\b[17] ), .b(\a[18] ), .o1(new_n216));
  nanb02aa1n02x5               g121(.a(new_n215), .b(new_n216), .out0(new_n217));
  xobna2aa1n03x5               g122(.a(new_n217), .b(new_n214), .c(new_n204), .out0(\s[18] ));
  aoai13aa1n06x5               g123(.a(new_n212), .b(new_n110), .c(new_n133), .d(new_n127), .o1(new_n219));
  inv040aa1d30x5               g124(.a(\a[17] ), .o1(new_n220));
  inv020aa1n04x5               g125(.a(\a[18] ), .o1(new_n221));
  xroi22aa1d06x4               g126(.a(new_n220), .b(\b[16] ), .c(new_n221), .d(\b[17] ), .out0(new_n222));
  inv000aa1n02x5               g127(.a(new_n222), .o1(new_n223));
  oaoi03aa1n02x5               g128(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n224));
  inv000aa1n02x5               g129(.a(new_n224), .o1(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n223), .c(new_n219), .d(new_n198), .o1(new_n226));
  xorb03aa1n02x5               g131(.a(new_n226), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g132(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g133(.a(\b[18] ), .b(\a[19] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  nand42aa1n16x5               g135(.a(\b[18] ), .b(\a[19] ), .o1(new_n231));
  nanb02aa1d24x5               g136(.a(new_n229), .b(new_n231), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n02x7               g138(.a(new_n233), .b(new_n224), .c(new_n201), .d(new_n222), .o1(new_n234));
  tech160nm_fixnrc02aa1n04x5   g139(.a(\b[19] ), .b(\a[20] ), .out0(new_n235));
  aoi012aa1n03x5               g140(.a(new_n235), .b(new_n234), .c(new_n230), .o1(new_n236));
  inv030aa1n02x5               g141(.a(new_n235), .o1(new_n237));
  aoi112aa1n03x4               g142(.a(new_n229), .b(new_n237), .c(new_n226), .d(new_n231), .o1(new_n238));
  norp02aa1n03x5               g143(.a(new_n236), .b(new_n238), .o1(\s[20] ));
  nona23aa1d18x5               g144(.a(new_n237), .b(new_n213), .c(new_n217), .d(new_n232), .out0(new_n240));
  oab012aa1n06x5               g145(.a(new_n229), .b(\a[20] ), .c(\b[19] ), .out0(new_n241));
  oai112aa1n06x5               g146(.a(new_n216), .b(new_n231), .c(new_n215), .d(new_n203), .o1(new_n242));
  aoi022aa1d18x5               g147(.a(new_n242), .b(new_n241), .c(\a[20] ), .d(\b[19] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n240), .c(new_n219), .d(new_n198), .o1(new_n245));
  xorb03aa1n02x5               g150(.a(new_n245), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g151(.a(\b[20] ), .b(\a[21] ), .o1(new_n247));
  inv040aa1n02x5               g152(.a(new_n247), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n240), .o1(new_n249));
  nand42aa1n03x5               g154(.a(\b[20] ), .b(\a[21] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n250), .b(new_n247), .out0(new_n251));
  aoai13aa1n02x7               g156(.a(new_n251), .b(new_n243), .c(new_n201), .d(new_n249), .o1(new_n252));
  inv040aa1d32x5               g157(.a(\a[22] ), .o1(new_n253));
  inv040aa1d28x5               g158(.a(\b[21] ), .o1(new_n254));
  nand22aa1n09x5               g159(.a(new_n254), .b(new_n253), .o1(new_n255));
  nand02aa1n08x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  nand22aa1n12x5               g161(.a(new_n255), .b(new_n256), .o1(new_n257));
  aoi012aa1n03x5               g162(.a(new_n257), .b(new_n252), .c(new_n248), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n257), .o1(new_n259));
  aoi112aa1n03x4               g164(.a(new_n247), .b(new_n259), .c(new_n245), .d(new_n251), .o1(new_n260));
  norp02aa1n03x5               g165(.a(new_n258), .b(new_n260), .o1(\s[22] ));
  nano22aa1n03x7               g166(.a(new_n257), .b(new_n248), .c(new_n250), .out0(new_n262));
  nona23aa1d18x5               g167(.a(new_n222), .b(new_n262), .c(new_n235), .d(new_n232), .out0(new_n263));
  nand02aa1d06x5               g168(.a(new_n242), .b(new_n241), .o1(new_n264));
  nanp02aa1n02x5               g169(.a(\b[19] ), .b(\a[20] ), .o1(new_n265));
  nano32aa1n03x7               g170(.a(new_n257), .b(new_n248), .c(new_n250), .d(new_n265), .out0(new_n266));
  oaoi03aa1n09x5               g171(.a(new_n253), .b(new_n254), .c(new_n247), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  aoi012aa1n12x5               g173(.a(new_n268), .b(new_n264), .c(new_n266), .o1(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n263), .c(new_n219), .d(new_n198), .o1(new_n270));
  xorb03aa1n02x5               g175(.a(new_n270), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g176(.a(\b[22] ), .b(\a[23] ), .o1(new_n272));
  inv000aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  inv040aa1n06x5               g178(.a(new_n263), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n269), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[23] ), .b(\b[22] ), .out0(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n275), .c(new_n201), .d(new_n274), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[24] ), .b(\b[23] ), .out0(new_n278));
  aobi12aa1n02x5               g183(.a(new_n278), .b(new_n277), .c(new_n273), .out0(new_n279));
  aoi112aa1n03x4               g184(.a(new_n272), .b(new_n278), .c(new_n270), .d(new_n276), .o1(new_n280));
  norp02aa1n03x5               g185(.a(new_n279), .b(new_n280), .o1(\s[24] ));
  nano32aa1n03x7               g186(.a(new_n240), .b(new_n278), .c(new_n262), .d(new_n276), .out0(new_n282));
  inv000aa1n02x5               g187(.a(new_n282), .o1(new_n283));
  inv020aa1n02x5               g188(.a(new_n241), .o1(new_n284));
  norp02aa1n02x5               g189(.a(new_n215), .b(new_n203), .o1(new_n285));
  nano22aa1n02x4               g190(.a(new_n285), .b(new_n216), .c(new_n231), .out0(new_n286));
  oai012aa1n06x5               g191(.a(new_n266), .b(new_n286), .c(new_n284), .o1(new_n287));
  nand02aa1d04x5               g192(.a(new_n278), .b(new_n276), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[24] ), .b(\b[23] ), .c(new_n273), .carry(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n288), .c(new_n287), .d(new_n267), .o1(new_n290));
  inv000aa1n02x5               g195(.a(new_n290), .o1(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n283), .c(new_n219), .d(new_n198), .o1(new_n292));
  xorb03aa1n02x5               g197(.a(new_n292), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n06x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  inv000aa1n02x5               g199(.a(new_n294), .o1(new_n295));
  xorc02aa1n03x5               g200(.a(\a[25] ), .b(\b[24] ), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n290), .c(new_n201), .d(new_n282), .o1(new_n297));
  xorc02aa1n03x5               g202(.a(\a[26] ), .b(\b[25] ), .out0(new_n298));
  aobi12aa1n02x5               g203(.a(new_n298), .b(new_n297), .c(new_n295), .out0(new_n299));
  aoi112aa1n03x4               g204(.a(new_n294), .b(new_n298), .c(new_n292), .d(new_n296), .o1(new_n300));
  norp02aa1n03x5               g205(.a(new_n299), .b(new_n300), .o1(\s[26] ));
  inv000aa1n02x5               g206(.a(new_n288), .o1(new_n302));
  and002aa1n06x5               g207(.a(new_n298), .b(new_n296), .o(new_n303));
  nano22aa1d15x5               g208(.a(new_n263), .b(new_n302), .c(new_n303), .out0(new_n304));
  aoai13aa1n06x5               g209(.a(new_n304), .b(new_n211), .c(new_n209), .d(new_n212), .o1(new_n305));
  oao003aa1n06x5               g210(.a(\a[26] ), .b(\b[25] ), .c(new_n295), .carry(new_n306));
  inv000aa1n02x5               g211(.a(new_n306), .o1(new_n307));
  aoi012aa1n06x5               g212(.a(new_n307), .b(new_n290), .c(new_n303), .o1(new_n308));
  xorc02aa1n12x5               g213(.a(\a[27] ), .b(\b[26] ), .out0(new_n309));
  xnbna2aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n308), .out0(\s[27] ));
  nor042aa1n03x5               g215(.a(\b[26] ), .b(\a[27] ), .o1(new_n311));
  inv040aa1n03x5               g216(.a(new_n311), .o1(new_n312));
  aoai13aa1n06x5               g217(.a(new_n302), .b(new_n268), .c(new_n264), .d(new_n266), .o1(new_n313));
  inv000aa1n02x5               g218(.a(new_n303), .o1(new_n314));
  aoai13aa1n12x5               g219(.a(new_n306), .b(new_n314), .c(new_n313), .d(new_n289), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n309), .b(new_n315), .c(new_n201), .d(new_n304), .o1(new_n316));
  xnrc02aa1n12x5               g221(.a(\b[27] ), .b(\a[28] ), .out0(new_n317));
  aoi012aa1n02x7               g222(.a(new_n317), .b(new_n316), .c(new_n312), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n309), .o1(new_n319));
  tech160nm_fiaoi012aa1n02p5x5 g224(.a(new_n319), .b(new_n305), .c(new_n308), .o1(new_n320));
  nano22aa1n03x5               g225(.a(new_n320), .b(new_n312), .c(new_n317), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n318), .b(new_n321), .o1(\s[28] ));
  norb02aa1n03x5               g227(.a(new_n309), .b(new_n317), .out0(new_n323));
  aoai13aa1n03x5               g228(.a(new_n323), .b(new_n315), .c(new_n201), .d(new_n304), .o1(new_n324));
  oao003aa1n02x5               g229(.a(\a[28] ), .b(\b[27] ), .c(new_n312), .carry(new_n325));
  xnrc02aa1n12x5               g230(.a(\b[28] ), .b(\a[29] ), .out0(new_n326));
  aoi012aa1n03x5               g231(.a(new_n326), .b(new_n324), .c(new_n325), .o1(new_n327));
  inv000aa1d42x5               g232(.a(new_n323), .o1(new_n328));
  tech160nm_fiaoi012aa1n03p5x5 g233(.a(new_n328), .b(new_n305), .c(new_n308), .o1(new_n329));
  nano22aa1n03x7               g234(.a(new_n329), .b(new_n325), .c(new_n326), .out0(new_n330));
  nor002aa1n02x5               g235(.a(new_n327), .b(new_n330), .o1(\s[29] ));
  xorb03aa1n02x5               g236(.a(new_n112), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1d15x5               g237(.a(new_n309), .b(new_n326), .c(new_n317), .out0(new_n333));
  aoai13aa1n02x7               g238(.a(new_n333), .b(new_n315), .c(new_n201), .d(new_n304), .o1(new_n334));
  oao003aa1n03x5               g239(.a(\a[29] ), .b(\b[28] ), .c(new_n325), .carry(new_n335));
  xnrc02aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .out0(new_n336));
  aoi012aa1n03x5               g241(.a(new_n336), .b(new_n334), .c(new_n335), .o1(new_n337));
  inv000aa1d42x5               g242(.a(new_n333), .o1(new_n338));
  tech160nm_fiaoi012aa1n03p5x5 g243(.a(new_n338), .b(new_n305), .c(new_n308), .o1(new_n339));
  nano22aa1n03x7               g244(.a(new_n339), .b(new_n335), .c(new_n336), .out0(new_n340));
  nor002aa1n02x5               g245(.a(new_n337), .b(new_n340), .o1(\s[30] ));
  nanb02aa1n02x5               g246(.a(\b[30] ), .b(\a[31] ), .out0(new_n342));
  nanb02aa1n02x5               g247(.a(\a[31] ), .b(\b[30] ), .out0(new_n343));
  norb02aa1n03x5               g248(.a(new_n333), .b(new_n336), .out0(new_n344));
  aoai13aa1n04x5               g249(.a(new_n344), .b(new_n315), .c(new_n201), .d(new_n304), .o1(new_n345));
  oao003aa1n02x5               g250(.a(\a[30] ), .b(\b[29] ), .c(new_n335), .carry(new_n346));
  aoi022aa1n03x5               g251(.a(new_n345), .b(new_n346), .c(new_n343), .d(new_n342), .o1(new_n347));
  nanp02aa1n02x5               g252(.a(new_n343), .b(new_n342), .o1(new_n348));
  inv000aa1n02x5               g253(.a(new_n346), .o1(new_n349));
  nona22aa1n02x4               g254(.a(new_n345), .b(new_n349), .c(new_n348), .out0(new_n350));
  norb02aa1n03x4               g255(.a(new_n350), .b(new_n347), .out0(\s[31] ));
  xnbna2aa1n03x5               g256(.a(new_n114), .b(new_n123), .c(new_n122), .out0(\s[3] ));
  aoai13aa1n02x5               g257(.a(new_n205), .b(new_n111), .c(new_n113), .d(new_n112), .o1(new_n353));
  aoi022aa1n02x5               g258(.a(new_n118), .b(new_n115), .c(new_n120), .d(new_n121), .o1(new_n354));
  aoi022aa1n02x5               g259(.a(new_n127), .b(new_n118), .c(new_n354), .d(new_n353), .o1(\s[4] ));
  xorb03aa1n02x5               g260(.a(new_n127), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n03x5               g261(.a(new_n105), .b(new_n129), .c(new_n206), .d(new_n126), .o1(new_n357));
  xorb03aa1n02x5               g262(.a(new_n357), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g263(.a(new_n130), .b(new_n131), .out0(new_n359));
  aoi012aa1n03x5               g264(.a(new_n106), .b(new_n357), .c(new_n359), .o1(new_n360));
  xnbna2aa1n03x5               g265(.a(new_n360), .b(new_n98), .c(new_n107), .out0(\s[7] ));
  aoai13aa1n02x5               g266(.a(new_n108), .b(new_n106), .c(new_n357), .d(new_n359), .o1(new_n362));
  xnbna2aa1n03x5               g267(.a(new_n102), .b(new_n362), .c(new_n98), .out0(\s[8] ));
  xnbna2aa1n03x5               g268(.a(new_n134), .b(new_n155), .c(new_n152), .out0(\s[9] ));
endmodule


