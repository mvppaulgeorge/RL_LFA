// Benchmark "adder" written by ABC on Wed Jul 17 19:49:45 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n337, new_n339,
    new_n340, new_n341, new_n342, new_n344, new_n346, new_n347, new_n348;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  tech160nm_fixorc02aa1n04x5   g002(.a(\a[3] ), .b(\b[2] ), .out0(new_n98));
  orn002aa1n03x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nand42aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n06x5               g005(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(new_n101));
  nand42aa1n02x5               g006(.a(new_n101), .b(new_n99), .o1(new_n102));
  nor042aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n08x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nona22aa1n03x5               g010(.a(new_n104), .b(new_n105), .c(new_n103), .out0(new_n106));
  tech160nm_fiaoi012aa1n04x5   g011(.a(new_n106), .b(new_n102), .c(new_n98), .o1(new_n107));
  nanp02aa1n09x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor042aa1n06x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1n06x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nano22aa1n06x5               g015(.a(new_n109), .b(new_n108), .c(new_n110), .out0(new_n111));
  xorc02aa1n12x5               g016(.a(\a[8] ), .b(\b[7] ), .out0(new_n112));
  nor002aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1n12x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand02aa1n06x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano23aa1n02x5               g020(.a(new_n114), .b(new_n113), .c(new_n115), .d(new_n104), .out0(new_n116));
  nand23aa1n03x5               g021(.a(new_n116), .b(new_n111), .c(new_n112), .o1(new_n117));
  orn002aa1n24x5               g022(.a(\a[6] ), .b(\b[5] ), .o(new_n118));
  oai112aa1n06x5               g023(.a(new_n118), .b(new_n108), .c(\b[4] ), .d(\a[5] ), .o1(new_n119));
  inv000aa1n02x5               g024(.a(new_n109), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  aoi013aa1n09x5               g026(.a(new_n121), .b(new_n111), .c(new_n119), .d(new_n112), .o1(new_n122));
  oai012aa1n18x5               g027(.a(new_n122), .b(new_n117), .c(new_n107), .o1(new_n123));
  nand42aa1n03x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  aoi012aa1n02x5               g029(.a(new_n97), .b(new_n123), .c(new_n124), .o1(new_n125));
  nor042aa1n06x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  inv000aa1n02x5               g031(.a(new_n126), .o1(new_n127));
  nand42aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  xnrc02aa1n02x5               g033(.a(\b[2] ), .b(\a[3] ), .out0(new_n129));
  norb03aa1n03x5               g034(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n129), .c(new_n101), .d(new_n99), .o1(new_n131));
  nanb03aa1n02x5               g036(.a(new_n109), .b(new_n110), .c(new_n108), .out0(new_n132));
  xnrc02aa1n02x5               g037(.a(\b[7] ), .b(\a[8] ), .out0(new_n133));
  nona23aa1n09x5               g038(.a(new_n104), .b(new_n115), .c(new_n114), .d(new_n113), .out0(new_n134));
  nona32aa1n03x5               g039(.a(new_n131), .b(new_n134), .c(new_n133), .d(new_n132), .out0(new_n135));
  nanb02aa1n12x5               g040(.a(new_n97), .b(new_n124), .out0(new_n136));
  norb03aa1d15x5               g041(.a(new_n128), .b(new_n97), .c(new_n126), .out0(new_n137));
  aoai13aa1n03x5               g042(.a(new_n137), .b(new_n136), .c(new_n135), .d(new_n122), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n125), .c(new_n128), .d(new_n127), .o1(\s[10] ));
  and002aa1n02x7               g044(.a(\b[10] ), .b(\a[11] ), .o(new_n140));
  nor002aa1d32x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norp02aa1n02x5               g046(.a(new_n140), .b(new_n141), .o1(new_n142));
  xobna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n128), .out0(\s[11] ));
  inv000aa1d42x5               g048(.a(new_n141), .o1(new_n144));
  nanp03aa1n03x5               g049(.a(new_n138), .b(new_n128), .c(new_n142), .o1(new_n145));
  nor002aa1n16x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand02aa1d20x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n03x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n145), .c(new_n144), .out0(\s[12] ));
  aoi112aa1n03x5               g054(.a(new_n140), .b(new_n141), .c(\a[10] ), .d(\b[9] ), .o1(new_n150));
  nona23aa1n03x5               g055(.a(new_n150), .b(new_n148), .c(new_n136), .d(new_n126), .out0(new_n151));
  aoi022aa1d18x5               g056(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n152));
  nona23aa1d18x5               g057(.a(new_n152), .b(new_n147), .c(new_n141), .d(new_n146), .out0(new_n153));
  oai012aa1d24x5               g058(.a(new_n147), .b(new_n146), .c(new_n141), .o1(new_n154));
  oai012aa1d24x5               g059(.a(new_n154), .b(new_n153), .c(new_n137), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n151), .c(new_n135), .d(new_n122), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n06x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n03x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g067(.a(new_n97), .o1(new_n163));
  nano32aa1n03x7               g068(.a(new_n153), .b(new_n127), .c(new_n124), .d(new_n163), .out0(new_n164));
  norp02aa1n04x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nanp02aa1n04x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nano23aa1n09x5               g071(.a(new_n159), .b(new_n165), .c(new_n166), .d(new_n160), .out0(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n155), .c(new_n123), .d(new_n164), .o1(new_n168));
  oai012aa1n06x5               g073(.a(new_n166), .b(new_n165), .c(new_n159), .o1(new_n169));
  nor022aa1n08x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand02aa1d04x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n168), .c(new_n169), .out0(\s[15] ));
  nanp02aa1n02x5               g078(.a(new_n168), .b(new_n169), .o1(new_n174));
  nor022aa1n06x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand02aa1n06x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  aoai13aa1n03x5               g082(.a(new_n177), .b(new_n170), .c(new_n174), .d(new_n172), .o1(new_n178));
  inv000aa1n06x5               g083(.a(new_n169), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n172), .b(new_n179), .c(new_n157), .d(new_n167), .o1(new_n180));
  nona22aa1n02x4               g085(.a(new_n180), .b(new_n177), .c(new_n170), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n178), .b(new_n181), .o1(\s[16] ));
  nanb02aa1n02x5               g087(.a(new_n159), .b(new_n160), .out0(new_n183));
  nanb02aa1n02x5               g088(.a(new_n165), .b(new_n166), .out0(new_n184));
  nona23aa1n09x5               g089(.a(new_n176), .b(new_n171), .c(new_n170), .d(new_n175), .out0(new_n185));
  nona32aa1n02x4               g090(.a(new_n164), .b(new_n185), .c(new_n184), .d(new_n183), .out0(new_n186));
  norp03aa1n02x5               g091(.a(new_n185), .b(new_n184), .c(new_n183), .o1(new_n187));
  tech160nm_fiao0012aa1n02p5x5 g092(.a(new_n175), .b(new_n170), .c(new_n176), .o(new_n188));
  oabi12aa1n03x5               g093(.a(new_n188), .b(new_n185), .c(new_n169), .out0(new_n189));
  aoi012aa1n06x5               g094(.a(new_n189), .b(new_n155), .c(new_n187), .o1(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n186), .c(new_n135), .d(new_n122), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[17] ), .o1(new_n193));
  nanb02aa1n02x5               g098(.a(\b[16] ), .b(new_n193), .out0(new_n194));
  nano23aa1n06x5               g099(.a(new_n170), .b(new_n175), .c(new_n176), .d(new_n171), .out0(new_n195));
  nand22aa1n03x5               g100(.a(new_n195), .b(new_n167), .o1(new_n196));
  nor042aa1n06x5               g101(.a(new_n151), .b(new_n196), .o1(new_n197));
  oai112aa1n02x5               g102(.a(new_n127), .b(new_n128), .c(\b[8] ), .d(\a[9] ), .o1(new_n198));
  nanp03aa1n03x5               g103(.a(new_n150), .b(new_n198), .c(new_n148), .o1(new_n199));
  tech160nm_fiaoi012aa1n04x5   g104(.a(new_n188), .b(new_n195), .c(new_n179), .o1(new_n200));
  aoai13aa1n09x5               g105(.a(new_n200), .b(new_n196), .c(new_n199), .d(new_n154), .o1(new_n201));
  xorc02aa1n12x5               g106(.a(\a[17] ), .b(\b[16] ), .out0(new_n202));
  aoai13aa1n03x5               g107(.a(new_n202), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n203));
  xnrc02aa1n02x5               g108(.a(\b[17] ), .b(\a[18] ), .out0(new_n204));
  xobna2aa1n03x5               g109(.a(new_n204), .b(new_n203), .c(new_n194), .out0(\s[18] ));
  inv000aa1d42x5               g110(.a(\a[18] ), .o1(new_n206));
  xroi22aa1d04x5               g111(.a(new_n193), .b(\b[16] ), .c(new_n206), .d(\b[17] ), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n208));
  oaih22aa1n04x5               g113(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n209));
  oaib12aa1n09x5               g114(.a(new_n209), .b(new_n206), .c(\b[17] ), .out0(new_n210));
  nor002aa1d24x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand42aa1d28x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nanb02aa1n18x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  xnbna2aa1n03x5               g119(.a(new_n214), .b(new_n208), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand22aa1n02x5               g121(.a(new_n208), .b(new_n210), .o1(new_n217));
  nor042aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand42aa1n16x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nanb02aa1n12x5               g124(.a(new_n218), .b(new_n219), .out0(new_n220));
  aoai13aa1n02x5               g125(.a(new_n220), .b(new_n211), .c(new_n217), .d(new_n214), .o1(new_n221));
  oaoi03aa1n02x5               g126(.a(\a[18] ), .b(\b[17] ), .c(new_n194), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n214), .b(new_n222), .c(new_n191), .d(new_n207), .o1(new_n223));
  nona22aa1n02x4               g128(.a(new_n223), .b(new_n220), .c(new_n211), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n221), .b(new_n224), .o1(\s[20] ));
  nano23aa1d12x5               g130(.a(new_n211), .b(new_n218), .c(new_n219), .d(new_n212), .out0(new_n226));
  nanb03aa1d24x5               g131(.a(new_n204), .b(new_n226), .c(new_n202), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n229));
  tech160nm_fioai012aa1n04x5   g134(.a(new_n219), .b(new_n218), .c(new_n211), .o1(new_n230));
  aobi12aa1n06x5               g135(.a(new_n230), .b(new_n226), .c(new_n222), .out0(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n229), .c(new_n231), .out0(\s[21] ));
  nanp02aa1n02x5               g139(.a(new_n229), .b(new_n231), .o1(new_n235));
  norp02aa1n04x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nor002aa1n02x5               g141(.a(\b[21] ), .b(\a[22] ), .o1(new_n237));
  nand42aa1n03x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nanb02aa1n06x5               g143(.a(new_n237), .b(new_n238), .out0(new_n239));
  aoai13aa1n02x5               g144(.a(new_n239), .b(new_n236), .c(new_n235), .d(new_n233), .o1(new_n240));
  oai013aa1d12x5               g145(.a(new_n230), .b(new_n210), .c(new_n213), .d(new_n220), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n233), .b(new_n241), .c(new_n191), .d(new_n228), .o1(new_n242));
  nona22aa1n03x5               g147(.a(new_n242), .b(new_n239), .c(new_n236), .out0(new_n243));
  nanp02aa1n02x5               g148(.a(new_n240), .b(new_n243), .o1(\s[22] ));
  nor042aa1n09x5               g149(.a(new_n232), .b(new_n239), .o1(new_n245));
  and003aa1n02x5               g150(.a(new_n207), .b(new_n245), .c(new_n226), .o(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n247));
  oaih12aa1n02x5               g152(.a(new_n238), .b(new_n237), .c(new_n236), .o1(new_n248));
  aobi12aa1n09x5               g153(.a(new_n248), .b(new_n241), .c(new_n245), .out0(new_n249));
  nor002aa1d32x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  nand02aa1n08x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  nanb02aa1d24x5               g156(.a(new_n250), .b(new_n251), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  xnbna2aa1n03x5               g158(.a(new_n253), .b(new_n247), .c(new_n249), .out0(\s[23] ));
  nand22aa1n03x5               g159(.a(new_n247), .b(new_n249), .o1(new_n255));
  nor002aa1d32x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nanp02aa1n04x5               g161(.a(\b[23] ), .b(\a[24] ), .o1(new_n257));
  nanb02aa1n02x5               g162(.a(new_n256), .b(new_n257), .out0(new_n258));
  aoai13aa1n02x5               g163(.a(new_n258), .b(new_n250), .c(new_n255), .d(new_n253), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n249), .o1(new_n260));
  aoai13aa1n04x5               g165(.a(new_n253), .b(new_n260), .c(new_n191), .d(new_n246), .o1(new_n261));
  nona22aa1n02x4               g166(.a(new_n261), .b(new_n258), .c(new_n250), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n259), .b(new_n262), .o1(\s[24] ));
  nona23aa1d18x5               g168(.a(new_n257), .b(new_n251), .c(new_n250), .d(new_n256), .out0(new_n264));
  inv040aa1n03x5               g169(.a(new_n264), .o1(new_n265));
  nano22aa1n03x7               g170(.a(new_n227), .b(new_n245), .c(new_n265), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n256), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(new_n250), .b(new_n257), .o1(new_n269));
  oai112aa1n04x5               g174(.a(new_n269), .b(new_n268), .c(new_n264), .d(new_n248), .o1(new_n270));
  aoi013aa1n09x5               g175(.a(new_n270), .b(new_n241), .c(new_n245), .d(new_n265), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n267), .c(new_n271), .out0(\s[25] ));
  nand22aa1n02x5               g178(.a(new_n267), .b(new_n271), .o1(new_n274));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  tech160nm_fixnrc02aa1n04x5   g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  aoai13aa1n02x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .d(new_n272), .o1(new_n277));
  inv000aa1n02x5               g182(.a(new_n271), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n272), .b(new_n278), .c(new_n191), .d(new_n266), .o1(new_n279));
  nona22aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n275), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n277), .b(new_n280), .o1(\s[26] ));
  norb02aa1n12x5               g186(.a(new_n272), .b(new_n276), .out0(new_n282));
  nano32aa1d15x5               g187(.a(new_n227), .b(new_n282), .c(new_n245), .d(new_n265), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n201), .c(new_n123), .d(new_n197), .o1(new_n284));
  nano22aa1n02x5               g189(.a(new_n231), .b(new_n245), .c(new_n265), .out0(new_n285));
  inv000aa1d42x5               g190(.a(\a[26] ), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\b[25] ), .o1(new_n287));
  oaoi03aa1n02x5               g192(.a(new_n286), .b(new_n287), .c(new_n275), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  oaoi13aa1n06x5               g194(.a(new_n289), .b(new_n282), .c(new_n285), .d(new_n270), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnbna2aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n284), .out0(\s[27] ));
  nanp02aa1n03x5               g197(.a(new_n290), .b(new_n284), .o1(new_n293));
  norp02aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  norp02aa1n02x5               g199(.a(\b[27] ), .b(\a[28] ), .o1(new_n295));
  nanp02aa1n02x5               g200(.a(\b[27] ), .b(\a[28] ), .o1(new_n296));
  norb02aa1n09x5               g201(.a(new_n296), .b(new_n295), .out0(new_n297));
  inv000aa1d42x5               g202(.a(new_n297), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n294), .c(new_n293), .d(new_n291), .o1(new_n299));
  norp03aa1n03x5               g204(.a(new_n248), .b(new_n252), .c(new_n258), .o1(new_n300));
  nano22aa1n03x7               g205(.a(new_n300), .b(new_n268), .c(new_n269), .out0(new_n301));
  nona32aa1n09x5               g206(.a(new_n241), .b(new_n264), .c(new_n239), .d(new_n232), .out0(new_n302));
  inv000aa1d42x5               g207(.a(new_n282), .o1(new_n303));
  aoai13aa1n12x5               g208(.a(new_n288), .b(new_n303), .c(new_n302), .d(new_n301), .o1(new_n304));
  aoai13aa1n02x7               g209(.a(new_n291), .b(new_n304), .c(new_n191), .d(new_n283), .o1(new_n305));
  nona22aa1n03x5               g210(.a(new_n305), .b(new_n298), .c(new_n294), .out0(new_n306));
  nanp02aa1n03x5               g211(.a(new_n299), .b(new_n306), .o1(\s[28] ));
  norb02aa1n02x5               g212(.a(new_n291), .b(new_n298), .out0(new_n308));
  aoai13aa1n06x5               g213(.a(new_n308), .b(new_n304), .c(new_n191), .d(new_n283), .o1(new_n309));
  oai012aa1n02x5               g214(.a(new_n296), .b(new_n295), .c(new_n294), .o1(new_n310));
  nanp02aa1n03x5               g215(.a(new_n309), .b(new_n310), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n02x7               g218(.a(new_n311), .b(new_n312), .c(new_n309), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g220(.a(new_n291), .b(new_n312), .c(new_n297), .o(new_n316));
  aoai13aa1n06x5               g221(.a(new_n316), .b(new_n304), .c(new_n191), .d(new_n283), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .carry(new_n318));
  nanp02aa1n03x5               g223(.a(new_n317), .b(new_n318), .o1(new_n319));
  xorc02aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .out0(new_n320));
  norp02aa1n02x5               g225(.a(\b[28] ), .b(\a[29] ), .o1(new_n321));
  aoi012aa1n02x5               g226(.a(new_n310), .b(\a[29] ), .c(\b[28] ), .o1(new_n322));
  norp03aa1n02x5               g227(.a(new_n322), .b(new_n320), .c(new_n321), .o1(new_n323));
  aoi022aa1n02x7               g228(.a(new_n319), .b(new_n320), .c(new_n317), .d(new_n323), .o1(\s[30] ));
  and003aa1n02x5               g229(.a(new_n308), .b(new_n320), .c(new_n312), .o(new_n325));
  aoai13aa1n04x5               g230(.a(new_n325), .b(new_n304), .c(new_n191), .d(new_n283), .o1(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n318), .carry(new_n327));
  nanb02aa1n02x5               g232(.a(\b[30] ), .b(\a[31] ), .out0(new_n328));
  nanb02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n326), .b(new_n327), .c(new_n329), .d(new_n328), .o1(new_n330));
  aobi12aa1n03x5               g235(.a(new_n325), .b(new_n290), .c(new_n284), .out0(new_n331));
  xnrc02aa1n02x5               g236(.a(\b[30] ), .b(\a[31] ), .out0(new_n332));
  nano22aa1n03x7               g237(.a(new_n331), .b(new_n327), .c(new_n332), .out0(new_n333));
  nor002aa1n02x5               g238(.a(new_n330), .b(new_n333), .o1(\s[31] ));
  xnbna2aa1n03x5               g239(.a(new_n98), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  norb02aa1n02x5               g240(.a(new_n104), .b(new_n105), .out0(new_n336));
  aoi012aa1n02x5               g241(.a(new_n103), .b(new_n102), .c(new_n98), .o1(new_n337));
  oai012aa1n02x5               g242(.a(new_n131), .b(new_n337), .c(new_n336), .o1(\s[4] ));
  nano22aa1n02x4               g243(.a(new_n114), .b(new_n104), .c(new_n115), .out0(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n106), .c(new_n102), .d(new_n98), .o1(new_n340));
  inv000aa1d42x5               g245(.a(new_n114), .o1(new_n341));
  aoi022aa1n02x5               g246(.a(new_n131), .b(new_n104), .c(new_n115), .d(new_n341), .o1(new_n342));
  norb02aa1n02x5               g247(.a(new_n340), .b(new_n342), .out0(\s[5] ));
  ao0022aa1n03x5               g248(.a(new_n340), .b(new_n341), .c(new_n118), .d(new_n108), .o(new_n344));
  oaib12aa1n02x5               g249(.a(new_n344), .b(new_n119), .c(new_n340), .out0(\s[6] ));
  norb02aa1n02x5               g250(.a(new_n110), .b(new_n109), .out0(new_n346));
  aoai13aa1n02x5               g251(.a(new_n111), .b(new_n119), .c(new_n131), .d(new_n339), .o1(new_n347));
  aboi22aa1n03x5               g252(.a(new_n119), .b(new_n340), .c(\a[6] ), .d(\b[5] ), .out0(new_n348));
  oa0012aa1n02x5               g253(.a(new_n347), .b(new_n348), .c(new_n346), .o(\s[7] ));
  xnbna2aa1n03x5               g254(.a(new_n112), .b(new_n347), .c(new_n120), .out0(\s[8] ));
  xorb03aa1n02x5               g255(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


