// Benchmark "adder" written by ABC on Wed Jul 17 21:04:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n318,
    new_n319, new_n320, new_n322, new_n323, new_n325, new_n326, new_n327,
    new_n328, new_n330, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  tech160nm_fixnrc02aa1n02p5x5 g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor042aa1n03x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  tech160nm_fioai012aa1n03p5x5 g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  tech160nm_fixnrc02aa1n05x5   g009(.a(\b[3] ), .b(\a[4] ), .out0(new_n105));
  nor042aa1n02x5               g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n103), .c(new_n99), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nor022aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand42aa1n20x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  norb02aa1n03x5               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  aoi022aa1d24x5               g016(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[5] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\b[4] ), .o1(new_n114));
  aoi022aa1d24x5               g019(.a(new_n114), .b(new_n113), .c(\a[4] ), .d(\b[3] ), .o1(new_n115));
  nor002aa1d24x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor022aa1n04x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nona22aa1n02x4               g022(.a(new_n115), .b(new_n116), .c(new_n117), .out0(new_n118));
  nano32aa1n03x7               g023(.a(new_n118), .b(new_n111), .c(new_n112), .d(new_n108), .out0(new_n119));
  oai012aa1n02x5               g024(.a(new_n110), .b(new_n116), .c(new_n109), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n112), .b(new_n110), .c(new_n116), .d(new_n109), .out0(new_n121));
  and002aa1n03x5               g026(.a(\b[5] ), .b(\a[6] ), .o(new_n122));
  aoi112aa1n06x5               g027(.a(new_n122), .b(new_n117), .c(new_n113), .d(new_n114), .o1(new_n123));
  oai012aa1n06x5               g028(.a(new_n120), .b(new_n121), .c(new_n123), .o1(new_n124));
  nand42aa1n08x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n97), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n124), .c(new_n107), .d(new_n119), .o1(new_n127));
  nor042aa1n03x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n129), .o1(new_n131));
  oai022aa1d24x5               g036(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n132));
  nona22aa1n02x4               g037(.a(new_n127), .b(new_n131), .c(new_n132), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n130), .c(new_n98), .d(new_n127), .o1(\s[10] ));
  nano23aa1d15x5               g039(.a(new_n97), .b(new_n128), .c(new_n129), .d(new_n125), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n124), .c(new_n107), .d(new_n119), .o1(new_n136));
  oaib12aa1n02x5               g041(.a(new_n136), .b(new_n131), .c(new_n132), .out0(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n02x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1n10x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nor042aa1n02x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanp02aa1n12x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n139), .c(new_n137), .d(new_n140), .o1(new_n144));
  oai022aa1n06x5               g049(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n140), .b(new_n139), .out0(new_n146));
  aob012aa1n02x5               g051(.a(new_n142), .b(new_n137), .c(new_n146), .out0(new_n147));
  oai012aa1n02x5               g052(.a(new_n144), .b(new_n147), .c(new_n145), .o1(\s[12] ));
  nano23aa1n06x5               g053(.a(new_n139), .b(new_n141), .c(new_n142), .d(new_n140), .out0(new_n149));
  nand22aa1n09x5               g054(.a(new_n149), .b(new_n135), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n124), .c(new_n107), .d(new_n119), .o1(new_n152));
  aoi022aa1n06x5               g057(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  aoai13aa1n04x5               g058(.a(new_n142), .b(new_n145), .c(new_n132), .d(new_n153), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(new_n152), .b(new_n154), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d24x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nand02aa1n03x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanp03aa1n02x5               g064(.a(new_n155), .b(new_n158), .c(new_n159), .o1(new_n160));
  nor002aa1n06x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  nona23aa1n02x4               g068(.a(new_n160), .b(new_n162), .c(new_n161), .d(new_n157), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n163), .c(new_n158), .d(new_n160), .o1(\s[14] ));
  nona23aa1n03x5               g070(.a(new_n162), .b(new_n159), .c(new_n157), .d(new_n161), .out0(new_n166));
  oaih12aa1n02x5               g071(.a(new_n162), .b(new_n161), .c(new_n157), .o1(new_n167));
  oai012aa1n03x5               g072(.a(new_n167), .b(new_n154), .c(new_n166), .o1(new_n168));
  oabi12aa1n02x5               g073(.a(new_n168), .b(new_n152), .c(new_n166), .out0(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand42aa1n03x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  nor042aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand42aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n171), .c(new_n169), .d(new_n172), .o1(new_n177));
  nona22aa1n02x4               g082(.a(new_n175), .b(new_n174), .c(new_n171), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n177), .b(new_n178), .c(new_n173), .d(new_n169), .o1(\s[16] ));
  nano23aa1n02x4               g084(.a(new_n157), .b(new_n161), .c(new_n162), .d(new_n159), .out0(new_n180));
  nano23aa1n03x7               g085(.a(new_n171), .b(new_n174), .c(new_n175), .d(new_n172), .out0(new_n181));
  nano22aa1n03x7               g086(.a(new_n150), .b(new_n180), .c(new_n181), .out0(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n124), .c(new_n107), .d(new_n119), .o1(new_n183));
  oai022aa1n02x5               g088(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n184));
  aoi022aa1n06x5               g089(.a(new_n168), .b(new_n181), .c(new_n175), .d(new_n184), .o1(new_n185));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n183), .out0(\s[17] ));
  nor042aa1n04x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n188), .o1(new_n189));
  nanp02aa1n12x5               g094(.a(new_n185), .b(new_n183), .o1(new_n190));
  nanp02aa1n06x5               g095(.a(new_n190), .b(new_n186), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[18] ), .b(\b[17] ), .out0(new_n192));
  nand42aa1n02x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  oai022aa1d18x5               g098(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n194));
  nanb03aa1n02x5               g099(.a(new_n194), .b(new_n191), .c(new_n193), .out0(new_n195));
  aoai13aa1n02x5               g100(.a(new_n195), .b(new_n192), .c(new_n189), .d(new_n191), .o1(\s[18] ));
  nanp02aa1n02x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  norp02aa1n02x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nano23aa1n06x5               g103(.a(new_n188), .b(new_n198), .c(new_n193), .d(new_n197), .out0(new_n199));
  oaoi03aa1n02x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n200));
  xorc02aa1n02x5               g105(.a(\a[19] ), .b(\b[18] ), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n202));
  aoi112aa1n02x5               g107(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n202), .b(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[18] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  xorc02aa1n02x5               g113(.a(\a[20] ), .b(\b[19] ), .out0(new_n209));
  nand02aa1d08x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  oai022aa1n03x5               g116(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n212));
  nona22aa1n02x5               g117(.a(new_n202), .b(new_n211), .c(new_n212), .out0(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n208), .d(new_n202), .o1(\s[20] ));
  nanp03aa1n02x5               g119(.a(new_n199), .b(new_n201), .c(new_n209), .o1(new_n215));
  oai112aa1n03x5               g120(.a(new_n194), .b(new_n193), .c(new_n207), .d(new_n206), .o1(new_n216));
  aoib12aa1n02x5               g121(.a(new_n211), .b(new_n216), .c(new_n212), .out0(new_n217));
  inv000aa1n02x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n215), .c(new_n185), .d(new_n183), .o1(new_n219));
  xorb03aa1n02x5               g124(.a(new_n219), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  xnrc02aa1n02x5               g128(.a(\b[21] ), .b(\a[22] ), .out0(new_n224));
  aoai13aa1n02x5               g129(.a(new_n224), .b(new_n221), .c(new_n219), .d(new_n223), .o1(new_n225));
  inv000aa1d42x5               g130(.a(\a[22] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[21] ), .o1(new_n227));
  nand42aa1n03x5               g132(.a(new_n219), .b(new_n223), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n221), .b(new_n226), .c(new_n227), .o1(new_n229));
  oai112aa1n03x5               g134(.a(new_n228), .b(new_n229), .c(new_n227), .d(new_n226), .o1(new_n230));
  nanp02aa1n03x5               g135(.a(new_n230), .b(new_n225), .o1(\s[22] ));
  inv030aa1n04x5               g136(.a(new_n221), .o1(new_n232));
  nano22aa1n02x4               g137(.a(new_n224), .b(new_n232), .c(new_n222), .out0(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n215), .out0(new_n234));
  nanb02aa1n02x5               g139(.a(new_n212), .b(new_n216), .out0(new_n235));
  nano32aa1n03x7               g140(.a(new_n224), .b(new_n232), .c(new_n222), .d(new_n210), .out0(new_n236));
  oaoi03aa1n12x5               g141(.a(\a[22] ), .b(\b[21] ), .c(new_n232), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aob012aa1n02x5               g143(.a(new_n238), .b(new_n235), .c(new_n236), .out0(new_n239));
  xorc02aa1n02x5               g144(.a(\a[23] ), .b(\b[22] ), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n239), .c(new_n190), .d(new_n234), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(new_n240), .b(new_n237), .c(new_n235), .d(new_n236), .o1(new_n242));
  aobi12aa1n02x5               g147(.a(new_n242), .b(new_n190), .c(new_n234), .out0(new_n243));
  norb02aa1n02x5               g148(.a(new_n241), .b(new_n243), .out0(\s[23] ));
  norp02aa1n02x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xorc02aa1n02x5               g151(.a(\a[24] ), .b(\b[23] ), .out0(new_n247));
  and002aa1n02x5               g152(.a(\b[23] ), .b(\a[24] ), .o(new_n248));
  oai022aa1n02x5               g153(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n249));
  nona22aa1n02x5               g154(.a(new_n241), .b(new_n248), .c(new_n249), .out0(new_n250));
  aoai13aa1n03x5               g155(.a(new_n250), .b(new_n247), .c(new_n246), .d(new_n241), .o1(\s[24] ));
  inv000aa1d42x5               g156(.a(\a[23] ), .o1(new_n252));
  inv000aa1d42x5               g157(.a(\a[24] ), .o1(new_n253));
  xroi22aa1d04x5               g158(.a(new_n252), .b(\b[22] ), .c(new_n253), .d(\b[23] ), .out0(new_n254));
  nano22aa1n02x4               g159(.a(new_n215), .b(new_n254), .c(new_n233), .out0(new_n255));
  aoai13aa1n03x5               g160(.a(new_n254), .b(new_n237), .c(new_n235), .d(new_n236), .o1(new_n256));
  oaib12aa1n02x5               g161(.a(new_n249), .b(new_n253), .c(\b[23] ), .out0(new_n257));
  nanp02aa1n02x5               g162(.a(new_n256), .b(new_n257), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[24] ), .b(\a[25] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n258), .c(new_n190), .d(new_n255), .o1(new_n261));
  aoi112aa1n02x5               g166(.a(new_n260), .b(new_n258), .c(new_n190), .d(new_n255), .o1(new_n262));
  norb02aa1n02x5               g167(.a(new_n261), .b(new_n262), .out0(\s[25] ));
  norp02aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n02x5               g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  and002aa1n02x5               g171(.a(\b[25] ), .b(\a[26] ), .o(new_n267));
  oai022aa1n02x5               g172(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n268));
  nona22aa1n03x5               g173(.a(new_n261), .b(new_n267), .c(new_n268), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n266), .c(new_n265), .d(new_n261), .o1(\s[26] ));
  norb02aa1n09x5               g175(.a(new_n266), .b(new_n259), .out0(new_n271));
  nano32aa1n03x7               g176(.a(new_n215), .b(new_n271), .c(new_n233), .d(new_n254), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n271), .o1(new_n273));
  aob012aa1n02x5               g178(.a(new_n268), .b(\b[25] ), .c(\a[26] ), .out0(new_n274));
  aoai13aa1n09x5               g179(.a(new_n274), .b(new_n273), .c(new_n256), .d(new_n257), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[27] ), .b(\b[26] ), .out0(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n275), .c(new_n190), .d(new_n272), .o1(new_n277));
  aoi112aa1n02x5               g182(.a(new_n276), .b(new_n275), .c(new_n190), .d(new_n272), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n277), .b(new_n278), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  xorc02aa1n02x5               g186(.a(\a[28] ), .b(\b[27] ), .out0(new_n282));
  and002aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .o(new_n283));
  oai022aa1d24x5               g188(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n284));
  nona22aa1n06x5               g189(.a(new_n277), .b(new_n283), .c(new_n284), .out0(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n282), .c(new_n281), .d(new_n277), .o1(\s[28] ));
  xorc02aa1n02x5               g191(.a(\a[29] ), .b(\b[28] ), .out0(new_n287));
  and002aa1n02x5               g192(.a(new_n282), .b(new_n276), .o(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n275), .c(new_n190), .d(new_n272), .o1(new_n289));
  inv000aa1d42x5               g194(.a(\b[27] ), .o1(new_n290));
  oaib12aa1n06x5               g195(.a(new_n284), .b(new_n290), .c(\a[28] ), .out0(new_n291));
  nanp03aa1n03x5               g196(.a(new_n289), .b(new_n291), .c(new_n287), .o1(new_n292));
  inv020aa1n03x5               g197(.a(new_n272), .o1(new_n293));
  tech160nm_fiaoi012aa1n04x5   g198(.a(new_n293), .b(new_n185), .c(new_n183), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n291), .o1(new_n295));
  oaoi13aa1n02x7               g200(.a(new_n295), .b(new_n288), .c(new_n294), .d(new_n275), .o1(new_n296));
  oai012aa1n03x5               g201(.a(new_n292), .b(new_n296), .c(new_n287), .o1(\s[29] ));
  xorb03aa1n02x5               g202(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g203(.a(new_n276), .b(new_n287), .c(new_n282), .o(new_n299));
  tech160nm_fioaoi03aa1n03p5x5 g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .o1(new_n300));
  oaoi13aa1n02x7               g205(.a(new_n300), .b(new_n299), .c(new_n294), .d(new_n275), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[30] ), .b(\b[29] ), .out0(new_n302));
  aoai13aa1n02x5               g207(.a(new_n299), .b(new_n275), .c(new_n190), .d(new_n272), .o1(new_n303));
  norb02aa1n03x5               g208(.a(new_n302), .b(new_n300), .out0(new_n304));
  nand02aa1n02x5               g209(.a(new_n303), .b(new_n304), .o1(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(new_n301), .c(new_n302), .o1(\s[30] ));
  and003aa1n02x5               g211(.a(new_n288), .b(new_n302), .c(new_n287), .o(new_n307));
  aoi012aa1n02x5               g212(.a(new_n304), .b(\a[30] ), .c(\b[29] ), .o1(new_n308));
  oaoi13aa1n02x7               g213(.a(new_n308), .b(new_n307), .c(new_n294), .d(new_n275), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[31] ), .b(\b[30] ), .out0(new_n310));
  aoai13aa1n02x5               g215(.a(new_n307), .b(new_n275), .c(new_n190), .d(new_n272), .o1(new_n311));
  norb02aa1n02x5               g216(.a(new_n310), .b(new_n308), .out0(new_n312));
  nand02aa1n02x5               g217(.a(new_n311), .b(new_n312), .o1(new_n313));
  tech160nm_fioai012aa1n02p5x5 g218(.a(new_n313), .b(new_n309), .c(new_n310), .o1(\s[31] ));
  xnrb03aa1n02x5               g219(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g220(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n316));
  aob012aa1n02x5               g221(.a(new_n107), .b(new_n316), .c(new_n105), .out0(\s[4] ));
  nanp02aa1n02x5               g222(.a(\b[3] ), .b(\a[4] ), .o1(new_n318));
  nanp02aa1n02x5               g223(.a(new_n114), .b(new_n113), .o1(new_n319));
  aoi022aa1n02x5               g224(.a(new_n107), .b(new_n318), .c(new_n319), .d(new_n108), .o1(new_n320));
  aoi013aa1n02x4               g225(.a(new_n320), .b(new_n115), .c(new_n108), .d(new_n107), .o1(\s[5] ));
  norp02aa1n02x5               g226(.a(new_n122), .b(new_n117), .o1(new_n322));
  nanp03aa1n02x5               g227(.a(new_n107), .b(new_n108), .c(new_n115), .o1(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n322), .b(new_n323), .c(new_n319), .out0(\s[6] ));
  norb02aa1n02x5               g229(.a(new_n112), .b(new_n116), .out0(new_n325));
  aob012aa1n02x5               g230(.a(new_n325), .b(new_n323), .c(new_n123), .out0(new_n326));
  xnrc02aa1n02x5               g231(.a(\b[6] ), .b(\a[7] ), .out0(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n122), .c(new_n323), .d(new_n123), .o1(new_n328));
  and002aa1n02x5               g233(.a(new_n328), .b(new_n326), .o(\s[7] ));
  inv000aa1d42x5               g234(.a(new_n116), .o1(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n111), .b(new_n326), .c(new_n330), .out0(\s[8] ));
  aoi112aa1n02x5               g236(.a(new_n126), .b(new_n124), .c(new_n107), .d(new_n119), .o1(new_n332));
  norb02aa1n02x5               g237(.a(new_n127), .b(new_n332), .out0(\s[9] ));
endmodule


