// Benchmark "adder" written by ABC on Thu Jul 18 07:34:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n327, new_n329, new_n332, new_n334,
    new_n336, new_n337, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n06x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  tech160nm_fiaoi012aa1n05x5   g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1d32x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n02x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  tech160nm_fioai012aa1n03p5x5 g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oaih12aa1n06x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  norp02aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1d04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n02x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  nor002aa1n12x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  tech160nm_finor002aa1n03p5x5 g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nona23aa1n02x5               g023(.a(new_n117), .b(new_n116), .c(new_n118), .d(new_n115), .out0(new_n119));
  nor042aa1n03x5               g024(.a(new_n119), .b(new_n114), .o1(new_n120));
  oai012aa1n02x7               g025(.a(new_n117), .b(new_n118), .c(new_n115), .o1(new_n121));
  oai012aa1n02x5               g026(.a(new_n111), .b(new_n112), .c(new_n110), .o1(new_n122));
  oai012aa1n04x7               g027(.a(new_n122), .b(new_n114), .c(new_n121), .o1(new_n123));
  tech160nm_fixorc02aa1n03p5x5 g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(new_n109), .d(new_n120), .o1(new_n125));
  tech160nm_fixorc02aa1n03p5x5 g030(.a(\a[10] ), .b(\b[9] ), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n126), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(new_n99), .o1(new_n128));
  aob012aa1n02x5               g033(.a(new_n128), .b(new_n100), .c(new_n101), .out0(new_n129));
  norb02aa1n02x7               g034(.a(new_n104), .b(new_n103), .out0(new_n130));
  norb02aa1n02x5               g035(.a(new_n106), .b(new_n105), .out0(new_n131));
  nanp03aa1n02x5               g036(.a(new_n129), .b(new_n130), .c(new_n131), .o1(new_n132));
  nano23aa1n02x4               g037(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n133));
  nanb02aa1n02x5               g038(.a(new_n115), .b(new_n116), .out0(new_n134));
  nanb02aa1n02x5               g039(.a(new_n118), .b(new_n117), .out0(new_n135));
  nona22aa1n02x4               g040(.a(new_n133), .b(new_n134), .c(new_n135), .out0(new_n136));
  inv000aa1d42x5               g041(.a(new_n115), .o1(new_n137));
  oaoi03aa1n02x5               g042(.a(\a[6] ), .b(\b[5] ), .c(new_n137), .o1(new_n138));
  aobi12aa1n02x5               g043(.a(new_n122), .b(new_n133), .c(new_n138), .out0(new_n139));
  aoai13aa1n06x5               g044(.a(new_n139), .b(new_n136), .c(new_n132), .d(new_n108), .o1(new_n140));
  and002aa1n02x5               g045(.a(new_n126), .b(new_n124), .o(new_n141));
  norp02aa1n04x5               g046(.a(\b[9] ), .b(\a[10] ), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(\b[9] ), .b(\a[10] ), .o1(new_n143));
  oai012aa1n12x5               g048(.a(new_n143), .b(new_n142), .c(new_n97), .o1(new_n144));
  aob012aa1n02x5               g049(.a(new_n144), .b(new_n140), .c(new_n141), .out0(new_n145));
  xorb03aa1n02x5               g050(.a(new_n145), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nanp02aa1n04x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  nor022aa1n06x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n147), .b(new_n148), .out0(new_n149));
  nor022aa1n08x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand42aa1n04x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nanb02aa1n02x5               g056(.a(new_n150), .b(new_n151), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n148), .c(new_n145), .d(new_n149), .o1(new_n153));
  nona22aa1n02x4               g058(.a(new_n151), .b(new_n150), .c(new_n148), .out0(new_n154));
  aoai13aa1n02x5               g059(.a(new_n153), .b(new_n154), .c(new_n149), .d(new_n145), .o1(\s[12] ));
  nona23aa1n02x4               g060(.a(new_n147), .b(new_n151), .c(new_n150), .d(new_n148), .out0(new_n156));
  nano22aa1n02x4               g061(.a(new_n156), .b(new_n124), .c(new_n126), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n123), .c(new_n109), .d(new_n120), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n144), .o1(new_n159));
  nano23aa1n03x7               g064(.a(new_n150), .b(new_n148), .c(new_n151), .d(new_n147), .out0(new_n160));
  oai012aa1n02x5               g065(.a(new_n151), .b(new_n150), .c(new_n148), .o1(new_n161));
  aobi12aa1n02x7               g066(.a(new_n161), .b(new_n160), .c(new_n159), .out0(new_n162));
  nand42aa1d28x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nor042aa1n04x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  xnbna2aa1n03x5               g070(.a(new_n165), .b(new_n158), .c(new_n162), .out0(\s[13] ));
  orn002aa1n24x5               g071(.a(\a[13] ), .b(\b[12] ), .o(new_n167));
  tech160nm_fioai012aa1n05x5   g072(.a(new_n161), .b(new_n156), .c(new_n144), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n165), .b(new_n168), .c(new_n140), .d(new_n157), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand42aa1n20x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n169), .c(new_n167), .out0(\s[14] ));
  oaoi03aa1n12x5               g078(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  nano23aa1d15x5               g080(.a(new_n170), .b(new_n164), .c(new_n171), .d(new_n163), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n175), .b(new_n177), .c(new_n158), .d(new_n162), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand42aa1n06x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  nor022aa1n08x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  nor022aa1n04x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nand42aa1n10x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n183), .b(new_n184), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n181), .c(new_n178), .d(new_n182), .o1(new_n186));
  nona22aa1n02x4               g091(.a(new_n184), .b(new_n183), .c(new_n181), .out0(new_n187));
  aoai13aa1n02x5               g092(.a(new_n186), .b(new_n187), .c(new_n178), .d(new_n182), .o1(\s[16] ));
  nano23aa1n06x5               g093(.a(new_n183), .b(new_n181), .c(new_n184), .d(new_n180), .out0(new_n189));
  nand02aa1d04x5               g094(.a(new_n189), .b(new_n176), .o1(new_n190));
  nano32aa1n09x5               g095(.a(new_n190), .b(new_n160), .c(new_n126), .d(new_n124), .out0(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n123), .c(new_n109), .d(new_n120), .o1(new_n192));
  aoi022aa1n09x5               g097(.a(new_n189), .b(new_n174), .c(new_n184), .d(new_n187), .o1(new_n193));
  inv030aa1n03x5               g098(.a(new_n193), .o1(new_n194));
  aoib12aa1n12x5               g099(.a(new_n194), .b(new_n168), .c(new_n190), .out0(new_n195));
  tech160nm_fixorc02aa1n03p5x5 g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n192), .c(new_n195), .out0(\s[17] ));
  nor042aa1n06x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  oai012aa1n02x7               g104(.a(new_n193), .b(new_n162), .c(new_n190), .o1(new_n200));
  aoai13aa1n02x5               g105(.a(new_n196), .b(new_n200), .c(new_n140), .d(new_n191), .o1(new_n201));
  xnrc02aa1n02x5               g106(.a(\b[17] ), .b(\a[18] ), .out0(new_n202));
  xobna2aa1n03x5               g107(.a(new_n202), .b(new_n201), .c(new_n199), .out0(\s[18] ));
  inv000aa1d42x5               g108(.a(\a[17] ), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\a[18] ), .o1(new_n205));
  xroi22aa1d04x5               g110(.a(new_n204), .b(\b[16] ), .c(new_n205), .d(\b[17] ), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  inv000aa1d42x5               g112(.a(\b[17] ), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(new_n205), .b(new_n208), .c(new_n198), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n207), .c(new_n192), .d(new_n195), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n04x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nor002aa1n04x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  norb02aa1n03x5               g120(.a(new_n210), .b(new_n215), .out0(new_n216));
  nor042aa1n02x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1n06x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n214), .c(new_n210), .d(new_n213), .o1(new_n220));
  nona22aa1n03x5               g125(.a(new_n218), .b(new_n217), .c(new_n214), .out0(new_n221));
  oai012aa1n03x5               g126(.a(new_n220), .b(new_n216), .c(new_n221), .o1(\s[20] ));
  nano23aa1n06x5               g127(.a(new_n217), .b(new_n214), .c(new_n218), .d(new_n213), .out0(new_n223));
  nanb03aa1n09x5               g128(.a(new_n202), .b(new_n223), .c(new_n196), .out0(new_n224));
  tech160nm_fioaoi03aa1n03p5x5 g129(.a(\a[18] ), .b(\b[17] ), .c(new_n199), .o1(new_n225));
  aoi022aa1n03x5               g130(.a(new_n223), .b(new_n225), .c(new_n218), .d(new_n221), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n224), .c(new_n192), .d(new_n195), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  xnrc02aa1n12x5               g133(.a(\b[20] ), .b(\a[21] ), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  norp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  tech160nm_fixnrc02aa1n05x5   g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n231), .c(new_n227), .d(new_n230), .o1(new_n233));
  oabi12aa1n02x5               g138(.a(new_n232), .b(\a[21] ), .c(\b[20] ), .out0(new_n234));
  aoai13aa1n03x5               g139(.a(new_n233), .b(new_n234), .c(new_n230), .d(new_n227), .o1(\s[22] ));
  nor042aa1n04x5               g140(.a(new_n232), .b(new_n229), .o1(new_n236));
  nanp03aa1n02x5               g141(.a(new_n206), .b(new_n236), .c(new_n223), .o1(new_n237));
  nona23aa1n09x5               g142(.a(new_n213), .b(new_n218), .c(new_n217), .d(new_n214), .out0(new_n238));
  oai012aa1n02x5               g143(.a(new_n218), .b(new_n217), .c(new_n214), .o1(new_n239));
  oai012aa1n04x7               g144(.a(new_n239), .b(new_n238), .c(new_n209), .o1(new_n240));
  orn002aa1n02x5               g145(.a(\a[21] ), .b(\b[20] ), .o(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n241), .o1(new_n242));
  aoi012aa1n02x5               g147(.a(new_n242), .b(new_n240), .c(new_n236), .o1(new_n243));
  aoai13aa1n04x5               g148(.a(new_n243), .b(new_n237), .c(new_n192), .d(new_n195), .o1(new_n244));
  xorb03aa1n02x5               g149(.a(new_n244), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[22] ), .b(\a[23] ), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  xnrc02aa1n12x5               g153(.a(\b[23] ), .b(\a[24] ), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n246), .c(new_n244), .d(new_n248), .o1(new_n250));
  norp02aa1n02x5               g155(.a(new_n249), .b(new_n246), .o1(new_n251));
  aob012aa1n03x5               g156(.a(new_n251), .b(new_n244), .c(new_n248), .out0(new_n252));
  nanp02aa1n03x5               g157(.a(new_n250), .b(new_n252), .o1(\s[24] ));
  nor042aa1n06x5               g158(.a(new_n249), .b(new_n247), .o1(new_n254));
  nanb03aa1n02x5               g159(.a(new_n224), .b(new_n254), .c(new_n236), .out0(new_n255));
  nanp02aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  nona22aa1n02x4               g161(.a(new_n242), .b(new_n247), .c(new_n249), .out0(new_n257));
  oaib12aa1n03x5               g162(.a(new_n257), .b(new_n251), .c(new_n256), .out0(new_n258));
  aoi013aa1n02x4               g163(.a(new_n258), .b(new_n240), .c(new_n236), .d(new_n254), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n255), .c(new_n192), .d(new_n195), .o1(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  xnrc02aa1n12x5               g166(.a(\b[24] ), .b(\a[25] ), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  norp02aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  tech160nm_fixnrc02aa1n04x5   g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n264), .c(new_n260), .d(new_n263), .o1(new_n266));
  oabi12aa1n02x5               g171(.a(new_n265), .b(\a[25] ), .c(\b[24] ), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n266), .b(new_n267), .c(new_n263), .d(new_n260), .o1(\s[26] ));
  nor042aa1n12x5               g173(.a(new_n265), .b(new_n262), .o1(new_n269));
  nano32aa1d15x5               g174(.a(new_n224), .b(new_n269), .c(new_n236), .d(new_n254), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n200), .c(new_n140), .d(new_n191), .o1(new_n271));
  nano22aa1n03x5               g176(.a(new_n226), .b(new_n236), .c(new_n254), .out0(new_n272));
  inv000aa1d42x5               g177(.a(\a[26] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(\b[25] ), .o1(new_n274));
  oao003aa1n02x5               g179(.a(new_n273), .b(new_n274), .c(new_n264), .carry(new_n275));
  oaoi13aa1n09x5               g180(.a(new_n275), .b(new_n269), .c(new_n272), .d(new_n258), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  xnbna2aa1n06x5               g182(.a(new_n277), .b(new_n276), .c(new_n271), .out0(\s[27] ));
  aobi12aa1n06x5               g183(.a(new_n277), .b(new_n276), .c(new_n271), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n270), .o1(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n192), .c(new_n195), .o1(new_n281));
  aboi22aa1n03x5               g186(.a(new_n251), .b(new_n256), .c(new_n254), .d(new_n242), .out0(new_n282));
  nanp03aa1n02x5               g187(.a(new_n240), .b(new_n236), .c(new_n254), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n269), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n275), .o1(new_n285));
  aoai13aa1n09x5               g190(.a(new_n285), .b(new_n284), .c(new_n283), .d(new_n282), .o1(new_n286));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  oaoi13aa1n03x5               g192(.a(new_n287), .b(new_n277), .c(new_n281), .d(new_n286), .o1(new_n288));
  xorc02aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .out0(new_n289));
  inv000aa1d42x5               g194(.a(\a[27] ), .o1(new_n290));
  oaib12aa1n02x5               g195(.a(new_n289), .b(\b[26] ), .c(new_n290), .out0(new_n291));
  oai022aa1n03x5               g196(.a(new_n288), .b(new_n289), .c(new_n291), .d(new_n279), .o1(\s[28] ));
  xorc02aa1n12x5               g197(.a(\a[29] ), .b(\b[28] ), .out0(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  inv000aa1d42x5               g199(.a(\a[28] ), .o1(new_n295));
  xroi22aa1d04x5               g200(.a(new_n290), .b(\b[26] ), .c(new_n295), .d(\b[27] ), .out0(new_n296));
  inv000aa1d42x5               g201(.a(new_n296), .o1(new_n297));
  inv000aa1d42x5               g202(.a(\b[27] ), .o1(new_n298));
  oao003aa1n06x5               g203(.a(new_n295), .b(new_n298), .c(new_n287), .carry(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  aoai13aa1n04x5               g205(.a(new_n300), .b(new_n297), .c(new_n276), .d(new_n271), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n301), .b(new_n294), .o1(new_n302));
  nand42aa1n04x5               g207(.a(new_n192), .b(new_n195), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n296), .b(new_n286), .c(new_n303), .d(new_n270), .o1(new_n304));
  nona22aa1n02x5               g209(.a(new_n304), .b(new_n299), .c(new_n294), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n302), .b(new_n305), .o1(\s[29] ));
  xorb03aa1n02x5               g211(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g212(.a(new_n294), .b(new_n277), .c(new_n289), .out0(new_n308));
  aoai13aa1n06x5               g213(.a(new_n308), .b(new_n286), .c(new_n303), .d(new_n270), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n310));
  xorc02aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .out0(new_n311));
  oai012aa1n02x5               g216(.a(new_n311), .b(\b[28] ), .c(\a[29] ), .o1(new_n312));
  aoi012aa1n02x5               g217(.a(new_n312), .b(new_n299), .c(new_n293), .o1(new_n313));
  tech160nm_finand02aa1n03p5x5 g218(.a(new_n309), .b(new_n313), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n311), .c(new_n309), .d(new_n310), .o1(\s[30] ));
  nano32aa1d15x5               g220(.a(new_n294), .b(new_n311), .c(new_n277), .d(new_n289), .out0(new_n316));
  inv000aa1d42x5               g221(.a(new_n316), .o1(new_n317));
  and002aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .o(new_n318));
  norp02aa1n02x5               g223(.a(new_n313), .b(new_n318), .o1(new_n319));
  inv000aa1n02x5               g224(.a(new_n319), .o1(new_n320));
  aoai13aa1n06x5               g225(.a(new_n320), .b(new_n317), .c(new_n276), .d(new_n271), .o1(new_n321));
  xnrc02aa1n02x5               g226(.a(\b[30] ), .b(\a[31] ), .out0(new_n322));
  nanp02aa1n03x5               g227(.a(new_n321), .b(new_n322), .o1(new_n323));
  aoai13aa1n03x5               g228(.a(new_n316), .b(new_n286), .c(new_n303), .d(new_n270), .o1(new_n324));
  nona22aa1n02x5               g229(.a(new_n324), .b(new_n319), .c(new_n322), .out0(new_n325));
  nanp02aa1n03x5               g230(.a(new_n323), .b(new_n325), .o1(\s[31] ));
  inv000aa1d42x5               g231(.a(new_n105), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n102), .b(new_n106), .c(new_n327), .out0(\s[3] ));
  aoai13aa1n02x5               g233(.a(new_n131), .b(new_n99), .c(new_n101), .d(new_n100), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n130), .b(new_n329), .c(new_n327), .out0(\s[4] ));
  xorb03aa1n02x5               g235(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g236(.a(new_n134), .b(new_n109), .out0(new_n332));
  xobna2aa1n03x5               g237(.a(new_n135), .b(new_n332), .c(new_n137), .out0(\s[6] ));
  aoai13aa1n02x5               g238(.a(new_n121), .b(new_n119), .c(new_n132), .d(new_n108), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  norb02aa1n02x5               g240(.a(new_n111), .b(new_n110), .out0(new_n336));
  inv000aa1d42x5               g241(.a(new_n112), .o1(new_n337));
  nanp03aa1n02x5               g242(.a(new_n334), .b(new_n337), .c(new_n113), .o1(new_n338));
  xnbna2aa1n03x5               g243(.a(new_n336), .b(new_n338), .c(new_n337), .out0(\s[8] ));
  xorb03aa1n02x5               g244(.a(new_n140), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


