// Benchmark "adder" written by ABC on Wed Jul 17 20:53:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n331, new_n332, new_n334, new_n335, new_n337, new_n338, new_n339,
    new_n340, new_n342, new_n344, new_n345, new_n346, new_n347, new_n350,
    new_n351, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor022aa1n16x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand42aa1n06x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nona22aa1n09x5               g005(.a(new_n99), .b(new_n98), .c(new_n100), .out0(new_n101));
  nand42aa1n06x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nor002aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nano22aa1n12x5               g008(.a(new_n103), .b(new_n99), .c(new_n102), .out0(new_n104));
  orn002aa1n24x5               g009(.a(\a[4] ), .b(\b[3] ), .o(new_n105));
  nand02aa1n06x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  oai112aa1n06x5               g011(.a(new_n105), .b(new_n106), .c(\b[2] ), .d(\a[3] ), .o1(new_n107));
  aoi012aa1d24x5               g012(.a(new_n107), .b(new_n104), .c(new_n101), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  oai022aa1d24x5               g014(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n110));
  norb02aa1n03x5               g015(.a(new_n109), .b(new_n110), .out0(new_n111));
  nor042aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  aoi012aa1n12x5               g017(.a(new_n112), .b(\a[4] ), .c(\b[3] ), .o1(new_n113));
  nand42aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  oai012aa1n02x5               g019(.a(new_n114), .b(\b[6] ), .c(\a[7] ), .o1(new_n115));
  tech160nm_finand02aa1n03p5x5 g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nanp02aa1n04x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nano22aa1n03x7               g022(.a(new_n115), .b(new_n116), .c(new_n117), .out0(new_n118));
  nand23aa1n06x5               g023(.a(new_n118), .b(new_n111), .c(new_n113), .o1(new_n119));
  nor042aa1d18x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  oai012aa1n02x5               g025(.a(new_n114), .b(new_n120), .c(new_n112), .o1(new_n121));
  nano22aa1d15x5               g026(.a(new_n120), .b(new_n116), .c(new_n117), .out0(new_n122));
  inv000aa1d42x5               g027(.a(new_n110), .o1(new_n123));
  nanb02aa1n06x5               g028(.a(new_n112), .b(new_n114), .out0(new_n124));
  nor042aa1n03x5               g029(.a(new_n124), .b(new_n123), .o1(new_n125));
  aobi12aa1n12x5               g030(.a(new_n121), .b(new_n125), .c(new_n122), .out0(new_n126));
  oai012aa1d24x5               g031(.a(new_n126), .b(new_n108), .c(new_n119), .o1(new_n127));
  nand42aa1n08x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  aoi012aa1n02x5               g033(.a(new_n97), .b(new_n127), .c(new_n128), .o1(new_n129));
  nor002aa1d32x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n16x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  norb02aa1n02x5               g037(.a(new_n128), .b(new_n97), .out0(new_n133));
  nanp02aa1n02x5               g038(.a(new_n127), .b(new_n133), .o1(new_n134));
  norp02aa1n06x5               g039(.a(new_n130), .b(new_n97), .o1(new_n135));
  nanp03aa1n02x5               g040(.a(new_n134), .b(new_n131), .c(new_n135), .o1(new_n136));
  oai012aa1n02x5               g041(.a(new_n136), .b(new_n129), .c(new_n132), .o1(\s[10] ));
  nano23aa1d15x5               g042(.a(new_n97), .b(new_n130), .c(new_n131), .d(new_n128), .out0(new_n138));
  nanp02aa1n02x5               g043(.a(new_n127), .b(new_n138), .o1(new_n139));
  oai012aa1n02x5               g044(.a(new_n131), .b(new_n130), .c(new_n97), .o1(new_n140));
  nor002aa1d32x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nand42aa1n06x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  norb02aa1n09x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  xnbna2aa1n03x5               g048(.a(new_n143), .b(new_n139), .c(new_n140), .out0(\s[11] ));
  inv040aa1n08x5               g049(.a(new_n141), .o1(new_n145));
  aob012aa1n02x5               g050(.a(new_n143), .b(new_n139), .c(new_n140), .out0(new_n146));
  nor022aa1n16x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand42aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n09x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  nona23aa1n02x4               g054(.a(new_n146), .b(new_n148), .c(new_n147), .d(new_n141), .out0(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n149), .c(new_n146), .d(new_n145), .o1(\s[12] ));
  nand23aa1d12x5               g056(.a(new_n138), .b(new_n143), .c(new_n149), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  nanb03aa1n12x5               g058(.a(new_n147), .b(new_n148), .c(new_n142), .out0(new_n154));
  oaih12aa1n12x5               g059(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .o1(new_n155));
  oaoi03aa1n09x5               g060(.a(\a[12] ), .b(\b[11] ), .c(new_n145), .o1(new_n156));
  inv040aa1n02x5               g061(.a(new_n156), .o1(new_n157));
  oai013aa1n09x5               g062(.a(new_n157), .b(new_n154), .c(new_n135), .d(new_n155), .o1(new_n158));
  nor042aa1d18x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n08x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  aoai13aa1n02x5               g066(.a(new_n161), .b(new_n158), .c(new_n127), .d(new_n153), .o1(new_n162));
  nano22aa1n03x7               g067(.a(new_n147), .b(new_n142), .c(new_n148), .out0(new_n163));
  oab012aa1n02x4               g068(.a(new_n155), .b(new_n97), .c(new_n130), .out0(new_n164));
  aoi112aa1n02x5               g069(.a(new_n156), .b(new_n161), .c(new_n164), .d(new_n163), .o1(new_n165));
  aobi12aa1n02x5               g070(.a(new_n165), .b(new_n127), .c(new_n153), .out0(new_n166));
  norb02aa1n02x5               g071(.a(new_n162), .b(new_n166), .out0(\s[13] ));
  inv030aa1n03x5               g072(.a(new_n159), .o1(new_n168));
  nor002aa1n04x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand42aa1n08x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  nona23aa1n02x4               g076(.a(new_n162), .b(new_n170), .c(new_n169), .d(new_n159), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n172), .b(new_n171), .c(new_n168), .d(new_n162), .o1(\s[14] ));
  nano23aa1d15x5               g078(.a(new_n159), .b(new_n169), .c(new_n170), .d(new_n160), .out0(new_n174));
  nand03aa1n02x5               g079(.a(new_n127), .b(new_n153), .c(new_n174), .o1(new_n175));
  aoai13aa1n03x5               g080(.a(new_n174), .b(new_n156), .c(new_n164), .d(new_n163), .o1(new_n176));
  oaoi03aa1n12x5               g081(.a(\a[14] ), .b(\b[13] ), .c(new_n168), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(new_n176), .b(new_n178), .o1(new_n179));
  xorc02aa1n12x5               g084(.a(\a[15] ), .b(\b[14] ), .out0(new_n180));
  oaib12aa1n02x5               g085(.a(new_n180), .b(new_n179), .c(new_n175), .out0(new_n181));
  aoi112aa1n02x5               g086(.a(new_n180), .b(new_n177), .c(new_n158), .d(new_n174), .o1(new_n182));
  aobi12aa1n02x5               g087(.a(new_n181), .b(new_n182), .c(new_n175), .out0(\s[15] ));
  nor042aa1n06x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n184), .o1(new_n185));
  xorc02aa1n12x5               g090(.a(\a[16] ), .b(\b[15] ), .out0(new_n186));
  and002aa1n02x5               g091(.a(\b[15] ), .b(\a[16] ), .o(new_n187));
  oai022aa1n02x5               g092(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n188));
  nona22aa1n03x5               g093(.a(new_n181), .b(new_n187), .c(new_n188), .out0(new_n189));
  aoai13aa1n02x5               g094(.a(new_n189), .b(new_n186), .c(new_n181), .d(new_n185), .o1(\s[16] ));
  and002aa1n18x5               g095(.a(new_n186), .b(new_n180), .o(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n177), .c(new_n158), .d(new_n174), .o1(new_n192));
  nano32aa1d12x5               g097(.a(new_n152), .b(new_n186), .c(new_n174), .d(new_n180), .out0(new_n193));
  nand02aa1d08x5               g098(.a(new_n127), .b(new_n193), .o1(new_n194));
  tech160nm_fioaoi03aa1n03p5x5 g099(.a(\a[16] ), .b(\b[15] ), .c(new_n185), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  nand23aa1d12x5               g101(.a(new_n194), .b(new_n192), .c(new_n196), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  aoi112aa1n02x5               g103(.a(new_n198), .b(new_n195), .c(new_n127), .d(new_n193), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n197), .b(new_n198), .c(new_n199), .d(new_n192), .o1(\s[17] ));
  nor002aa1n03x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  nor022aa1n08x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand42aa1n06x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nanb02aa1n06x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  aoai13aa1n02x5               g109(.a(new_n204), .b(new_n201), .c(new_n197), .d(new_n198), .o1(new_n205));
  nona22aa1n02x4               g110(.a(new_n203), .b(new_n202), .c(new_n201), .out0(new_n206));
  aoai13aa1n02x5               g111(.a(new_n205), .b(new_n206), .c(new_n198), .d(new_n197), .o1(\s[18] ));
  norb02aa1n06x5               g112(.a(new_n198), .b(new_n204), .out0(new_n208));
  oa0012aa1n02x5               g113(.a(new_n203), .b(new_n202), .c(new_n201), .o(new_n209));
  xorc02aa1n12x5               g114(.a(\a[19] ), .b(\b[18] ), .out0(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n209), .c(new_n197), .d(new_n208), .o1(new_n211));
  aoi112aa1n02x5               g116(.a(new_n210), .b(new_n209), .c(new_n197), .d(new_n208), .o1(new_n212));
  norb02aa1n03x4               g117(.a(new_n211), .b(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g119(.a(\a[19] ), .o1(new_n215));
  inv000aa1d42x5               g120(.a(\b[18] ), .o1(new_n216));
  nand02aa1n03x5               g121(.a(new_n216), .b(new_n215), .o1(new_n217));
  nor042aa1n02x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand42aa1n04x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  norb02aa1n03x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  nano22aa1n02x4               g125(.a(new_n218), .b(new_n217), .c(new_n219), .out0(new_n221));
  nanp02aa1n03x5               g126(.a(new_n211), .b(new_n221), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n222), .b(new_n220), .c(new_n217), .d(new_n211), .o1(\s[20] ));
  and003aa1n06x5               g128(.a(new_n208), .b(new_n220), .c(new_n210), .o(new_n224));
  nanp02aa1n02x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  nano22aa1n03x7               g130(.a(new_n218), .b(new_n225), .c(new_n219), .out0(new_n226));
  tech160nm_fioai012aa1n03p5x5 g131(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .o1(new_n227));
  oab012aa1n06x5               g132(.a(new_n227), .b(new_n201), .c(new_n202), .out0(new_n228));
  oaoi03aa1n02x5               g133(.a(\a[20] ), .b(\b[19] ), .c(new_n217), .o1(new_n229));
  tech160nm_fiao0012aa1n02p5x5 g134(.a(new_n229), .b(new_n228), .c(new_n226), .o(new_n230));
  nor042aa1n09x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  nand42aa1n03x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n230), .c(new_n197), .d(new_n224), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n229), .b(new_n233), .c(new_n228), .d(new_n226), .o1(new_n235));
  aobi12aa1n02x5               g140(.a(new_n235), .b(new_n197), .c(new_n224), .out0(new_n236));
  norb02aa1n03x4               g141(.a(new_n234), .b(new_n236), .out0(\s[21] ));
  inv000aa1d42x5               g142(.a(new_n231), .o1(new_n238));
  nor042aa1n03x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nand42aa1n04x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  norb03aa1n02x5               g146(.a(new_n240), .b(new_n231), .c(new_n239), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n234), .b(new_n242), .o1(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n241), .c(new_n238), .d(new_n234), .o1(\s[22] ));
  nano23aa1n09x5               g149(.a(new_n231), .b(new_n239), .c(new_n240), .d(new_n232), .out0(new_n245));
  inv020aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  nano32aa1n02x4               g151(.a(new_n246), .b(new_n208), .c(new_n210), .d(new_n220), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n245), .b(new_n229), .c(new_n228), .d(new_n226), .o1(new_n248));
  oai012aa1n12x5               g153(.a(new_n240), .b(new_n239), .c(new_n231), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(new_n248), .b(new_n249), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n250), .c(new_n197), .d(new_n247), .o1(new_n252));
  nanb02aa1n02x5               g157(.a(new_n251), .b(new_n249), .out0(new_n253));
  aoi122aa1n06x5               g158(.a(new_n253), .b(new_n230), .c(new_n245), .d(new_n197), .e(new_n247), .o1(new_n254));
  norb02aa1n02x7               g159(.a(new_n252), .b(new_n254), .out0(\s[23] ));
  norp02aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  tech160nm_fixorc02aa1n05x5   g162(.a(\a[24] ), .b(\b[23] ), .out0(new_n258));
  oai022aa1n02x5               g163(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n259));
  aoi012aa1n02x5               g164(.a(new_n259), .b(\a[24] ), .c(\b[23] ), .o1(new_n260));
  nanp02aa1n03x5               g165(.a(new_n252), .b(new_n260), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n258), .c(new_n257), .d(new_n252), .o1(\s[24] ));
  nano22aa1n06x5               g167(.a(new_n246), .b(new_n251), .c(new_n258), .out0(new_n263));
  and002aa1n02x5               g168(.a(new_n224), .b(new_n263), .o(new_n264));
  and002aa1n02x5               g169(.a(new_n258), .b(new_n251), .o(new_n265));
  inv020aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  aob012aa1n02x5               g171(.a(new_n259), .b(\b[23] ), .c(\a[24] ), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n266), .c(new_n248), .d(new_n249), .o1(new_n268));
  tech160nm_fixorc02aa1n03p5x5 g173(.a(\a[25] ), .b(\b[24] ), .out0(new_n269));
  aoai13aa1n09x5               g174(.a(new_n269), .b(new_n268), .c(new_n197), .d(new_n264), .o1(new_n270));
  nanb02aa1n02x5               g175(.a(new_n269), .b(new_n267), .out0(new_n271));
  aoi122aa1n06x5               g176(.a(new_n271), .b(new_n250), .c(new_n265), .d(new_n197), .e(new_n264), .o1(new_n272));
  norb02aa1n02x7               g177(.a(new_n270), .b(new_n272), .out0(\s[25] ));
  norp02aa1n02x5               g178(.a(\b[24] ), .b(\a[25] ), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n274), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .out0(new_n276));
  nanp02aa1n02x5               g181(.a(\b[25] ), .b(\a[26] ), .o1(new_n277));
  oai022aa1n02x5               g182(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n278));
  norb02aa1n02x5               g183(.a(new_n277), .b(new_n278), .out0(new_n279));
  nanp02aa1n03x5               g184(.a(new_n270), .b(new_n279), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n276), .c(new_n275), .d(new_n270), .o1(\s[26] ));
  and002aa1n02x5               g186(.a(new_n276), .b(new_n269), .o(new_n282));
  nand23aa1n09x5               g187(.a(new_n224), .b(new_n263), .c(new_n282), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  nand42aa1n08x5               g189(.a(new_n197), .b(new_n284), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n191), .o1(new_n286));
  tech160nm_fiaoi012aa1n05x5   g191(.a(new_n286), .b(new_n176), .c(new_n178), .o1(new_n287));
  aoi112aa1n06x5               g192(.a(new_n287), .b(new_n195), .c(new_n127), .d(new_n193), .o1(new_n288));
  aoi022aa1n09x5               g193(.a(new_n268), .b(new_n282), .c(new_n277), .d(new_n278), .o1(new_n289));
  oai012aa1n12x5               g194(.a(new_n289), .b(new_n288), .c(new_n283), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  aoi122aa1n02x5               g196(.a(new_n291), .b(new_n277), .c(new_n278), .d(new_n268), .e(new_n282), .o1(new_n292));
  aoi022aa1n02x5               g197(.a(new_n290), .b(new_n291), .c(new_n292), .d(new_n285), .o1(\s[27] ));
  norp02aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n294), .o1(new_n295));
  nanp02aa1n06x5               g200(.a(new_n290), .b(new_n291), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .out0(new_n297));
  inv000aa1d42x5               g202(.a(new_n291), .o1(new_n298));
  oai022aa1n02x5               g203(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n299));
  aoi012aa1n02x5               g204(.a(new_n299), .b(\a[28] ), .c(\b[27] ), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n298), .c(new_n285), .d(new_n289), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n297), .c(new_n296), .d(new_n295), .o1(\s[28] ));
  and002aa1n06x5               g207(.a(new_n297), .b(new_n291), .o(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  inv000aa1d42x5               g209(.a(\b[27] ), .o1(new_n305));
  oaib12aa1n09x5               g210(.a(new_n299), .b(new_n305), .c(\a[28] ), .out0(new_n306));
  inv000aa1d42x5               g211(.a(new_n306), .o1(new_n307));
  tech160nm_fixorc02aa1n03p5x5 g212(.a(\a[29] ), .b(\b[28] ), .out0(new_n308));
  norb02aa1n02x5               g213(.a(new_n308), .b(new_n307), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n285), .d(new_n289), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n308), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n307), .c(new_n290), .d(new_n303), .o1(new_n312));
  nanp02aa1n03x5               g217(.a(new_n312), .b(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g219(.a(new_n311), .b(new_n291), .c(new_n297), .out0(new_n315));
  oaoi03aa1n02x5               g220(.a(\a[29] ), .b(\b[28] ), .c(new_n306), .o1(new_n316));
  xnrc02aa1n02x5               g221(.a(\b[29] ), .b(\a[30] ), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n316), .c(new_n290), .d(new_n315), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n315), .o1(new_n319));
  norp02aa1n02x5               g224(.a(new_n316), .b(new_n317), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n285), .d(new_n289), .o1(new_n321));
  nanp02aa1n03x5               g226(.a(new_n318), .b(new_n321), .o1(\s[30] ));
  nano32aa1n03x7               g227(.a(new_n317), .b(new_n308), .c(new_n297), .d(new_n291), .out0(new_n323));
  aoi012aa1n02x5               g228(.a(new_n320), .b(\a[30] ), .c(\b[29] ), .o1(new_n324));
  xnrc02aa1n02x5               g229(.a(\b[30] ), .b(\a[31] ), .out0(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n324), .c(new_n290), .d(new_n323), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n323), .o1(new_n327));
  norp02aa1n02x5               g232(.a(new_n324), .b(new_n325), .o1(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n327), .c(new_n285), .d(new_n289), .o1(new_n329));
  nanp02aa1n03x5               g234(.a(new_n326), .b(new_n329), .o1(\s[31] ));
  nanb02aa1n02x5               g235(.a(new_n103), .b(new_n102), .out0(new_n331));
  oai012aa1n02x5               g236(.a(new_n99), .b(new_n98), .c(new_n100), .o1(new_n332));
  aoi022aa1n02x5               g237(.a(new_n104), .b(new_n101), .c(new_n332), .d(new_n331), .o1(\s[3] ));
  inv000aa1d42x5               g238(.a(new_n108), .o1(new_n334));
  aoi012aa1n02x5               g239(.a(new_n103), .b(new_n104), .c(new_n101), .o1(new_n335));
  aoai13aa1n02x5               g240(.a(new_n334), .b(new_n335), .c(new_n106), .d(new_n105), .o1(\s[4] ));
  norp02aa1n04x5               g241(.a(\b[4] ), .b(\a[5] ), .o1(new_n337));
  nona23aa1n03x5               g242(.a(new_n106), .b(new_n109), .c(new_n108), .d(new_n337), .out0(new_n338));
  inv000aa1d42x5               g243(.a(new_n337), .o1(new_n339));
  aboi22aa1n03x5               g244(.a(new_n108), .b(new_n106), .c(new_n339), .d(new_n109), .out0(new_n340));
  norb02aa1n02x5               g245(.a(new_n338), .b(new_n340), .out0(\s[5] ));
  xorc02aa1n02x5               g246(.a(\a[6] ), .b(\b[5] ), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n342), .b(new_n338), .c(new_n339), .out0(\s[6] ));
  nand23aa1n03x5               g248(.a(new_n338), .b(new_n339), .c(new_n342), .o1(new_n344));
  nanp02aa1n03x5               g249(.a(new_n344), .b(new_n122), .o1(new_n345));
  inv000aa1d42x5               g250(.a(new_n120), .o1(new_n346));
  aoi022aa1n02x5               g251(.a(new_n344), .b(new_n117), .c(new_n346), .d(new_n116), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n345), .b(new_n347), .out0(\s[7] ));
  xobna2aa1n03x5               g253(.a(new_n124), .b(new_n345), .c(new_n346), .out0(\s[8] ));
  norp02aa1n02x5               g254(.a(new_n108), .b(new_n119), .o1(new_n350));
  oaib12aa1n02x5               g255(.a(new_n121), .b(new_n97), .c(new_n128), .out0(new_n351));
  aoi012aa1n02x5               g256(.a(new_n351), .b(new_n125), .c(new_n122), .o1(new_n352));
  aboi22aa1n03x5               g257(.a(new_n350), .b(new_n352), .c(new_n127), .d(new_n133), .out0(\s[9] ));
endmodule


