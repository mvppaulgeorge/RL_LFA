// Benchmark "adder" written by ABC on Thu Jul 18 15:07:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n307, new_n310, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[6] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[5] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[4] ), .b(\a[5] ), .o1(new_n102));
  oao003aa1n03x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .carry(new_n103));
  nor042aa1n02x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  nand22aa1n12x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nor042aa1n12x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  nand22aa1n09x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nano23aa1n06x5               g012(.a(new_n104), .b(new_n106), .c(new_n107), .d(new_n105), .out0(new_n108));
  inv000aa1n02x5               g013(.a(new_n106), .o1(new_n109));
  oaoi03aa1n03x5               g014(.a(\a[8] ), .b(\b[7] ), .c(new_n109), .o1(new_n110));
  tech160nm_fiaoi012aa1n03p5x5 g015(.a(new_n110), .b(new_n108), .c(new_n103), .o1(new_n111));
  nor042aa1d18x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  inv000aa1n02x5               g017(.a(new_n112), .o1(new_n113));
  oao003aa1n06x5               g018(.a(\a[4] ), .b(\b[3] ), .c(new_n113), .carry(new_n114));
  tech160nm_fixorc02aa1n02p5x5 g019(.a(\a[4] ), .b(\b[3] ), .out0(new_n115));
  nand42aa1n04x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  norb02aa1n03x5               g021(.a(new_n116), .b(new_n112), .out0(new_n117));
  and002aa1n12x5               g022(.a(\b[1] ), .b(\a[2] ), .o(new_n118));
  nand22aa1n12x5               g023(.a(\b[0] ), .b(\a[1] ), .o1(new_n119));
  nor042aa1n03x5               g024(.a(\b[1] ), .b(\a[2] ), .o1(new_n120));
  oab012aa1n09x5               g025(.a(new_n118), .b(new_n120), .c(new_n119), .out0(new_n121));
  nand03aa1n06x5               g026(.a(new_n121), .b(new_n115), .c(new_n117), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[6] ), .b(\b[5] ), .out0(new_n123));
  nand02aa1d06x5               g028(.a(\b[4] ), .b(\a[5] ), .o1(new_n124));
  norb02aa1n03x5               g029(.a(new_n124), .b(new_n102), .out0(new_n125));
  nand03aa1n02x5               g030(.a(new_n108), .b(new_n123), .c(new_n125), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n111), .b(new_n126), .c(new_n122), .d(new_n114), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  nanp02aa1n02x5               g033(.a(new_n127), .b(new_n128), .o1(new_n129));
  nor042aa1n06x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand02aa1n06x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nanb02aa1d24x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  xobna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  norb02aa1n02x5               g038(.a(new_n128), .b(new_n132), .out0(new_n134));
  aoai13aa1n02x5               g039(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n135));
  aob012aa1n03x5               g040(.a(new_n135), .b(new_n127), .c(new_n134), .out0(new_n136));
  xorb03aa1n02x5               g041(.a(new_n136), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n12x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand42aa1d28x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  aoi012aa1n02x5               g044(.a(new_n138), .b(new_n136), .c(new_n139), .o1(new_n140));
  xnrb03aa1n03x5               g045(.a(new_n140), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1n08x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand42aa1n16x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nona23aa1n03x5               g048(.a(new_n143), .b(new_n139), .c(new_n138), .d(new_n142), .out0(new_n144));
  oa0012aa1n06x5               g049(.a(new_n143), .b(new_n142), .c(new_n138), .o(new_n145));
  oabi12aa1n06x5               g050(.a(new_n145), .b(new_n135), .c(new_n144), .out0(new_n146));
  nano23aa1d15x5               g051(.a(new_n138), .b(new_n142), .c(new_n143), .d(new_n139), .out0(new_n147));
  nanb03aa1d24x5               g052(.a(new_n132), .b(new_n147), .c(new_n128), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  xnrc02aa1n12x5               g054(.a(\b[12] ), .b(\a[13] ), .out0(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n146), .c(new_n127), .d(new_n149), .o1(new_n152));
  aoi112aa1n02x5               g057(.a(new_n146), .b(new_n151), .c(new_n127), .d(new_n149), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n152), .b(new_n153), .out0(\s[13] ));
  norp02aa1n02x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  inv000aa1n03x5               g060(.a(new_n155), .o1(new_n156));
  tech160nm_fixnrc02aa1n04x5   g061(.a(\b[13] ), .b(\a[14] ), .out0(new_n157));
  xobna2aa1n03x5               g062(.a(new_n157), .b(new_n152), .c(new_n156), .out0(\s[14] ));
  nor042aa1n06x5               g063(.a(new_n157), .b(new_n150), .o1(new_n159));
  oaoi03aa1n02x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n160));
  aoi012aa1n06x5               g065(.a(new_n160), .b(new_n146), .c(new_n159), .o1(new_n161));
  nona32aa1n02x4               g066(.a(new_n127), .b(new_n157), .c(new_n150), .d(new_n148), .out0(new_n162));
  xnrc02aa1n12x5               g067(.a(\b[14] ), .b(\a[15] ), .out0(new_n163));
  xobna2aa1n03x5               g068(.a(new_n163), .b(new_n162), .c(new_n161), .out0(\s[15] ));
  nor042aa1n06x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  inv000aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  aoai13aa1n03x5               g071(.a(new_n166), .b(new_n163), .c(new_n162), .d(new_n161), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  inv040aa1d32x5               g073(.a(\a[17] ), .o1(new_n169));
  tech160nm_fixnrc02aa1n02p5x5 g074(.a(\b[15] ), .b(\a[16] ), .out0(new_n170));
  nor002aa1n03x5               g075(.a(new_n170), .b(new_n163), .o1(new_n171));
  nano22aa1d15x5               g076(.a(new_n148), .b(new_n159), .c(new_n171), .out0(new_n172));
  oaoi03aa1n12x5               g077(.a(\a[16] ), .b(\b[15] ), .c(new_n166), .o1(new_n173));
  oaoi03aa1n02x5               g078(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n174));
  aoai13aa1n03x5               g079(.a(new_n159), .b(new_n145), .c(new_n147), .d(new_n174), .o1(new_n175));
  inv000aa1n02x5               g080(.a(new_n160), .o1(new_n176));
  inv000aa1n02x5               g081(.a(new_n171), .o1(new_n177));
  tech160nm_fiaoi012aa1n05x5   g082(.a(new_n177), .b(new_n175), .c(new_n176), .o1(new_n178));
  aoi112aa1n09x5               g083(.a(new_n178), .b(new_n173), .c(new_n127), .d(new_n172), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(new_n169), .out0(\s[17] ));
  oaoi03aa1n03x5               g085(.a(\a[17] ), .b(\b[16] ), .c(new_n179), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g087(.a(\a[18] ), .o1(new_n183));
  xroi22aa1d06x4               g088(.a(new_n169), .b(\b[16] ), .c(new_n183), .d(\b[17] ), .out0(new_n184));
  inv000aa1n03x5               g089(.a(new_n184), .o1(new_n185));
  oaih22aa1n04x5               g090(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n186));
  oaib12aa1n09x5               g091(.a(new_n186), .b(new_n183), .c(\b[17] ), .out0(new_n187));
  tech160nm_fioai012aa1n05x5   g092(.a(new_n187), .b(new_n179), .c(new_n185), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g094(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n09x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nand42aa1n06x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  nor042aa1n06x5               g099(.a(\b[19] ), .b(\a[20] ), .o1(new_n195));
  nand42aa1n08x5               g100(.a(\b[19] ), .b(\a[20] ), .o1(new_n196));
  nanb02aa1n02x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  aoai13aa1n03x5               g102(.a(new_n197), .b(new_n191), .c(new_n188), .d(new_n194), .o1(new_n198));
  tech160nm_finand02aa1n03p5x5 g103(.a(new_n127), .b(new_n172), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n173), .o1(new_n200));
  oai112aa1n06x5               g105(.a(new_n199), .b(new_n200), .c(new_n161), .d(new_n177), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(\b[16] ), .b(new_n169), .out0(new_n202));
  oaoi03aa1n02x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n194), .b(new_n203), .c(new_n201), .d(new_n184), .o1(new_n204));
  nona22aa1n03x5               g109(.a(new_n204), .b(new_n197), .c(new_n191), .out0(new_n205));
  nanp02aa1n03x5               g110(.a(new_n198), .b(new_n205), .o1(\s[20] ));
  nona23aa1n09x5               g111(.a(new_n196), .b(new_n192), .c(new_n191), .d(new_n195), .out0(new_n207));
  oa0012aa1n03x5               g112(.a(new_n196), .b(new_n195), .c(new_n191), .o(new_n208));
  inv040aa1n03x5               g113(.a(new_n208), .o1(new_n209));
  oai012aa1d24x5               g114(.a(new_n209), .b(new_n207), .c(new_n187), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  nano23aa1n09x5               g116(.a(new_n191), .b(new_n195), .c(new_n196), .d(new_n192), .out0(new_n212));
  nand22aa1n12x5               g117(.a(new_n184), .b(new_n212), .o1(new_n213));
  tech160nm_fioai012aa1n05x5   g118(.a(new_n211), .b(new_n179), .c(new_n213), .o1(new_n214));
  xorb03aa1n02x5               g119(.a(new_n214), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  xnrc02aa1n12x5               g121(.a(\b[20] ), .b(\a[21] ), .out0(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  tech160nm_fixnrc02aa1n05x5   g123(.a(\b[21] ), .b(\a[22] ), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n216), .c(new_n214), .d(new_n218), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n213), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n218), .b(new_n210), .c(new_n201), .d(new_n221), .o1(new_n222));
  nona22aa1n02x4               g127(.a(new_n222), .b(new_n219), .c(new_n216), .out0(new_n223));
  nanp02aa1n03x5               g128(.a(new_n220), .b(new_n223), .o1(\s[22] ));
  nor042aa1n06x5               g129(.a(new_n219), .b(new_n217), .o1(new_n225));
  inv040aa1d32x5               g130(.a(\a[22] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\b[21] ), .o1(new_n227));
  oao003aa1n06x5               g132(.a(new_n226), .b(new_n227), .c(new_n216), .carry(new_n228));
  aoi012aa1d18x5               g133(.a(new_n228), .b(new_n210), .c(new_n225), .o1(new_n229));
  nano22aa1n02x4               g134(.a(new_n185), .b(new_n225), .c(new_n212), .out0(new_n230));
  inv000aa1n02x5               g135(.a(new_n230), .o1(new_n231));
  tech160nm_fioai012aa1n05x5   g136(.a(new_n229), .b(new_n179), .c(new_n231), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  xorc02aa1n12x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[23] ), .b(\a[24] ), .out0(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n234), .c(new_n232), .d(new_n235), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n229), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n235), .b(new_n238), .c(new_n201), .d(new_n230), .o1(new_n239));
  nona22aa1n02x4               g144(.a(new_n239), .b(new_n236), .c(new_n234), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n237), .b(new_n240), .o1(\s[24] ));
  norb02aa1n02x7               g146(.a(new_n235), .b(new_n236), .out0(new_n242));
  inv020aa1n06x5               g147(.a(new_n242), .o1(new_n243));
  nano32aa1n03x5               g148(.a(new_n243), .b(new_n184), .c(new_n225), .d(new_n212), .out0(new_n244));
  inv020aa1n02x5               g149(.a(new_n244), .o1(new_n245));
  aoai13aa1n06x5               g150(.a(new_n225), .b(new_n208), .c(new_n212), .d(new_n203), .o1(new_n246));
  inv030aa1n02x5               g151(.a(new_n228), .o1(new_n247));
  oai022aa1n02x5               g152(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n248));
  aob012aa1n02x5               g153(.a(new_n248), .b(\b[23] ), .c(\a[24] ), .out0(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n243), .c(new_n246), .d(new_n247), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  tech160nm_fioai012aa1n05x5   g156(.a(new_n251), .b(new_n179), .c(new_n245), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g158(.a(\b[24] ), .b(\a[25] ), .o1(new_n254));
  xorc02aa1n03x5               g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  xnrc02aa1n12x5               g160(.a(\b[25] ), .b(\a[26] ), .out0(new_n256));
  aoai13aa1n03x5               g161(.a(new_n256), .b(new_n254), .c(new_n252), .d(new_n255), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n255), .b(new_n250), .c(new_n201), .d(new_n244), .o1(new_n258));
  nona22aa1n02x4               g163(.a(new_n258), .b(new_n256), .c(new_n254), .out0(new_n259));
  nanp02aa1n03x5               g164(.a(new_n257), .b(new_n259), .o1(\s[26] ));
  nanp02aa1n02x5               g165(.a(\b[25] ), .b(\a[26] ), .o1(new_n261));
  norb02aa1n06x5               g166(.a(new_n255), .b(new_n256), .out0(new_n262));
  oai022aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n263));
  aoi022aa1n09x5               g168(.a(new_n250), .b(new_n262), .c(new_n261), .d(new_n263), .o1(new_n264));
  nano23aa1n06x5               g169(.a(new_n213), .b(new_n243), .c(new_n262), .d(new_n225), .out0(new_n265));
  inv020aa1n03x5               g170(.a(new_n265), .o1(new_n266));
  tech160nm_fioai012aa1n05x5   g171(.a(new_n264), .b(new_n179), .c(new_n266), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g173(.a(\b[26] ), .b(\a[27] ), .o1(new_n269));
  xorc02aa1n02x5               g174(.a(\a[27] ), .b(\b[26] ), .out0(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[27] ), .b(\a[28] ), .out0(new_n271));
  aoai13aa1n03x5               g176(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n270), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n242), .b(new_n228), .c(new_n210), .d(new_n225), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n262), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(new_n263), .b(new_n261), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n275), .b(new_n274), .c(new_n273), .d(new_n249), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n270), .b(new_n276), .c(new_n201), .d(new_n265), .o1(new_n277));
  nona22aa1n02x4               g182(.a(new_n277), .b(new_n271), .c(new_n269), .out0(new_n278));
  nanp02aa1n03x5               g183(.a(new_n272), .b(new_n278), .o1(\s[28] ));
  norb02aa1n02x5               g184(.a(new_n270), .b(new_n271), .out0(new_n280));
  aoai13aa1n02x5               g185(.a(new_n280), .b(new_n276), .c(new_n201), .d(new_n265), .o1(new_n281));
  inv000aa1n03x5               g186(.a(new_n269), .o1(new_n282));
  oaoi03aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .o1(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[28] ), .b(\a[29] ), .out0(new_n284));
  nona22aa1n02x4               g189(.a(new_n281), .b(new_n283), .c(new_n284), .out0(new_n285));
  aoai13aa1n03x5               g190(.a(new_n284), .b(new_n283), .c(new_n267), .d(new_n280), .o1(new_n286));
  nanp02aa1n03x5               g191(.a(new_n286), .b(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n119), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g193(.a(new_n270), .b(new_n284), .c(new_n271), .out0(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .carry(new_n290));
  oaoi03aa1n02x5               g195(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .o1(new_n291));
  tech160nm_fixorc02aa1n03p5x5 g196(.a(\a[30] ), .b(\b[29] ), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n291), .c(new_n267), .d(new_n289), .o1(new_n294));
  aoai13aa1n02x5               g199(.a(new_n289), .b(new_n276), .c(new_n201), .d(new_n265), .o1(new_n295));
  nona22aa1n03x5               g200(.a(new_n295), .b(new_n291), .c(new_n293), .out0(new_n296));
  nanp02aa1n03x5               g201(.a(new_n294), .b(new_n296), .o1(\s[30] ));
  nanp02aa1n02x5               g202(.a(new_n291), .b(new_n292), .o1(new_n298));
  oai012aa1n02x5               g203(.a(new_n298), .b(\b[29] ), .c(\a[30] ), .o1(new_n299));
  nano23aa1n03x7               g204(.a(new_n284), .b(new_n271), .c(new_n292), .d(new_n270), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n276), .c(new_n201), .d(new_n265), .o1(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[30] ), .b(\a[31] ), .out0(new_n302));
  nona22aa1n03x5               g207(.a(new_n301), .b(new_n302), .c(new_n299), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n302), .b(new_n299), .c(new_n267), .d(new_n300), .o1(new_n304));
  nanp02aa1n03x5               g209(.a(new_n304), .b(new_n303), .o1(\s[31] ));
  xobna2aa1n03x5               g210(.a(new_n121), .b(new_n116), .c(new_n113), .out0(\s[3] ));
  oai012aa1n02x5               g211(.a(new_n116), .b(new_n121), .c(new_n112), .o1(new_n307));
  xnrb03aa1n02x5               g212(.a(new_n307), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnbna2aa1n03x5               g213(.a(new_n125), .b(new_n122), .c(new_n114), .out0(\s[5] ));
  nanp03aa1n02x5               g214(.a(new_n122), .b(new_n114), .c(new_n125), .o1(new_n310));
  xobna2aa1n03x5               g215(.a(new_n123), .b(new_n310), .c(new_n124), .out0(\s[6] ));
  norb02aa1n02x5               g216(.a(new_n107), .b(new_n106), .out0(new_n312));
  nanp02aa1n02x5               g217(.a(new_n310), .b(new_n124), .o1(new_n313));
  nanp02aa1n02x5               g218(.a(new_n313), .b(new_n123), .o1(new_n314));
  oai112aa1n02x5               g219(.a(new_n314), .b(new_n312), .c(new_n101), .d(new_n100), .o1(new_n315));
  oaoi13aa1n02x5               g220(.a(new_n312), .b(new_n314), .c(new_n100), .d(new_n101), .o1(new_n316));
  norb02aa1n02x5               g221(.a(new_n315), .b(new_n316), .out0(\s[7] ));
  norb02aa1n02x5               g222(.a(new_n105), .b(new_n104), .out0(new_n318));
  xnbna2aa1n03x5               g223(.a(new_n318), .b(new_n315), .c(new_n109), .out0(\s[8] ));
  xorb03aa1n02x5               g224(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


