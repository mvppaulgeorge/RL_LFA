// Benchmark "adder" written by ABC on Thu Jul 18 02:24:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n331,
    new_n334, new_n335, new_n337, new_n338, new_n339, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d28x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\b[8] ), .o1(new_n98));
  orn002aa1n12x5               g003(.a(\a[3] ), .b(\b[2] ), .o(new_n99));
  oao003aa1n03x5               g004(.a(\a[4] ), .b(\b[3] ), .c(new_n99), .carry(new_n100));
  nand42aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanp03aa1n03x5               g007(.a(new_n99), .b(new_n101), .c(new_n102), .o1(new_n103));
  xnrc02aa1n12x5               g008(.a(\b[3] ), .b(\a[4] ), .out0(new_n104));
  nanp02aa1n04x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  norb03aa1n03x5               g011(.a(new_n101), .b(new_n106), .c(new_n105), .out0(new_n107));
  oai013aa1n06x5               g012(.a(new_n100), .b(new_n103), .c(new_n107), .d(new_n104), .o1(new_n108));
  xnrc02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .out0(new_n109));
  xnrc02aa1n02x5               g014(.a(\b[4] ), .b(\a[5] ), .out0(new_n110));
  nor022aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand22aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n03x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  nor043aa1n03x5               g020(.a(new_n115), .b(new_n110), .c(new_n109), .o1(new_n116));
  inv040aa1d32x5               g021(.a(\a[6] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\b[5] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(new_n118), .b(new_n117), .o1(new_n119));
  aoi112aa1n03x5               g024(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n120));
  norb02aa1n09x5               g025(.a(new_n119), .b(new_n120), .out0(new_n121));
  tech160nm_fiao0012aa1n02p5x5 g026(.a(new_n111), .b(new_n113), .c(new_n112), .o(new_n122));
  oabi12aa1n18x5               g027(.a(new_n122), .b(new_n115), .c(new_n121), .out0(new_n123));
  inv000aa1d42x5               g028(.a(new_n123), .o1(new_n124));
  aob012aa1d15x5               g029(.a(new_n124), .b(new_n108), .c(new_n116), .out0(new_n125));
  oaoi03aa1n02x5               g030(.a(new_n97), .b(new_n98), .c(new_n125), .o1(new_n126));
  xnrb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  tech160nm_fixnrc02aa1n04x5   g032(.a(\b[8] ), .b(\a[9] ), .out0(new_n128));
  nor002aa1d32x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nanb02aa1n06x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  nona22aa1n03x5               g036(.a(new_n125), .b(new_n128), .c(new_n131), .out0(new_n132));
  aoai13aa1n12x5               g037(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n133));
  nor002aa1n16x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1d28x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n132), .c(new_n133), .out0(\s[11] ));
  nanp02aa1n03x5               g042(.a(new_n132), .b(new_n133), .o1(new_n138));
  norp02aa1n24x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand02aa1d28x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n134), .c(new_n138), .d(new_n135), .o1(new_n142));
  aoi112aa1n02x5               g047(.a(new_n134), .b(new_n141), .c(new_n138), .d(new_n135), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(\s[12] ));
  nano23aa1d15x5               g049(.a(new_n134), .b(new_n139), .c(new_n140), .d(new_n135), .out0(new_n145));
  nona22aa1d30x5               g050(.a(new_n145), .b(new_n128), .c(new_n131), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  aoai13aa1n02x5               g052(.a(new_n147), .b(new_n123), .c(new_n108), .d(new_n116), .o1(new_n148));
  nona23aa1d18x5               g053(.a(new_n140), .b(new_n135), .c(new_n134), .d(new_n139), .out0(new_n149));
  aoi012aa1d18x5               g054(.a(new_n139), .b(new_n134), .c(new_n140), .o1(new_n150));
  oai012aa1d24x5               g055(.a(new_n150), .b(new_n149), .c(new_n133), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nor022aa1n06x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanp02aa1n04x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(new_n155));
  xobna2aa1n03x5               g060(.a(new_n155), .b(new_n148), .c(new_n152), .out0(\s[13] ));
  nanp02aa1n02x5               g061(.a(new_n148), .b(new_n152), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n153), .b(new_n157), .c(new_n154), .o1(new_n158));
  xnrb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n02x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand02aa1n03x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nona23aa1n02x4               g066(.a(new_n161), .b(new_n154), .c(new_n153), .d(new_n160), .out0(new_n162));
  nona22aa1n02x4               g067(.a(new_n125), .b(new_n146), .c(new_n162), .out0(new_n163));
  nano23aa1n06x5               g068(.a(new_n153), .b(new_n160), .c(new_n161), .d(new_n154), .out0(new_n164));
  oai012aa1n02x7               g069(.a(new_n161), .b(new_n160), .c(new_n153), .o1(new_n165));
  inv000aa1n02x5               g070(.a(new_n165), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n166), .b(new_n151), .c(new_n164), .o1(new_n167));
  xnrc02aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .out0(new_n168));
  tech160nm_fiaoi012aa1n04x5   g073(.a(new_n168), .b(new_n163), .c(new_n167), .o1(new_n169));
  oaoi13aa1n06x5               g074(.a(new_n162), .b(new_n150), .c(new_n149), .d(new_n133), .o1(new_n170));
  nano22aa1n02x4               g075(.a(new_n170), .b(new_n165), .c(new_n168), .out0(new_n171));
  aoi012aa1n02x5               g076(.a(new_n169), .b(new_n163), .c(new_n171), .o1(\s[15] ));
  nor002aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  xnrc02aa1n12x5               g078(.a(\b[15] ), .b(\a[16] ), .out0(new_n174));
  oai012aa1n02x5               g079(.a(new_n174), .b(new_n169), .c(new_n173), .o1(new_n175));
  orn003aa1n03x7               g080(.a(new_n169), .b(new_n173), .c(new_n174), .o(new_n176));
  nanp02aa1n02x5               g081(.a(new_n176), .b(new_n175), .o1(\s[16] ));
  nor042aa1n09x5               g082(.a(new_n174), .b(new_n168), .o1(new_n178));
  nano22aa1d15x5               g083(.a(new_n146), .b(new_n178), .c(new_n164), .out0(new_n179));
  aoai13aa1n12x5               g084(.a(new_n179), .b(new_n123), .c(new_n108), .d(new_n116), .o1(new_n180));
  aoai13aa1n09x5               g085(.a(new_n178), .b(new_n166), .c(new_n151), .d(new_n164), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[16] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[15] ), .o1(new_n183));
  oaoi03aa1n12x5               g088(.a(new_n182), .b(new_n183), .c(new_n173), .o1(new_n184));
  nand23aa1d12x5               g089(.a(new_n180), .b(new_n181), .c(new_n184), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nand02aa1d28x5               g091(.a(\b[17] ), .b(\a[18] ), .o1(new_n187));
  nor042aa1d18x5               g092(.a(\b[17] ), .b(\a[18] ), .o1(new_n188));
  nanb02aa1n02x5               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  nor042aa1d18x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nand42aa1n03x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  oai012aa1n02x5               g096(.a(new_n191), .b(new_n185), .c(new_n190), .o1(new_n192));
  oai122aa1n03x5               g097(.a(new_n191), .b(new_n185), .c(new_n190), .d(\a[18] ), .e(\b[17] ), .o1(new_n193));
  aboi22aa1n02x7               g098(.a(new_n193), .b(new_n187), .c(new_n189), .d(new_n192), .out0(\s[18] ));
  inv000aa1d42x5               g099(.a(new_n184), .o1(new_n195));
  oaoi13aa1n06x5               g100(.a(new_n195), .b(new_n178), .c(new_n170), .d(new_n166), .o1(new_n196));
  nano23aa1d15x5               g101(.a(new_n188), .b(new_n190), .c(new_n191), .d(new_n187), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  nand22aa1n09x5               g104(.a(new_n190), .b(new_n187), .o1(new_n200));
  oaib12aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n199), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  aoai13aa1n02x7               g107(.a(new_n202), .b(new_n198), .c(new_n196), .d(new_n180), .o1(new_n203));
  nor002aa1d32x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nand02aa1n03x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  norb02aa1n06x4               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  aoi112aa1n03x4               g111(.a(new_n206), .b(new_n201), .c(new_n185), .d(new_n197), .o1(new_n207));
  tech160nm_fiaoi012aa1n02p5x5 g112(.a(new_n207), .b(new_n203), .c(new_n206), .o1(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n04x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nanp02aa1n02x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nanb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  aoai13aa1n02x5               g117(.a(new_n212), .b(new_n204), .c(new_n203), .d(new_n205), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n206), .b(new_n201), .c(new_n185), .d(new_n197), .o1(new_n214));
  nona22aa1n02x5               g119(.a(new_n214), .b(new_n212), .c(new_n204), .out0(new_n215));
  nanp02aa1n03x5               g120(.a(new_n213), .b(new_n215), .o1(\s[20] ));
  nano22aa1n03x7               g121(.a(new_n212), .b(new_n197), .c(new_n206), .out0(new_n217));
  inv030aa1n04x5               g122(.a(new_n217), .o1(new_n218));
  nona22aa1n09x5               g123(.a(new_n200), .b(new_n204), .c(new_n188), .out0(new_n219));
  aoai13aa1n12x5               g124(.a(new_n211), .b(new_n210), .c(new_n219), .d(new_n205), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n220), .b(new_n218), .c(new_n196), .d(new_n180), .o1(new_n221));
  xorb03aa1n03x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  xnrc02aa1n12x5               g128(.a(\b[20] ), .b(\a[21] ), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  tech160nm_fixnrc02aa1n04x5   g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n221), .d(new_n225), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n220), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n225), .b(new_n228), .c(new_n185), .d(new_n217), .o1(new_n229));
  nona22aa1n02x5               g134(.a(new_n229), .b(new_n226), .c(new_n223), .out0(new_n230));
  nanp02aa1n03x5               g135(.a(new_n227), .b(new_n230), .o1(\s[22] ));
  inv000aa1n02x5               g136(.a(new_n133), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n150), .o1(new_n233));
  aoai13aa1n02x5               g138(.a(new_n164), .b(new_n233), .c(new_n145), .d(new_n232), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n178), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n184), .b(new_n235), .c(new_n234), .d(new_n165), .o1(new_n236));
  nor042aa1n06x5               g141(.a(new_n226), .b(new_n224), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  nano23aa1n03x7               g143(.a(new_n238), .b(new_n212), .c(new_n206), .d(new_n197), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n236), .c(new_n125), .d(new_n179), .o1(new_n240));
  orn002aa1n02x5               g145(.a(\a[21] ), .b(\b[20] ), .o(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n241), .o1(new_n242));
  oab012aa1n02x5               g147(.a(new_n242), .b(new_n220), .c(new_n238), .out0(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[22] ), .b(\a[23] ), .out0(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  xnbna2aa1n03x5               g150(.a(new_n245), .b(new_n240), .c(new_n243), .out0(\s[23] ));
  xnrc02aa1n02x5               g151(.a(\b[23] ), .b(\a[24] ), .out0(new_n247));
  nanp02aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  norp02aa1n02x5               g153(.a(new_n220), .b(new_n238), .o1(new_n249));
  nona32aa1n02x4               g154(.a(new_n240), .b(new_n244), .c(new_n242), .d(new_n249), .out0(new_n250));
  nanp02aa1n02x5               g155(.a(new_n250), .b(new_n248), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n243), .o1(new_n252));
  aoi112aa1n06x5               g157(.a(new_n244), .b(new_n252), .c(new_n185), .d(new_n239), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\a[24] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(\b[23] ), .o1(new_n256));
  aoi022aa1n02x5               g161(.a(new_n256), .b(new_n255), .c(\a[23] ), .d(\b[22] ), .o1(new_n257));
  nano22aa1n03x7               g162(.a(new_n253), .b(new_n254), .c(new_n257), .out0(new_n258));
  aoi012aa1n02x7               g163(.a(new_n258), .b(new_n251), .c(new_n247), .o1(\s[24] ));
  nor002aa1n04x5               g164(.a(new_n247), .b(new_n244), .o1(new_n260));
  nano22aa1n03x7               g165(.a(new_n218), .b(new_n237), .c(new_n260), .out0(new_n261));
  aoai13aa1n02x5               g166(.a(new_n261), .b(new_n236), .c(new_n125), .d(new_n179), .o1(new_n262));
  inv020aa1n02x5               g167(.a(new_n261), .o1(new_n263));
  nand22aa1n04x5               g168(.a(new_n260), .b(new_n237), .o1(new_n264));
  norp02aa1n02x5               g169(.a(\b[22] ), .b(\a[23] ), .o1(new_n265));
  oao003aa1n02x5               g170(.a(new_n255), .b(new_n256), .c(new_n265), .carry(new_n266));
  tech160nm_fiaoi012aa1n05x5   g171(.a(new_n266), .b(new_n260), .c(new_n242), .o1(new_n267));
  oai012aa1d24x5               g172(.a(new_n267), .b(new_n220), .c(new_n264), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  aoai13aa1n04x5               g174(.a(new_n269), .b(new_n263), .c(new_n196), .d(new_n180), .o1(new_n270));
  xorc02aa1n06x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  aoi112aa1n02x5               g176(.a(new_n266), .b(new_n271), .c(new_n260), .d(new_n242), .o1(new_n272));
  oa0012aa1n02x5               g177(.a(new_n272), .b(new_n264), .c(new_n220), .o(new_n273));
  aoi022aa1n02x5               g178(.a(new_n270), .b(new_n271), .c(new_n262), .d(new_n273), .o1(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  tech160nm_fixnrc02aa1n04x5   g180(.a(\b[25] ), .b(\a[26] ), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n270), .d(new_n271), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n271), .b(new_n268), .c(new_n185), .d(new_n261), .o1(new_n278));
  nona22aa1n03x5               g183(.a(new_n278), .b(new_n276), .c(new_n275), .out0(new_n279));
  nanp02aa1n03x5               g184(.a(new_n277), .b(new_n279), .o1(\s[26] ));
  norb02aa1n06x5               g185(.a(new_n271), .b(new_n276), .out0(new_n281));
  nano32aa1n03x7               g186(.a(new_n218), .b(new_n281), .c(new_n237), .d(new_n260), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n236), .c(new_n125), .d(new_n179), .o1(new_n283));
  aob012aa1n02x5               g188(.a(new_n275), .b(\b[25] ), .c(\a[26] ), .out0(new_n284));
  oai012aa1n02x5               g189(.a(new_n284), .b(\b[25] ), .c(\a[26] ), .o1(new_n285));
  aoi012aa1d18x5               g190(.a(new_n285), .b(new_n268), .c(new_n281), .o1(new_n286));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  nand42aa1n03x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  nanb02aa1n06x5               g193(.a(new_n287), .b(new_n288), .out0(new_n289));
  xobna2aa1n03x5               g194(.a(new_n289), .b(new_n283), .c(new_n286), .out0(\s[27] ));
  oai012aa1n02x5               g195(.a(new_n288), .b(\b[27] ), .c(\a[28] ), .o1(new_n291));
  aoi012aa1n02x5               g196(.a(new_n291), .b(\a[28] ), .c(\b[27] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n281), .o1(new_n293));
  oaoi13aa1n02x5               g198(.a(new_n293), .b(new_n267), .c(new_n220), .d(new_n264), .o1(new_n294));
  nona32aa1n03x5               g199(.a(new_n283), .b(new_n287), .c(new_n285), .d(new_n294), .out0(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  nanp02aa1n03x5               g201(.a(new_n295), .b(new_n288), .o1(new_n297));
  aoi022aa1n02x7               g202(.a(new_n297), .b(new_n296), .c(new_n292), .d(new_n295), .o1(\s[28] ));
  inv040aa1n09x5               g203(.a(new_n286), .o1(new_n299));
  nor042aa1n03x5               g204(.a(new_n296), .b(new_n289), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n299), .c(new_n185), .d(new_n282), .o1(new_n301));
  inv000aa1n02x5               g206(.a(new_n300), .o1(new_n302));
  orn002aa1n02x5               g207(.a(\a[27] ), .b(\b[26] ), .o(new_n303));
  oao003aa1n03x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n303), .carry(new_n304));
  aoai13aa1n02x7               g209(.a(new_n304), .b(new_n302), .c(new_n283), .d(new_n286), .o1(new_n305));
  xorc02aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n304), .b(new_n306), .out0(new_n307));
  aoi022aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n301), .d(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g213(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g214(.a(new_n306), .b(new_n289), .c(new_n296), .out0(new_n310));
  aoai13aa1n06x5               g215(.a(new_n310), .b(new_n299), .c(new_n185), .d(new_n282), .o1(new_n311));
  inv000aa1n02x5               g216(.a(new_n310), .o1(new_n312));
  oaoi03aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .o1(new_n313));
  inv000aa1n03x5               g218(.a(new_n313), .o1(new_n314));
  aoai13aa1n02x7               g219(.a(new_n314), .b(new_n312), .c(new_n283), .d(new_n286), .o1(new_n315));
  xorc02aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n304), .b(\a[29] ), .c(\b[28] ), .o1(new_n317));
  oabi12aa1n02x5               g222(.a(new_n316), .b(\a[29] ), .c(\b[28] ), .out0(new_n318));
  norp02aa1n02x5               g223(.a(new_n317), .b(new_n318), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n315), .b(new_n316), .c(new_n311), .d(new_n319), .o1(\s[30] ));
  nano22aa1n06x5               g225(.a(new_n302), .b(new_n306), .c(new_n316), .out0(new_n321));
  aoai13aa1n06x5               g226(.a(new_n321), .b(new_n299), .c(new_n185), .d(new_n282), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[31] ), .b(\b[30] ), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n314), .carry(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(new_n325));
  inv000aa1d42x5               g230(.a(new_n321), .o1(new_n326));
  aoai13aa1n02x7               g231(.a(new_n324), .b(new_n326), .c(new_n283), .d(new_n286), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n323), .c(new_n322), .d(new_n325), .o1(\s[31] ));
  oai012aa1n02x5               g233(.a(new_n101), .b(new_n106), .c(new_n105), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n329), .b(new_n99), .c(new_n102), .out0(\s[3] ));
  oaoi03aa1n02x5               g235(.a(\a[3] ), .b(\b[2] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g237(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanp02aa1n02x5               g238(.a(\b[4] ), .b(\a[5] ), .o1(new_n334));
  oai012aa1n02x5               g239(.a(new_n334), .b(new_n108), .c(new_n110), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[5] ), .c(new_n117), .out0(\s[6] ));
  nanb02aa1n02x5               g241(.a(new_n113), .b(new_n114), .out0(new_n337));
  oaoi13aa1n03x5               g242(.a(new_n337), .b(new_n119), .c(new_n335), .d(new_n109), .o1(new_n338));
  oai112aa1n02x5               g243(.a(new_n119), .b(new_n337), .c(new_n335), .d(new_n109), .o1(new_n339));
  norb02aa1n02x5               g244(.a(new_n339), .b(new_n338), .out0(\s[7] ));
  norp02aa1n02x5               g245(.a(new_n338), .b(new_n113), .o1(new_n341));
  xnrb03aa1n03x5               g246(.a(new_n341), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g247(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


