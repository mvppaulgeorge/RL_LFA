// Benchmark "adder" written by ABC on Wed Jul 17 15:12:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n347, new_n350, new_n352, new_n353, new_n355, new_n356,
    new_n357, new_n358;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d30x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  norp02aa1n04x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n04x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  aoi012aa1d18x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nand02aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n12x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n104), .b(new_n107), .c(new_n106), .d(new_n105), .out0(new_n108));
  oa0012aa1n03x5               g013(.a(new_n104), .b(new_n105), .c(new_n106), .o(new_n109));
  inv000aa1n02x5               g014(.a(new_n109), .o1(new_n110));
  oai012aa1n06x5               g015(.a(new_n110), .b(new_n108), .c(new_n103), .o1(new_n111));
  nand02aa1d10x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  inv020aa1n04x5               g018(.a(new_n113), .o1(new_n114));
  oai112aa1n06x5               g019(.a(new_n114), .b(new_n112), .c(\b[6] ), .d(\a[7] ), .o1(new_n115));
  nor042aa1n06x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nand42aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nanb02aa1n09x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  nand22aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nand02aa1n06x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nor042aa1n06x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nanb03aa1n03x5               g026(.a(new_n121), .b(new_n119), .c(new_n120), .out0(new_n122));
  nor043aa1n03x5               g027(.a(new_n115), .b(new_n122), .c(new_n118), .o1(new_n123));
  inv040aa1n03x5               g028(.a(new_n115), .o1(new_n124));
  tech160nm_fiao0012aa1n05x5   g029(.a(new_n121), .b(new_n116), .c(new_n119), .o(new_n125));
  nor042aa1n09x5               g030(.a(\b[6] ), .b(\a[7] ), .o1(new_n126));
  nano23aa1n06x5               g031(.a(new_n126), .b(new_n113), .c(new_n120), .d(new_n112), .out0(new_n127));
  nanp02aa1n02x5               g032(.a(new_n127), .b(new_n125), .o1(new_n128));
  oaib12aa1n06x5               g033(.a(new_n128), .b(new_n124), .c(new_n112), .out0(new_n129));
  xorc02aa1n02x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n129), .c(new_n111), .d(new_n123), .o1(new_n131));
  nor002aa1d32x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nand42aa1d28x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norb02aa1n03x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n131), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g040(.a(new_n132), .o1(new_n136));
  inv000aa1n02x5               g041(.a(new_n133), .o1(new_n137));
  nor042aa1d18x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand02aa1d04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  inv000aa1n02x5               g045(.a(new_n140), .o1(new_n141));
  aoi113aa1n02x5               g046(.a(new_n141), .b(new_n137), .c(new_n131), .d(new_n136), .e(new_n99), .o1(new_n142));
  inv000aa1n02x5               g047(.a(new_n103), .o1(new_n143));
  nano23aa1n03x5               g048(.a(new_n106), .b(new_n105), .c(new_n107), .d(new_n104), .out0(new_n144));
  aoai13aa1n06x5               g049(.a(new_n123), .b(new_n109), .c(new_n143), .d(new_n144), .o1(new_n145));
  aoi022aa1n06x5               g050(.a(new_n127), .b(new_n125), .c(new_n112), .d(new_n115), .o1(new_n146));
  and002aa1n02x5               g051(.a(\b[8] ), .b(\a[9] ), .o(new_n147));
  aoai13aa1n03x5               g052(.a(new_n99), .b(new_n147), .c(new_n145), .d(new_n146), .o1(new_n148));
  aoai13aa1n12x5               g053(.a(new_n133), .b(new_n132), .c(new_n97), .d(new_n98), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoi112aa1n02x5               g055(.a(new_n150), .b(new_n140), .c(new_n148), .d(new_n134), .o1(new_n151));
  norp02aa1n02x5               g056(.a(new_n151), .b(new_n142), .o1(\s[11] ));
  inv000aa1n02x5               g057(.a(new_n138), .o1(new_n153));
  nor042aa1n09x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  nand42aa1d28x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  norb02aa1n12x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  nano22aa1n03x5               g062(.a(new_n142), .b(new_n153), .c(new_n157), .out0(new_n158));
  aoai13aa1n03x5               g063(.a(new_n140), .b(new_n150), .c(new_n148), .d(new_n134), .o1(new_n159));
  aoi012aa1n03x5               g064(.a(new_n157), .b(new_n159), .c(new_n153), .o1(new_n160));
  nor002aa1n02x5               g065(.a(new_n160), .b(new_n158), .o1(\s[12] ));
  oai112aa1n02x5               g066(.a(new_n153), .b(new_n139), .c(new_n98), .d(new_n97), .o1(new_n162));
  nano32aa1n02x4               g067(.a(new_n162), .b(new_n156), .c(new_n134), .d(new_n99), .out0(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n129), .c(new_n111), .d(new_n123), .o1(new_n164));
  tech160nm_fioai012aa1n03p5x5 g069(.a(new_n155), .b(new_n154), .c(new_n138), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n155), .b(new_n139), .c(new_n138), .d(new_n154), .out0(new_n166));
  oai012aa1d24x5               g071(.a(new_n165), .b(new_n166), .c(new_n149), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  nor002aa1d32x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nand02aa1n04x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n164), .c(new_n168), .out0(\s[13] ));
  inv000aa1d42x5               g077(.a(new_n169), .o1(new_n173));
  nanp02aa1n02x5               g078(.a(new_n144), .b(new_n143), .o1(new_n174));
  nona22aa1n02x4               g079(.a(new_n124), .b(new_n122), .c(new_n118), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n146), .b(new_n175), .c(new_n174), .d(new_n110), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n171), .b(new_n167), .c(new_n176), .d(new_n163), .o1(new_n177));
  nor002aa1d32x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nand22aa1n09x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  xobna2aa1n03x5               g085(.a(new_n180), .b(new_n177), .c(new_n173), .out0(\s[14] ));
  oai012aa1n18x5               g086(.a(new_n179), .b(new_n178), .c(new_n169), .o1(new_n182));
  nona23aa1n03x5               g087(.a(new_n179), .b(new_n170), .c(new_n169), .d(new_n178), .out0(new_n183));
  aoai13aa1n03x5               g088(.a(new_n182), .b(new_n183), .c(new_n164), .d(new_n168), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  nand02aa1n06x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  nor042aa1n04x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  nand02aa1d04x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  norb02aa1n02x5               g094(.a(new_n189), .b(new_n188), .out0(new_n190));
  aoi112aa1n03x4               g095(.a(new_n186), .b(new_n190), .c(new_n184), .d(new_n187), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n186), .o1(new_n192));
  aoi112aa1n02x7               g097(.a(new_n137), .b(new_n132), .c(new_n97), .d(new_n98), .o1(new_n193));
  nanb03aa1n02x5               g098(.a(new_n162), .b(new_n193), .c(new_n156), .out0(new_n194));
  aoai13aa1n03x5               g099(.a(new_n168), .b(new_n194), .c(new_n145), .d(new_n146), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n182), .o1(new_n196));
  nano23aa1n03x7               g101(.a(new_n169), .b(new_n178), .c(new_n179), .d(new_n170), .out0(new_n197));
  norb02aa1n02x5               g102(.a(new_n187), .b(new_n186), .out0(new_n198));
  aoai13aa1n03x5               g103(.a(new_n198), .b(new_n196), .c(new_n195), .d(new_n197), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n190), .o1(new_n200));
  tech160nm_fiaoi012aa1n03p5x5 g105(.a(new_n200), .b(new_n199), .c(new_n192), .o1(new_n201));
  nor042aa1n03x5               g106(.a(new_n201), .b(new_n191), .o1(\s[16] ));
  xorc02aa1n02x5               g107(.a(\a[17] ), .b(\b[16] ), .out0(new_n203));
  nona23aa1n03x5               g108(.a(new_n156), .b(new_n139), .c(new_n147), .d(new_n138), .out0(new_n204));
  nona23aa1d18x5               g109(.a(new_n189), .b(new_n187), .c(new_n186), .d(new_n188), .out0(new_n205));
  nano23aa1n03x7               g110(.a(new_n204), .b(new_n205), .c(new_n197), .d(new_n193), .out0(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n129), .c(new_n111), .d(new_n123), .o1(new_n207));
  nor002aa1n03x5               g112(.a(new_n205), .b(new_n183), .o1(new_n208));
  oai012aa1n02x7               g113(.a(new_n189), .b(new_n188), .c(new_n186), .o1(new_n209));
  tech160nm_fioai012aa1n04x5   g114(.a(new_n209), .b(new_n205), .c(new_n182), .o1(new_n210));
  aoi012aa1d24x5               g115(.a(new_n210), .b(new_n167), .c(new_n208), .o1(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n203), .b(new_n207), .c(new_n211), .out0(\s[17] ));
  orn002aa1n24x5               g117(.a(\a[17] ), .b(\b[16] ), .o(new_n213));
  nanp02aa1n03x5               g118(.a(new_n167), .b(new_n208), .o1(new_n214));
  inv000aa1n02x5               g119(.a(new_n210), .o1(new_n215));
  nanp02aa1n03x5               g120(.a(new_n214), .b(new_n215), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n203), .b(new_n216), .c(new_n176), .d(new_n206), .o1(new_n217));
  xnrc02aa1n12x5               g122(.a(\b[17] ), .b(\a[18] ), .out0(new_n218));
  xobna2aa1n03x5               g123(.a(new_n218), .b(new_n217), .c(new_n213), .out0(\s[18] ));
  nanp02aa1n02x5               g124(.a(\b[16] ), .b(\a[17] ), .o1(new_n220));
  nano22aa1n12x5               g125(.a(new_n218), .b(new_n213), .c(new_n220), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oaoi03aa1n12x5               g127(.a(\a[18] ), .b(\b[17] ), .c(new_n213), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n02x5               g129(.a(new_n224), .b(new_n222), .c(new_n207), .d(new_n211), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g131(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g132(.a(\b[18] ), .b(\a[19] ), .o1(new_n228));
  nand42aa1n08x5               g133(.a(\b[18] ), .b(\a[19] ), .o1(new_n229));
  nor002aa1n03x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  nand42aa1n06x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  nanb02aa1n02x5               g136(.a(new_n230), .b(new_n231), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoi112aa1n02x5               g138(.a(new_n228), .b(new_n233), .c(new_n225), .d(new_n229), .o1(new_n234));
  inv000aa1n02x5               g139(.a(new_n228), .o1(new_n235));
  nand02aa1n02x5               g140(.a(new_n163), .b(new_n208), .o1(new_n236));
  aoai13aa1n09x5               g141(.a(new_n211), .b(new_n236), .c(new_n145), .d(new_n146), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n229), .b(new_n228), .out0(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n223), .c(new_n237), .d(new_n221), .o1(new_n239));
  aoi012aa1n03x5               g144(.a(new_n232), .b(new_n239), .c(new_n235), .o1(new_n240));
  norp02aa1n03x5               g145(.a(new_n240), .b(new_n234), .o1(\s[20] ));
  nano23aa1d12x5               g146(.a(new_n228), .b(new_n230), .c(new_n231), .d(new_n229), .out0(new_n242));
  nand02aa1d06x5               g147(.a(new_n221), .b(new_n242), .o1(new_n243));
  oaoi03aa1n06x5               g148(.a(\a[20] ), .b(\b[19] ), .c(new_n235), .o1(new_n244));
  aoi012aa1d24x5               g149(.a(new_n244), .b(new_n242), .c(new_n223), .o1(new_n245));
  aoai13aa1n02x7               g150(.a(new_n245), .b(new_n243), .c(new_n207), .d(new_n211), .o1(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n06x5               g152(.a(\b[20] ), .b(\a[21] ), .o1(new_n248));
  nand02aa1n06x5               g153(.a(\b[20] ), .b(\a[21] ), .o1(new_n249));
  nor022aa1n08x5               g154(.a(\b[21] ), .b(\a[22] ), .o1(new_n250));
  nand42aa1n03x5               g155(.a(\b[21] ), .b(\a[22] ), .o1(new_n251));
  norb02aa1n02x5               g156(.a(new_n251), .b(new_n250), .out0(new_n252));
  aoi112aa1n02x5               g157(.a(new_n248), .b(new_n252), .c(new_n246), .d(new_n249), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n248), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n243), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n245), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n249), .b(new_n248), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n256), .c(new_n237), .d(new_n255), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n252), .o1(new_n259));
  aoi012aa1n03x5               g164(.a(new_n259), .b(new_n258), .c(new_n254), .o1(new_n260));
  norp02aa1n03x5               g165(.a(new_n260), .b(new_n253), .o1(\s[22] ));
  nona23aa1n09x5               g166(.a(new_n251), .b(new_n249), .c(new_n248), .d(new_n250), .out0(new_n262));
  nano22aa1n09x5               g167(.a(new_n262), .b(new_n221), .c(new_n242), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  oaoi03aa1n09x5               g169(.a(\a[22] ), .b(\b[21] ), .c(new_n254), .o1(new_n265));
  oab012aa1n06x5               g170(.a(new_n265), .b(new_n245), .c(new_n262), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n264), .c(new_n207), .d(new_n211), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n16x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  nand02aa1n02x5               g174(.a(\b[22] ), .b(\a[23] ), .o1(new_n270));
  nor002aa1n03x5               g175(.a(\b[23] ), .b(\a[24] ), .o1(new_n271));
  nanp02aa1n04x5               g176(.a(\b[23] ), .b(\a[24] ), .o1(new_n272));
  nanb02aa1n02x5               g177(.a(new_n271), .b(new_n272), .out0(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  aoi112aa1n02x5               g179(.a(new_n269), .b(new_n274), .c(new_n267), .d(new_n270), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n269), .o1(new_n276));
  inv040aa1n03x5               g181(.a(new_n266), .o1(new_n277));
  norb02aa1n02x5               g182(.a(new_n270), .b(new_n269), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n237), .d(new_n263), .o1(new_n279));
  tech160nm_fiaoi012aa1n05x5   g184(.a(new_n273), .b(new_n279), .c(new_n276), .o1(new_n280));
  norp02aa1n03x5               g185(.a(new_n280), .b(new_n275), .o1(\s[24] ));
  nona23aa1n03x5               g186(.a(new_n272), .b(new_n270), .c(new_n269), .d(new_n271), .out0(new_n282));
  nor042aa1n02x5               g187(.a(new_n282), .b(new_n262), .o1(new_n283));
  norb02aa1n02x5               g188(.a(new_n283), .b(new_n243), .out0(new_n284));
  inv000aa1n02x5               g189(.a(new_n284), .o1(new_n285));
  nona22aa1n02x4               g190(.a(new_n272), .b(new_n271), .c(new_n269), .out0(new_n286));
  aboi22aa1n09x5               g191(.a(new_n282), .b(new_n265), .c(new_n272), .d(new_n286), .out0(new_n287));
  oaib12aa1n18x5               g192(.a(new_n287), .b(new_n245), .c(new_n283), .out0(new_n288));
  inv020aa1n04x5               g193(.a(new_n288), .o1(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n285), .c(new_n207), .d(new_n211), .o1(new_n290));
  xorb03aa1n02x5               g195(.a(new_n290), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor002aa1n02x5               g196(.a(\b[24] ), .b(\a[25] ), .o1(new_n292));
  nanp02aa1n02x5               g197(.a(\b[24] ), .b(\a[25] ), .o1(new_n293));
  tech160nm_fixorc02aa1n05x5   g198(.a(\a[26] ), .b(\b[25] ), .out0(new_n294));
  aoi112aa1n02x5               g199(.a(new_n292), .b(new_n294), .c(new_n290), .d(new_n293), .o1(new_n295));
  inv000aa1n02x5               g200(.a(new_n292), .o1(new_n296));
  norb02aa1n02x5               g201(.a(new_n293), .b(new_n292), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n288), .c(new_n237), .d(new_n284), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n294), .o1(new_n299));
  aoi012aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n296), .o1(new_n300));
  nor002aa1n02x5               g205(.a(new_n300), .b(new_n295), .o1(\s[26] ));
  nano22aa1n12x5               g206(.a(new_n299), .b(new_n296), .c(new_n293), .out0(new_n302));
  nano22aa1n02x5               g207(.a(new_n243), .b(new_n302), .c(new_n283), .out0(new_n303));
  aoai13aa1n04x5               g208(.a(new_n303), .b(new_n216), .c(new_n176), .d(new_n206), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[26] ), .b(\b[25] ), .c(new_n296), .carry(new_n305));
  aobi12aa1n12x5               g210(.a(new_n305), .b(new_n288), .c(new_n302), .out0(new_n306));
  norp02aa1n02x5               g211(.a(\b[26] ), .b(\a[27] ), .o1(new_n307));
  nanp02aa1n02x5               g212(.a(\b[26] ), .b(\a[27] ), .o1(new_n308));
  norb02aa1n02x5               g213(.a(new_n308), .b(new_n307), .out0(new_n309));
  xnbna2aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n306), .out0(\s[27] ));
  inv000aa1n06x5               g215(.a(new_n307), .o1(new_n311));
  aobi12aa1n02x7               g216(.a(new_n309), .b(new_n304), .c(new_n306), .out0(new_n312));
  xnrc02aa1n02x5               g217(.a(\b[27] ), .b(\a[28] ), .out0(new_n313));
  nano22aa1n03x5               g218(.a(new_n312), .b(new_n311), .c(new_n313), .out0(new_n314));
  aoai13aa1n03x5               g219(.a(new_n283), .b(new_n244), .c(new_n223), .d(new_n242), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n302), .o1(new_n316));
  aoai13aa1n04x5               g221(.a(new_n305), .b(new_n316), .c(new_n315), .d(new_n287), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n309), .b(new_n317), .c(new_n237), .d(new_n303), .o1(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n313), .b(new_n318), .c(new_n311), .o1(new_n319));
  norp02aa1n03x5               g224(.a(new_n319), .b(new_n314), .o1(\s[28] ));
  xnrc02aa1n02x5               g225(.a(\b[28] ), .b(\a[29] ), .out0(new_n321));
  nano22aa1n02x4               g226(.a(new_n313), .b(new_n311), .c(new_n308), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n317), .c(new_n237), .d(new_n303), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[28] ), .b(\b[27] ), .c(new_n311), .carry(new_n324));
  tech160nm_fiaoi012aa1n02p5x5 g229(.a(new_n321), .b(new_n323), .c(new_n324), .o1(new_n325));
  aobi12aa1n02x7               g230(.a(new_n322), .b(new_n304), .c(new_n306), .out0(new_n326));
  nano22aa1n03x5               g231(.a(new_n326), .b(new_n321), .c(new_n324), .out0(new_n327));
  norp02aa1n03x5               g232(.a(new_n325), .b(new_n327), .o1(\s[29] ));
  xorb03aa1n02x5               g233(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  oao003aa1n02x5               g234(.a(\a[29] ), .b(\b[28] ), .c(new_n324), .carry(new_n330));
  nano23aa1n02x4               g235(.a(new_n321), .b(new_n313), .c(new_n308), .d(new_n311), .out0(new_n331));
  aoai13aa1n03x5               g236(.a(new_n331), .b(new_n317), .c(new_n237), .d(new_n303), .o1(new_n332));
  xnrc02aa1n02x5               g237(.a(\b[29] ), .b(\a[30] ), .out0(new_n333));
  tech160nm_fiaoi012aa1n02p5x5 g238(.a(new_n333), .b(new_n332), .c(new_n330), .o1(new_n334));
  aobi12aa1n02x7               g239(.a(new_n331), .b(new_n304), .c(new_n306), .out0(new_n335));
  nano22aa1n03x5               g240(.a(new_n335), .b(new_n330), .c(new_n333), .out0(new_n336));
  norp02aa1n03x5               g241(.a(new_n334), .b(new_n336), .o1(\s[30] ));
  norb03aa1n02x5               g242(.a(new_n322), .b(new_n321), .c(new_n333), .out0(new_n338));
  aobi12aa1n06x5               g243(.a(new_n338), .b(new_n304), .c(new_n306), .out0(new_n339));
  oao003aa1n02x5               g244(.a(\a[30] ), .b(\b[29] ), .c(new_n330), .carry(new_n340));
  xnrc02aa1n02x5               g245(.a(\b[30] ), .b(\a[31] ), .out0(new_n341));
  nano22aa1n02x4               g246(.a(new_n339), .b(new_n340), .c(new_n341), .out0(new_n342));
  aoai13aa1n03x5               g247(.a(new_n338), .b(new_n317), .c(new_n237), .d(new_n303), .o1(new_n343));
  tech160nm_fiaoi012aa1n02p5x5 g248(.a(new_n341), .b(new_n343), .c(new_n340), .o1(new_n344));
  norp02aa1n03x5               g249(.a(new_n344), .b(new_n342), .o1(\s[31] ));
  xnrb03aa1n02x5               g250(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g251(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n347));
  xorb03aa1n02x5               g252(.a(new_n347), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g253(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fiaoi012aa1n05x5   g254(.a(new_n116), .b(new_n111), .c(new_n117), .o1(new_n350));
  xnrb03aa1n02x5               g255(.a(new_n350), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g256(.a(new_n126), .o1(new_n352));
  oaib12aa1n03x5               g257(.a(new_n119), .b(new_n121), .c(new_n350), .out0(new_n353));
  xnbna2aa1n03x5               g258(.a(new_n353), .b(new_n352), .c(new_n120), .out0(\s[7] ));
  nanb02aa1n02x5               g259(.a(new_n113), .b(new_n112), .out0(new_n355));
  nanb02aa1n02x5               g260(.a(new_n126), .b(new_n120), .out0(new_n356));
  oaoi13aa1n02x7               g261(.a(new_n355), .b(new_n352), .c(new_n353), .d(new_n356), .o1(new_n357));
  oai112aa1n03x5               g262(.a(new_n355), .b(new_n352), .c(new_n353), .d(new_n356), .o1(new_n358));
  norb02aa1n02x7               g263(.a(new_n358), .b(new_n357), .out0(\s[8] ));
  xnbna2aa1n03x5               g264(.a(new_n130), .b(new_n145), .c(new_n146), .out0(\s[9] ));
endmodule


