// Benchmark "adder" written by ABC on Thu Jul 18 01:12:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n336, new_n338, new_n340,
    new_n341, new_n342, new_n343, new_n346;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1d18x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n08x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n09x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  norp02aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanb02aa1n03x5               g009(.a(new_n103), .b(new_n104), .out0(new_n105));
  inv040aa1d32x5               g010(.a(\a[3] ), .o1(new_n106));
  inv040aa1d28x5               g011(.a(\b[2] ), .o1(new_n107));
  nand02aa1d16x5               g012(.a(new_n107), .b(new_n106), .o1(new_n108));
  nand02aa1n04x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(new_n108), .b(new_n109), .o1(new_n110));
  nor043aa1n02x5               g015(.a(new_n102), .b(new_n105), .c(new_n110), .o1(new_n111));
  oaoi03aa1n06x5               g016(.a(\a[4] ), .b(\b[3] ), .c(new_n108), .o1(new_n112));
  nor042aa1n06x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand02aa1d28x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor042aa1d18x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n03x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nona23aa1n03x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nor042aa1n04x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1d28x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nor042aa1n04x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nand42aa1n06x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nona23aa1n03x5               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  nor042aa1n02x5               g027(.a(new_n122), .b(new_n117), .o1(new_n123));
  tech160nm_fioai012aa1n05x5   g028(.a(new_n123), .b(new_n111), .c(new_n112), .o1(new_n124));
  nano23aa1d15x5               g029(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n125));
  inv040aa1n06x5               g030(.a(new_n113), .o1(new_n126));
  aob012aa1d24x5               g031(.a(new_n126), .b(new_n115), .c(new_n114), .out0(new_n127));
  oai022aa1n06x5               g032(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n128));
  aoi022aa1d24x5               g033(.a(new_n125), .b(new_n127), .c(new_n119), .d(new_n128), .o1(new_n129));
  nanp02aa1n04x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  norb02aa1d21x5               g035(.a(new_n130), .b(new_n97), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  aoai13aa1n02x5               g037(.a(new_n98), .b(new_n132), .c(new_n124), .d(new_n129), .o1(new_n133));
  xorb03aa1n02x5               g038(.a(new_n133), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  inv000aa1d42x5               g039(.a(new_n99), .o1(new_n135));
  aob012aa1n03x5               g040(.a(new_n135), .b(new_n100), .c(new_n101), .out0(new_n136));
  norb02aa1n06x5               g041(.a(new_n104), .b(new_n103), .out0(new_n137));
  nor042aa1n02x5               g042(.a(\b[2] ), .b(\a[3] ), .o1(new_n138));
  norb02aa1n03x5               g043(.a(new_n109), .b(new_n138), .out0(new_n139));
  nand23aa1n06x5               g044(.a(new_n136), .b(new_n137), .c(new_n139), .o1(new_n140));
  inv030aa1n02x5               g045(.a(new_n112), .o1(new_n141));
  nano23aa1n03x7               g046(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n142));
  nand02aa1d04x5               g047(.a(new_n125), .b(new_n142), .o1(new_n143));
  aoai13aa1n12x5               g048(.a(new_n129), .b(new_n143), .c(new_n140), .d(new_n141), .o1(new_n144));
  nor002aa1n06x5               g049(.a(\b[9] ), .b(\a[10] ), .o1(new_n145));
  nand02aa1n06x5               g050(.a(\b[9] ), .b(\a[10] ), .o1(new_n146));
  norb02aa1n09x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  aoai13aa1n06x5               g052(.a(new_n147), .b(new_n97), .c(new_n144), .d(new_n130), .o1(new_n148));
  oai012aa1n06x5               g053(.a(new_n148), .b(\b[9] ), .c(\a[10] ), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n12x5               g055(.a(\b[10] ), .b(\a[11] ), .o1(new_n151));
  nand02aa1d06x5               g056(.a(\b[10] ), .b(\a[11] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  nor002aa1n16x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  nand02aa1n08x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n154), .b(new_n155), .out0(new_n156));
  aoai13aa1n03x5               g061(.a(new_n156), .b(new_n151), .c(new_n149), .d(new_n153), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n153), .b(new_n145), .c(new_n133), .d(new_n146), .o1(new_n158));
  nona22aa1n02x4               g063(.a(new_n158), .b(new_n156), .c(new_n151), .out0(new_n159));
  nanp02aa1n02x5               g064(.a(new_n157), .b(new_n159), .o1(\s[12] ));
  nona23aa1d18x5               g065(.a(new_n155), .b(new_n152), .c(new_n151), .d(new_n154), .out0(new_n161));
  nano22aa1d15x5               g066(.a(new_n161), .b(new_n131), .c(new_n147), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nano23aa1n09x5               g068(.a(new_n151), .b(new_n154), .c(new_n155), .d(new_n152), .out0(new_n164));
  aoi012aa1n09x5               g069(.a(new_n145), .b(new_n97), .c(new_n146), .o1(new_n165));
  inv040aa1n03x5               g070(.a(new_n165), .o1(new_n166));
  tech160nm_fioai012aa1n03p5x5 g071(.a(new_n155), .b(new_n154), .c(new_n151), .o1(new_n167));
  aobi12aa1n02x5               g072(.a(new_n167), .b(new_n164), .c(new_n166), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n163), .c(new_n124), .d(new_n129), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n06x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nand22aa1n03x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n173));
  xnrb03aa1n02x5               g078(.a(new_n173), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  oai012aa1n06x5               g079(.a(new_n167), .b(new_n161), .c(new_n165), .o1(new_n175));
  nor042aa1n06x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  nand02aa1n03x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nano23aa1n06x5               g082(.a(new_n171), .b(new_n176), .c(new_n177), .d(new_n172), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n175), .c(new_n144), .d(new_n162), .o1(new_n179));
  aoi012aa1n02x7               g084(.a(new_n176), .b(new_n171), .c(new_n177), .o1(new_n180));
  nor002aa1n16x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  nand02aa1n04x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n182), .b(new_n181), .out0(new_n183));
  xnbna2aa1n03x5               g088(.a(new_n183), .b(new_n179), .c(new_n180), .out0(\s[15] ));
  nanp02aa1n03x5               g089(.a(new_n179), .b(new_n180), .o1(new_n185));
  nor022aa1n16x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nanp02aa1n04x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nanb02aa1n02x5               g092(.a(new_n186), .b(new_n187), .out0(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n181), .c(new_n185), .d(new_n183), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n185), .b(new_n183), .o1(new_n190));
  nona22aa1n02x4               g095(.a(new_n190), .b(new_n188), .c(new_n181), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(new_n191), .b(new_n189), .o1(\s[16] ));
  nona23aa1n03x5               g097(.a(new_n177), .b(new_n172), .c(new_n171), .d(new_n176), .out0(new_n193));
  nona23aa1d18x5               g098(.a(new_n187), .b(new_n182), .c(new_n181), .d(new_n186), .out0(new_n194));
  nor042aa1n02x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  nand22aa1n03x5               g100(.a(new_n162), .b(new_n195), .o1(new_n196));
  oai012aa1n02x5               g101(.a(new_n187), .b(new_n186), .c(new_n181), .o1(new_n197));
  oaih12aa1n02x5               g102(.a(new_n197), .b(new_n194), .c(new_n180), .o1(new_n198));
  aoi012aa1n06x5               g103(.a(new_n198), .b(new_n175), .c(new_n195), .o1(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n196), .c(new_n124), .d(new_n129), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g106(.a(\a[18] ), .o1(new_n202));
  inv000aa1d42x5               g107(.a(\a[17] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(\b[16] ), .o1(new_n204));
  oaoi03aa1n03x5               g109(.a(new_n203), .b(new_n204), .c(new_n200), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[17] ), .c(new_n202), .out0(\s[18] ));
  nanb02aa1n06x5               g111(.a(new_n194), .b(new_n178), .out0(new_n207));
  nano32aa1n03x7               g112(.a(new_n207), .b(new_n164), .c(new_n147), .d(new_n131), .out0(new_n208));
  oabi12aa1n06x5               g113(.a(new_n198), .b(new_n168), .c(new_n207), .out0(new_n209));
  xroi22aa1d06x4               g114(.a(new_n203), .b(\b[16] ), .c(new_n202), .d(\b[17] ), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n209), .c(new_n144), .d(new_n208), .o1(new_n211));
  nor042aa1n02x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  aoi112aa1n09x5               g117(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n213));
  norp02aa1n02x5               g118(.a(new_n213), .b(new_n212), .o1(new_n214));
  nor042aa1n04x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand42aa1n08x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n12x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n211), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n03x5               g124(.a(new_n211), .b(new_n214), .o1(new_n220));
  nor002aa1n10x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand42aa1d28x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1d21x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n04x5               g129(.a(new_n224), .b(new_n215), .c(new_n220), .d(new_n216), .o1(new_n225));
  inv000aa1n02x5               g130(.a(new_n214), .o1(new_n226));
  aoai13aa1n02x5               g131(.a(new_n217), .b(new_n226), .c(new_n200), .d(new_n210), .o1(new_n227));
  nona22aa1n02x4               g132(.a(new_n227), .b(new_n224), .c(new_n215), .out0(new_n228));
  nanp02aa1n03x5               g133(.a(new_n225), .b(new_n228), .o1(\s[20] ));
  nanp02aa1n06x5               g134(.a(new_n144), .b(new_n208), .o1(new_n230));
  nano23aa1n02x5               g135(.a(new_n215), .b(new_n221), .c(new_n222), .d(new_n216), .out0(new_n231));
  nanp02aa1n02x5               g136(.a(new_n210), .b(new_n231), .o1(new_n232));
  oai112aa1n06x5               g137(.a(new_n217), .b(new_n223), .c(new_n213), .d(new_n212), .o1(new_n233));
  oai012aa1n06x5               g138(.a(new_n222), .b(new_n221), .c(new_n215), .o1(new_n234));
  nanp02aa1n12x5               g139(.a(new_n233), .b(new_n234), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n232), .c(new_n230), .d(new_n199), .o1(new_n237));
  xorb03aa1n02x5               g142(.a(new_n237), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n04x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[20] ), .b(\a[21] ), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  tech160nm_fixnrc02aa1n04x5   g146(.a(\b[21] ), .b(\a[22] ), .out0(new_n242));
  aoai13aa1n02x7               g147(.a(new_n242), .b(new_n239), .c(new_n237), .d(new_n241), .o1(new_n243));
  tech160nm_finand02aa1n03p5x5 g148(.a(new_n237), .b(new_n241), .o1(new_n244));
  nona22aa1n02x4               g149(.a(new_n244), .b(new_n242), .c(new_n239), .out0(new_n245));
  nanp02aa1n03x5               g150(.a(new_n245), .b(new_n243), .o1(\s[22] ));
  nor042aa1n06x5               g151(.a(new_n242), .b(new_n240), .o1(new_n247));
  nand23aa1n03x5               g152(.a(new_n210), .b(new_n247), .c(new_n231), .o1(new_n248));
  norp02aa1n02x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[21] ), .b(\a[22] ), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n249), .b(new_n239), .c(new_n250), .o1(new_n251));
  aobi12aa1n06x5               g156(.a(new_n251), .b(new_n235), .c(new_n247), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n248), .c(new_n230), .d(new_n199), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n04x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  nand22aa1n04x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  nanb02aa1n12x5               g161(.a(new_n255), .b(new_n256), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  nor002aa1d24x5               g163(.a(\b[23] ), .b(\a[24] ), .o1(new_n259));
  nanp02aa1n04x5               g164(.a(\b[23] ), .b(\a[24] ), .o1(new_n260));
  nanb02aa1n02x5               g165(.a(new_n259), .b(new_n260), .out0(new_n261));
  aoai13aa1n02x7               g166(.a(new_n261), .b(new_n255), .c(new_n253), .d(new_n258), .o1(new_n262));
  tech160nm_finand02aa1n03p5x5 g167(.a(new_n253), .b(new_n258), .o1(new_n263));
  nona22aa1n03x5               g168(.a(new_n263), .b(new_n261), .c(new_n255), .out0(new_n264));
  nanp02aa1n03x5               g169(.a(new_n264), .b(new_n262), .o1(\s[24] ));
  nona23aa1n09x5               g170(.a(new_n260), .b(new_n256), .c(new_n255), .d(new_n259), .out0(new_n266));
  inv000aa1n02x5               g171(.a(new_n266), .o1(new_n267));
  nano22aa1n02x4               g172(.a(new_n232), .b(new_n247), .c(new_n267), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n209), .c(new_n144), .d(new_n208), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n247), .o1(new_n270));
  aoi112aa1n03x5               g175(.a(new_n270), .b(new_n266), .c(new_n233), .d(new_n234), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n259), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(new_n255), .b(new_n260), .o1(new_n273));
  oai112aa1n02x5               g178(.a(new_n273), .b(new_n272), .c(new_n266), .d(new_n251), .o1(new_n274));
  nona22aa1n03x5               g179(.a(new_n269), .b(new_n271), .c(new_n274), .out0(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  xnrc02aa1n12x5               g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  aoai13aa1n02x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  nona32aa1n09x5               g185(.a(new_n235), .b(new_n266), .c(new_n242), .d(new_n240), .out0(new_n281));
  norp03aa1n02x5               g186(.a(new_n251), .b(new_n257), .c(new_n261), .o1(new_n282));
  nano22aa1n02x4               g187(.a(new_n282), .b(new_n272), .c(new_n273), .out0(new_n283));
  nanp02aa1n02x5               g188(.a(new_n281), .b(new_n283), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n278), .b(new_n284), .c(new_n200), .d(new_n268), .o1(new_n285));
  nona22aa1n02x4               g190(.a(new_n285), .b(new_n279), .c(new_n277), .out0(new_n286));
  nanp02aa1n02x5               g191(.a(new_n280), .b(new_n286), .o1(\s[26] ));
  norb02aa1n09x5               g192(.a(new_n278), .b(new_n279), .out0(new_n288));
  nano22aa1n03x7               g193(.a(new_n248), .b(new_n267), .c(new_n288), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n209), .c(new_n144), .d(new_n208), .o1(new_n290));
  inv000aa1d42x5               g195(.a(\a[26] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\b[25] ), .o1(new_n292));
  oao003aa1n02x5               g197(.a(new_n291), .b(new_n292), .c(new_n277), .carry(new_n293));
  oaoi13aa1n09x5               g198(.a(new_n293), .b(new_n288), .c(new_n271), .d(new_n274), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  xnbna2aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n290), .out0(\s[27] ));
  nanp02aa1n03x5               g201(.a(new_n294), .b(new_n290), .o1(new_n297));
  norp02aa1n02x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  tech160nm_fixorc02aa1n03p5x5 g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n298), .c(new_n297), .d(new_n295), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n288), .o1(new_n302));
  inv000aa1n02x5               g207(.a(new_n293), .o1(new_n303));
  aoai13aa1n06x5               g208(.a(new_n303), .b(new_n302), .c(new_n281), .d(new_n283), .o1(new_n304));
  aoai13aa1n02x5               g209(.a(new_n295), .b(new_n304), .c(new_n200), .d(new_n289), .o1(new_n305));
  nona22aa1n03x5               g210(.a(new_n305), .b(new_n300), .c(new_n298), .out0(new_n306));
  nanp02aa1n03x5               g211(.a(new_n301), .b(new_n306), .o1(\s[28] ));
  and002aa1n02x5               g212(.a(new_n299), .b(new_n295), .o(new_n308));
  aoai13aa1n02x5               g213(.a(new_n308), .b(new_n304), .c(new_n200), .d(new_n289), .o1(new_n309));
  aoi112aa1n02x5               g214(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n310));
  oab012aa1n02x4               g215(.a(new_n310), .b(\a[28] ), .c(\b[27] ), .out0(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[28] ), .b(\a[29] ), .out0(new_n312));
  aoi012aa1n02x5               g217(.a(new_n312), .b(new_n309), .c(new_n311), .o1(new_n313));
  aobi12aa1n03x5               g218(.a(new_n308), .b(new_n294), .c(new_n290), .out0(new_n314));
  nano22aa1n03x7               g219(.a(new_n314), .b(new_n311), .c(new_n312), .out0(new_n315));
  nor002aa1n02x5               g220(.a(new_n313), .b(new_n315), .o1(\s[29] ));
  xorb03aa1n02x5               g221(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g222(.a(new_n312), .b(new_n295), .c(new_n299), .out0(new_n318));
  aoai13aa1n02x5               g223(.a(new_n318), .b(new_n304), .c(new_n200), .d(new_n289), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .carry(new_n320));
  xnrc02aa1n02x5               g225(.a(\b[29] ), .b(\a[30] ), .out0(new_n321));
  aoi012aa1n02x5               g226(.a(new_n321), .b(new_n319), .c(new_n320), .o1(new_n322));
  aobi12aa1n03x5               g227(.a(new_n318), .b(new_n294), .c(new_n290), .out0(new_n323));
  nano22aa1n03x7               g228(.a(new_n323), .b(new_n320), .c(new_n321), .out0(new_n324));
  nor002aa1n02x5               g229(.a(new_n322), .b(new_n324), .o1(\s[30] ));
  nano23aa1n02x4               g230(.a(new_n321), .b(new_n312), .c(new_n299), .d(new_n295), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n304), .c(new_n200), .d(new_n289), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n320), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  aoi012aa1n03x5               g234(.a(new_n329), .b(new_n327), .c(new_n328), .o1(new_n330));
  aobi12aa1n03x5               g235(.a(new_n326), .b(new_n294), .c(new_n290), .out0(new_n331));
  nano22aa1n03x7               g236(.a(new_n331), .b(new_n328), .c(new_n329), .out0(new_n332));
  norp02aa1n03x5               g237(.a(new_n330), .b(new_n332), .o1(\s[31] ));
  xnbna2aa1n03x5               g238(.a(new_n102), .b(new_n109), .c(new_n108), .out0(\s[3] ));
  orn002aa1n02x5               g239(.a(\a[4] ), .b(\b[3] ), .o(new_n335));
  aoi112aa1n02x5               g240(.a(new_n138), .b(new_n137), .c(new_n136), .d(new_n139), .o1(new_n336));
  oaoi13aa1n02x5               g241(.a(new_n336), .b(new_n335), .c(new_n111), .d(new_n112), .o1(\s[4] ));
  nanb02aa1n02x5               g242(.a(new_n115), .b(new_n116), .out0(new_n338));
  xobna2aa1n03x5               g243(.a(new_n338), .b(new_n140), .c(new_n141), .out0(\s[5] ));
  oabi12aa1n02x5               g244(.a(new_n338), .b(new_n111), .c(new_n112), .out0(new_n340));
  aoi012aa1n02x5               g245(.a(new_n115), .b(new_n126), .c(new_n114), .o1(new_n341));
  inv000aa1d42x5               g246(.a(new_n127), .o1(new_n342));
  aoai13aa1n02x5               g247(.a(new_n342), .b(new_n117), .c(new_n140), .d(new_n141), .o1(new_n343));
  aoi022aa1n02x5               g248(.a(new_n343), .b(new_n126), .c(new_n340), .d(new_n341), .o1(\s[6] ));
  xorb03aa1n02x5               g249(.a(new_n343), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g250(.a(new_n120), .b(new_n343), .c(new_n121), .o1(new_n346));
  xnrb03aa1n02x5               g251(.a(new_n346), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g252(.a(new_n144), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


