// Benchmark "adder" written by ABC on Thu Jul 18 06:25:34 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n338, new_n339, new_n340, new_n341, new_n343, new_n344, new_n345,
    new_n346, new_n348, new_n349, new_n351, new_n352, new_n353, new_n355,
    new_n356, new_n358, new_n359, new_n361, new_n362, new_n363;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv030aa1d32x5               g003(.a(\a[2] ), .o1(new_n99));
  inv040aa1d30x5               g004(.a(\b[1] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n12x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor022aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  tech160nm_fioai012aa1n03p5x5 g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oai012aa1n18x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  xnrc02aa1n03x5               g014(.a(\b[7] ), .b(\a[8] ), .out0(new_n110));
  norp02aa1n12x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n16x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanb02aa1n06x5               g017(.a(new_n111), .b(new_n112), .out0(new_n113));
  nand02aa1n06x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor002aa1d24x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nona23aa1n09x5               g022(.a(new_n114), .b(new_n117), .c(new_n116), .d(new_n115), .out0(new_n118));
  nor003aa1n12x5               g023(.a(new_n118), .b(new_n113), .c(new_n110), .o1(new_n119));
  nand42aa1n06x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nano22aa1n02x4               g025(.a(new_n111), .b(new_n120), .c(new_n112), .out0(new_n121));
  oai122aa1n02x5               g026(.a(new_n114), .b(new_n115), .c(new_n116), .d(\b[7] ), .e(\a[8] ), .o1(new_n122));
  norp02aa1n02x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  oai012aa1n02x5               g028(.a(new_n120), .b(new_n111), .c(new_n123), .o1(new_n124));
  oaib12aa1n06x5               g029(.a(new_n124), .b(new_n122), .c(new_n121), .out0(new_n125));
  nand42aa1n16x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1d21x5               g031(.a(new_n126), .b(new_n97), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n128));
  nor002aa1n10x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1n16x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  norp02aa1n02x5               g036(.a(new_n129), .b(new_n97), .o1(new_n132));
  nanp03aa1n02x5               g037(.a(new_n128), .b(new_n130), .c(new_n132), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n131), .c(new_n98), .d(new_n128), .o1(\s[10] ));
  nano23aa1n02x5               g039(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n126), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n136));
  oai012aa1n02x5               g041(.a(new_n130), .b(new_n129), .c(new_n97), .o1(new_n137));
  nor002aa1n10x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand42aa1n10x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n136), .c(new_n137), .out0(\s[11] ));
  inv040aa1n02x5               g046(.a(new_n138), .o1(new_n142));
  aob012aa1n02x5               g047(.a(new_n140), .b(new_n136), .c(new_n137), .out0(new_n143));
  nor042aa1n06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanp02aa1n12x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  nona23aa1n02x4               g051(.a(new_n143), .b(new_n145), .c(new_n144), .d(new_n138), .out0(new_n147));
  aoai13aa1n02x5               g052(.a(new_n147), .b(new_n146), .c(new_n143), .d(new_n142), .o1(\s[12] ));
  inv000aa1d42x5               g053(.a(new_n127), .o1(new_n149));
  nano32aa1n03x7               g054(.a(new_n149), .b(new_n146), .c(new_n131), .d(new_n140), .out0(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n151));
  nano22aa1n03x7               g056(.a(new_n144), .b(new_n139), .c(new_n145), .out0(new_n152));
  oai112aa1n06x5               g057(.a(new_n142), .b(new_n130), .c(new_n129), .d(new_n97), .o1(new_n153));
  oai012aa1n12x5               g058(.a(new_n145), .b(new_n144), .c(new_n138), .o1(new_n154));
  oaib12aa1n18x5               g059(.a(new_n154), .b(new_n153), .c(new_n152), .out0(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nand02aa1d04x5               g061(.a(new_n151), .b(new_n156), .o1(new_n157));
  nor042aa1d18x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand42aa1n04x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n159), .b(new_n158), .out0(new_n160));
  oaib12aa1n02x5               g065(.a(new_n154), .b(new_n158), .c(new_n159), .out0(new_n161));
  aoib12aa1n02x5               g066(.a(new_n161), .b(new_n152), .c(new_n153), .out0(new_n162));
  aoi022aa1n02x5               g067(.a(new_n157), .b(new_n160), .c(new_n151), .d(new_n162), .o1(\s[13] ));
  inv000aa1d42x5               g068(.a(new_n158), .o1(new_n164));
  nanp02aa1n03x5               g069(.a(new_n157), .b(new_n160), .o1(new_n165));
  nor042aa1n06x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanp02aa1n06x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  nona23aa1n02x4               g073(.a(new_n165), .b(new_n167), .c(new_n166), .d(new_n158), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n168), .c(new_n164), .d(new_n165), .o1(\s[14] ));
  nano23aa1n06x5               g075(.a(new_n158), .b(new_n166), .c(new_n167), .d(new_n159), .out0(new_n171));
  oaoi03aa1n02x5               g076(.a(\a[14] ), .b(\b[13] ), .c(new_n164), .o1(new_n172));
  nor022aa1n16x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n08x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x7               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n172), .c(new_n157), .d(new_n171), .o1(new_n176));
  aoi112aa1n02x5               g081(.a(new_n175), .b(new_n172), .c(new_n157), .d(new_n171), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(\s[15] ));
  inv000aa1d42x5               g083(.a(new_n173), .o1(new_n179));
  nor042aa1n02x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nand42aa1n03x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  norb02aa1n03x4               g086(.a(new_n181), .b(new_n180), .out0(new_n182));
  norb03aa1n02x5               g087(.a(new_n181), .b(new_n173), .c(new_n180), .out0(new_n183));
  nand22aa1n03x5               g088(.a(new_n176), .b(new_n183), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n182), .c(new_n176), .d(new_n179), .o1(\s[16] ));
  nano23aa1n02x4               g090(.a(new_n138), .b(new_n144), .c(new_n145), .d(new_n139), .out0(new_n186));
  nano23aa1n03x5               g091(.a(new_n173), .b(new_n180), .c(new_n181), .d(new_n174), .out0(new_n187));
  nand02aa1n02x5               g092(.a(new_n187), .b(new_n171), .o1(new_n188));
  nano22aa1n03x7               g093(.a(new_n188), .b(new_n135), .c(new_n186), .out0(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n190));
  nona23aa1n03x5               g095(.a(new_n167), .b(new_n159), .c(new_n158), .d(new_n166), .out0(new_n191));
  nano22aa1n03x7               g096(.a(new_n191), .b(new_n175), .c(new_n182), .out0(new_n192));
  nanb03aa1n03x5               g097(.a(new_n180), .b(new_n181), .c(new_n174), .out0(new_n193));
  oai112aa1n02x7               g098(.a(new_n179), .b(new_n167), .c(new_n166), .d(new_n158), .o1(new_n194));
  oaih12aa1n02x5               g099(.a(new_n181), .b(new_n180), .c(new_n173), .o1(new_n195));
  oai012aa1n02x7               g100(.a(new_n195), .b(new_n194), .c(new_n193), .o1(new_n196));
  aoi012aa1d18x5               g101(.a(new_n196), .b(new_n155), .c(new_n192), .o1(new_n197));
  nand02aa1d12x5               g102(.a(new_n190), .b(new_n197), .o1(new_n198));
  xorc02aa1n02x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  xnrc02aa1n02x5               g104(.a(\b[16] ), .b(\a[17] ), .out0(new_n200));
  oai112aa1n02x5               g105(.a(new_n195), .b(new_n200), .c(new_n194), .d(new_n193), .o1(new_n201));
  aoi012aa1n02x5               g106(.a(new_n201), .b(new_n155), .c(new_n192), .o1(new_n202));
  aoi022aa1n02x5               g107(.a(new_n198), .b(new_n199), .c(new_n202), .d(new_n190), .o1(\s[17] ));
  nor042aa1n03x5               g108(.a(\b[16] ), .b(\a[17] ), .o1(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  nanp02aa1n06x5               g110(.a(new_n198), .b(new_n199), .o1(new_n206));
  tech160nm_fixorc02aa1n03p5x5 g111(.a(\a[18] ), .b(\b[17] ), .out0(new_n207));
  nand02aa1n03x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  oai022aa1d24x5               g113(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n209));
  nanb03aa1n03x5               g114(.a(new_n209), .b(new_n206), .c(new_n208), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n205), .d(new_n206), .o1(\s[18] ));
  norb02aa1n02x5               g116(.a(new_n207), .b(new_n200), .out0(new_n212));
  oaoi03aa1n02x5               g117(.a(\a[18] ), .b(\b[17] ), .c(new_n205), .o1(new_n213));
  tech160nm_fixorc02aa1n03p5x5 g118(.a(\a[19] ), .b(\b[18] ), .out0(new_n214));
  aoai13aa1n06x5               g119(.a(new_n214), .b(new_n213), .c(new_n198), .d(new_n212), .o1(new_n215));
  aoi112aa1n02x7               g120(.a(new_n214), .b(new_n213), .c(new_n198), .d(new_n212), .o1(new_n216));
  norb02aa1n03x4               g121(.a(new_n215), .b(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  inv000aa1n02x5               g124(.a(new_n219), .o1(new_n220));
  tech160nm_fixorc02aa1n03p5x5 g125(.a(\a[20] ), .b(\b[19] ), .out0(new_n221));
  nand02aa1d28x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  oai022aa1n03x5               g128(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n224));
  nona22aa1n03x5               g129(.a(new_n215), .b(new_n223), .c(new_n224), .out0(new_n225));
  aoai13aa1n03x5               g130(.a(new_n225), .b(new_n221), .c(new_n220), .d(new_n215), .o1(\s[20] ));
  nano32aa1n06x5               g131(.a(new_n200), .b(new_n221), .c(new_n207), .d(new_n214), .out0(new_n227));
  inv000aa1d42x5               g132(.a(\a[19] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\b[18] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\a[20] ), .o1(new_n230));
  nanb02aa1n03x5               g135(.a(\b[19] ), .b(new_n230), .out0(new_n231));
  oai112aa1n04x5               g136(.a(new_n231), .b(new_n222), .c(new_n229), .d(new_n228), .o1(new_n232));
  oai112aa1n03x5               g137(.a(new_n209), .b(new_n208), .c(\b[18] ), .d(\a[19] ), .o1(new_n233));
  nand42aa1n02x5               g138(.a(new_n224), .b(new_n222), .o1(new_n234));
  oai012aa1n06x5               g139(.a(new_n234), .b(new_n233), .c(new_n232), .o1(new_n235));
  xorc02aa1n02x5               g140(.a(\a[21] ), .b(\b[20] ), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n235), .c(new_n198), .d(new_n227), .o1(new_n237));
  nano32aa1n02x4               g142(.a(new_n232), .b(new_n209), .c(new_n220), .d(new_n208), .out0(new_n238));
  nona22aa1n02x4               g143(.a(new_n234), .b(new_n238), .c(new_n236), .out0(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n198), .c(new_n227), .o1(new_n240));
  norb02aa1n03x4               g145(.a(new_n237), .b(new_n240), .out0(\s[21] ));
  inv000aa1d42x5               g146(.a(\a[21] ), .o1(new_n242));
  nanb02aa1n02x5               g147(.a(\b[20] ), .b(new_n242), .out0(new_n243));
  xorc02aa1n02x5               g148(.a(\a[22] ), .b(\b[21] ), .out0(new_n244));
  and002aa1n02x5               g149(.a(\b[21] ), .b(\a[22] ), .o(new_n245));
  oai022aa1n02x5               g150(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n246));
  nona22aa1n03x5               g151(.a(new_n237), .b(new_n245), .c(new_n246), .out0(new_n247));
  aoai13aa1n03x5               g152(.a(new_n247), .b(new_n244), .c(new_n243), .d(new_n237), .o1(\s[22] ));
  inv000aa1n02x5               g153(.a(new_n227), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\a[22] ), .o1(new_n250));
  xroi22aa1d06x4               g155(.a(new_n242), .b(\b[20] ), .c(new_n250), .d(\b[21] ), .out0(new_n251));
  norb02aa1n02x5               g156(.a(new_n251), .b(new_n249), .out0(new_n252));
  oaoi03aa1n02x5               g157(.a(\a[22] ), .b(\b[21] ), .c(new_n243), .o1(new_n253));
  tech160nm_fiao0012aa1n02p5x5 g158(.a(new_n253), .b(new_n235), .c(new_n251), .o(new_n254));
  xorc02aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n198), .d(new_n252), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n255), .b(new_n253), .c(new_n235), .d(new_n251), .o1(new_n257));
  aobi12aa1n02x5               g162(.a(new_n257), .b(new_n198), .c(new_n252), .out0(new_n258));
  norb02aa1n03x4               g163(.a(new_n256), .b(new_n258), .out0(\s[23] ));
  norp02aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  and002aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .o(new_n263));
  oai022aa1n02x5               g168(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n264));
  nona22aa1n03x5               g169(.a(new_n256), .b(new_n263), .c(new_n264), .out0(new_n265));
  aoai13aa1n03x5               g170(.a(new_n265), .b(new_n262), .c(new_n261), .d(new_n256), .o1(\s[24] ));
  inv000aa1d42x5               g171(.a(\a[23] ), .o1(new_n267));
  inv040aa1d32x5               g172(.a(\a[24] ), .o1(new_n268));
  xroi22aa1d06x4               g173(.a(new_n267), .b(\b[22] ), .c(new_n268), .d(\b[23] ), .out0(new_n269));
  nano22aa1n02x4               g174(.a(new_n249), .b(new_n251), .c(new_n269), .out0(new_n270));
  oaib12aa1n02x5               g175(.a(new_n264), .b(new_n268), .c(\b[23] ), .out0(new_n271));
  aoai13aa1n02x5               g176(.a(new_n269), .b(new_n253), .c(new_n235), .d(new_n251), .o1(new_n272));
  nanp02aa1n02x5               g177(.a(new_n272), .b(new_n271), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n198), .d(new_n270), .o1(new_n275));
  nanb02aa1n02x5               g180(.a(new_n274), .b(new_n271), .out0(new_n276));
  aoi122aa1n02x7               g181(.a(new_n276), .b(new_n254), .c(new_n269), .d(new_n198), .e(new_n270), .o1(new_n277));
  norb02aa1n03x4               g182(.a(new_n275), .b(new_n277), .out0(\s[25] ));
  norp02aa1n02x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  tech160nm_fixorc02aa1n05x5   g185(.a(\a[26] ), .b(\b[25] ), .out0(new_n281));
  and002aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .o(new_n282));
  oai022aa1n02x5               g187(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n283));
  nona22aa1n03x5               g188(.a(new_n275), .b(new_n282), .c(new_n283), .out0(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n281), .c(new_n280), .d(new_n275), .o1(\s[26] ));
  nanp02aa1n02x5               g190(.a(new_n244), .b(new_n236), .o1(new_n286));
  nand22aa1n03x5               g191(.a(new_n281), .b(new_n274), .o1(new_n287));
  nona23aa1n03x5               g192(.a(new_n227), .b(new_n269), .c(new_n287), .d(new_n286), .out0(new_n288));
  nanb02aa1n02x5               g193(.a(new_n288), .b(new_n198), .out0(new_n289));
  aoi012aa1n12x5               g194(.a(new_n288), .b(new_n190), .c(new_n197), .o1(new_n290));
  aob012aa1n02x5               g195(.a(new_n283), .b(\b[25] ), .c(\a[26] ), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n287), .c(new_n272), .d(new_n271), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  oai012aa1n06x5               g198(.a(new_n293), .b(new_n292), .c(new_n290), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n282), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n287), .o1(new_n296));
  aoi122aa1n02x5               g201(.a(new_n293), .b(new_n295), .c(new_n283), .d(new_n273), .e(new_n296), .o1(new_n297));
  aobi12aa1n02x7               g202(.a(new_n294), .b(new_n297), .c(new_n289), .out0(\s[27] ));
  norp02aa1n02x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .out0(new_n301));
  oai022aa1n02x5               g206(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n302));
  aoi012aa1n02x5               g207(.a(new_n302), .b(\a[28] ), .c(\b[27] ), .o1(new_n303));
  nanp02aa1n06x5               g208(.a(new_n294), .b(new_n303), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n294), .d(new_n300), .o1(\s[28] ));
  xorc02aa1n12x5               g210(.a(\a[29] ), .b(\b[28] ), .out0(new_n306));
  and002aa1n02x5               g211(.a(new_n301), .b(new_n293), .o(new_n307));
  tech160nm_fioai012aa1n02p5x5 g212(.a(new_n307), .b(new_n292), .c(new_n290), .o1(new_n308));
  aob012aa1n02x5               g213(.a(new_n302), .b(\b[27] ), .c(\a[28] ), .out0(new_n309));
  inv000aa1d42x5               g214(.a(new_n309), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n306), .o1(new_n311));
  nona22aa1n03x5               g216(.a(new_n308), .b(new_n310), .c(new_n311), .out0(new_n312));
  oaoi13aa1n02x7               g217(.a(new_n310), .b(new_n307), .c(new_n292), .d(new_n290), .o1(new_n313));
  oai012aa1n03x5               g218(.a(new_n312), .b(new_n313), .c(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g220(.a(new_n311), .b(new_n293), .c(new_n301), .out0(new_n316));
  oaoi03aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .o1(new_n317));
  oaoi13aa1n02x7               g222(.a(new_n317), .b(new_n316), .c(new_n292), .d(new_n290), .o1(new_n318));
  norp02aa1n02x5               g223(.a(\b[29] ), .b(\a[30] ), .o1(new_n319));
  nanp02aa1n02x5               g224(.a(\b[29] ), .b(\a[30] ), .o1(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(new_n321));
  tech160nm_fioai012aa1n02p5x5 g226(.a(new_n316), .b(new_n292), .c(new_n290), .o1(new_n322));
  and002aa1n02x5               g227(.a(\b[29] ), .b(\a[30] ), .o(new_n323));
  nona32aa1n03x5               g228(.a(new_n322), .b(new_n323), .c(new_n319), .d(new_n317), .out0(new_n324));
  tech160nm_fioai012aa1n02p5x5 g229(.a(new_n324), .b(new_n318), .c(new_n321), .o1(\s[30] ));
  nano32aa1n02x4               g230(.a(new_n311), .b(new_n301), .c(new_n293), .d(new_n321), .out0(new_n326));
  oaih12aa1n02x5               g231(.a(new_n326), .b(new_n292), .c(new_n290), .o1(new_n327));
  oai012aa1n02x5               g232(.a(new_n309), .b(\b[28] ), .c(\a[29] ), .o1(new_n328));
  nanp02aa1n02x5               g233(.a(\b[28] ), .b(\a[29] ), .o1(new_n329));
  nano22aa1n02x4               g234(.a(new_n319), .b(new_n329), .c(new_n320), .out0(new_n330));
  aoi012aa1n02x5               g235(.a(new_n319), .b(\a[31] ), .c(\b[30] ), .o1(new_n331));
  oai012aa1n02x5               g236(.a(new_n331), .b(\b[30] ), .c(\a[31] ), .o1(new_n332));
  aoi012aa1n02x5               g237(.a(new_n332), .b(new_n328), .c(new_n330), .o1(new_n333));
  nanp02aa1n03x5               g238(.a(new_n327), .b(new_n333), .o1(new_n334));
  aoi012aa1n02x5               g239(.a(new_n319), .b(new_n328), .c(new_n330), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n334), .b(new_n336), .c(new_n327), .d(new_n335), .o1(\s[31] ));
  nanp02aa1n02x5               g242(.a(new_n100), .b(new_n99), .o1(new_n338));
  nanp02aa1n02x5               g243(.a(\b[1] ), .b(\a[2] ), .o1(new_n339));
  nanp03aa1n02x5               g244(.a(new_n338), .b(new_n101), .c(new_n339), .o1(new_n340));
  norb02aa1n02x5               g245(.a(new_n106), .b(new_n105), .out0(new_n341));
  xnbna2aa1n03x5               g246(.a(new_n341), .b(new_n340), .c(new_n338), .out0(\s[3] ));
  inv000aa1d42x5               g247(.a(new_n102), .o1(new_n343));
  oaoi03aa1n02x5               g248(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n344));
  oaib12aa1n02x5               g249(.a(new_n344), .b(new_n103), .c(new_n104), .out0(new_n345));
  nona22aa1n02x4               g250(.a(new_n104), .b(new_n105), .c(new_n103), .out0(new_n346));
  aoai13aa1n02x5               g251(.a(new_n345), .b(new_n346), .c(new_n341), .d(new_n343), .o1(\s[4] ));
  nanb02aa1n02x5               g252(.a(new_n107), .b(new_n343), .out0(new_n348));
  norb02aa1n02x5               g253(.a(new_n117), .b(new_n116), .out0(new_n349));
  xnbna2aa1n03x5               g254(.a(new_n349), .b(new_n348), .c(new_n108), .out0(\s[5] ));
  nanb02aa1n02x5               g255(.a(new_n115), .b(new_n114), .out0(new_n351));
  aoai13aa1n02x5               g256(.a(new_n351), .b(new_n116), .c(new_n109), .d(new_n117), .o1(new_n352));
  nona22aa1n02x4               g257(.a(new_n114), .b(new_n115), .c(new_n116), .out0(new_n353));
  aoai13aa1n02x5               g258(.a(new_n352), .b(new_n353), .c(new_n349), .d(new_n109), .o1(\s[6] ));
  oai012aa1n02x5               g259(.a(new_n114), .b(new_n116), .c(new_n115), .o1(new_n355));
  nanb02aa1n02x5               g260(.a(new_n118), .b(new_n109), .out0(new_n356));
  xobna2aa1n03x5               g261(.a(new_n113), .b(new_n356), .c(new_n355), .out0(\s[7] ));
  orn002aa1n02x5               g262(.a(\a[7] ), .b(\b[6] ), .o(new_n358));
  tech160nm_fiao0012aa1n02p5x5 g263(.a(new_n113), .b(new_n356), .c(new_n355), .o(new_n359));
  xobna2aa1n03x5               g264(.a(new_n110), .b(new_n359), .c(new_n358), .out0(\s[8] ));
  oaoi13aa1n02x5               g265(.a(new_n127), .b(new_n120), .c(new_n123), .d(new_n111), .o1(new_n361));
  oaib12aa1n02x5               g266(.a(new_n361), .b(new_n122), .c(new_n121), .out0(new_n362));
  aoi012aa1n02x5               g267(.a(new_n362), .b(new_n109), .c(new_n119), .o1(new_n363));
  norb02aa1n02x5               g268(.a(new_n128), .b(new_n363), .out0(\s[9] ));
endmodule


