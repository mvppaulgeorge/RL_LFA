// Benchmark "adder" written by ABC on Thu Jul 18 15:02:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n317, new_n318, new_n320,
    new_n321, new_n322, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand02aa1d04x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  tech160nm_fioai012aa1n05x5   g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  nor022aa1n08x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  tech160nm_fiaoi012aa1n03p5x5 g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  oaih12aa1n06x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  nor022aa1n04x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nanp02aa1n04x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n09x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .out0(new_n113));
  tech160nm_fixnrc02aa1n02p5x5 g018(.a(\b[7] ), .b(\a[8] ), .out0(new_n114));
  nor043aa1n03x5               g019(.a(new_n112), .b(new_n113), .c(new_n114), .o1(new_n115));
  oai022aa1n02x5               g020(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n116));
  nano22aa1n03x7               g021(.a(new_n110), .b(new_n109), .c(new_n111), .out0(new_n117));
  nand02aa1n03x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  oab012aa1d30x5               g023(.a(new_n110), .b(\a[8] ), .c(\b[7] ), .out0(new_n119));
  aoi022aa1n06x5               g024(.a(new_n118), .b(new_n119), .c(\b[7] ), .d(\a[8] ), .o1(new_n120));
  tech160nm_fiaoi012aa1n05x5   g025(.a(new_n120), .b(new_n107), .c(new_n115), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .c(new_n121), .o1(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  tech160nm_fixnrc02aa1n04x5   g028(.a(\b[8] ), .b(\a[9] ), .out0(new_n124));
  and002aa1n02x5               g029(.a(\b[9] ), .b(\a[10] ), .o(new_n125));
  inv000aa1d42x5               g030(.a(\a[10] ), .o1(new_n126));
  inv040aa1d32x5               g031(.a(\b[9] ), .o1(new_n127));
  nor002aa1d32x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  aoi012aa1n02x7               g033(.a(new_n128), .b(new_n126), .c(new_n127), .o1(new_n129));
  oaoi13aa1n04x5               g034(.a(new_n125), .b(new_n129), .c(new_n121), .d(new_n124), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  aoi012aa1n02x5               g038(.a(new_n132), .b(new_n130), .c(new_n133), .o1(new_n134));
  xnrb03aa1n03x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nand22aa1n06x5               g040(.a(new_n107), .b(new_n115), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(\b[7] ), .b(\a[8] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n119), .o1(new_n138));
  aoai13aa1n06x5               g043(.a(new_n137), .b(new_n138), .c(new_n117), .d(new_n116), .o1(new_n139));
  xnrc02aa1n02x5               g044(.a(\b[9] ), .b(\a[10] ), .out0(new_n140));
  nor022aa1n16x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanp02aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nano23aa1n03x7               g047(.a(new_n132), .b(new_n141), .c(new_n142), .d(new_n133), .out0(new_n143));
  nona22aa1n02x4               g048(.a(new_n143), .b(new_n140), .c(new_n124), .out0(new_n144));
  nona23aa1n09x5               g049(.a(new_n142), .b(new_n133), .c(new_n132), .d(new_n141), .out0(new_n145));
  oaoi03aa1n06x5               g050(.a(new_n126), .b(new_n127), .c(new_n128), .o1(new_n146));
  oa0012aa1n06x5               g051(.a(new_n142), .b(new_n141), .c(new_n132), .o(new_n147));
  oabi12aa1n18x5               g052(.a(new_n147), .b(new_n145), .c(new_n146), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n144), .c(new_n136), .d(new_n139), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1n10x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n152), .b(new_n150), .c(new_n153), .o1(new_n154));
  xnrb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor043aa1n03x5               g060(.a(new_n145), .b(new_n140), .c(new_n124), .o1(new_n156));
  aoai13aa1n03x5               g061(.a(new_n156), .b(new_n120), .c(new_n107), .d(new_n115), .o1(new_n157));
  nor042aa1n04x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand42aa1n16x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nano23aa1d15x5               g064(.a(new_n152), .b(new_n158), .c(new_n159), .d(new_n153), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoi012aa1d18x5               g066(.a(new_n158), .b(new_n152), .c(new_n159), .o1(new_n162));
  aoai13aa1n04x5               g067(.a(new_n162), .b(new_n161), .c(new_n157), .d(new_n149), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand42aa1n04x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nor042aa1n04x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nanp02aa1n06x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  nanb02aa1n02x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n170));
  aoi112aa1n02x7               g075(.a(new_n165), .b(new_n169), .c(new_n163), .d(new_n166), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(\s[16] ));
  nano23aa1d15x5               g077(.a(new_n165), .b(new_n167), .c(new_n168), .d(new_n166), .out0(new_n173));
  nano22aa1n03x7               g078(.a(new_n144), .b(new_n160), .c(new_n173), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n120), .c(new_n107), .d(new_n115), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n162), .o1(new_n176));
  aoai13aa1n12x5               g081(.a(new_n173), .b(new_n176), .c(new_n148), .d(new_n160), .o1(new_n177));
  oaih12aa1n06x5               g082(.a(new_n168), .b(new_n167), .c(new_n165), .o1(new_n178));
  nand23aa1n06x5               g083(.a(new_n175), .b(new_n177), .c(new_n178), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g085(.a(\a[18] ), .o1(new_n181));
  nand23aa1n03x5               g086(.a(new_n156), .b(new_n160), .c(new_n173), .o1(new_n182));
  aoi012aa1d18x5               g087(.a(new_n182), .b(new_n136), .c(new_n139), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n173), .o1(new_n184));
  norp02aa1n02x5               g089(.a(new_n129), .b(new_n125), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n160), .b(new_n147), .c(new_n143), .d(new_n185), .o1(new_n186));
  aoai13aa1n12x5               g091(.a(new_n178), .b(new_n184), .c(new_n186), .d(new_n162), .o1(new_n187));
  nor042aa1n02x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  tech160nm_fixorc02aa1n03p5x5 g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  oaoi13aa1n06x5               g094(.a(new_n188), .b(new_n189), .c(new_n187), .d(new_n183), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  nor002aa1n06x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nand22aa1n04x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  nano22aa1n06x5               g098(.a(new_n192), .b(new_n189), .c(new_n193), .out0(new_n194));
  tech160nm_fioai012aa1n05x5   g099(.a(new_n194), .b(new_n187), .c(new_n183), .o1(new_n195));
  aoi012aa1n12x5               g100(.a(new_n192), .b(new_n188), .c(new_n193), .o1(new_n196));
  nor042aa1n06x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanp02aa1n04x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n195), .c(new_n196), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g106(.a(new_n195), .b(new_n196), .o1(new_n202));
  nor022aa1n16x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  nand02aa1n08x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(new_n205));
  aoai13aa1n03x5               g110(.a(new_n205), .b(new_n197), .c(new_n202), .d(new_n199), .o1(new_n206));
  inv040aa1n03x5               g111(.a(new_n196), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n199), .b(new_n207), .c(new_n179), .d(new_n194), .o1(new_n208));
  nona22aa1n02x5               g113(.a(new_n208), .b(new_n205), .c(new_n197), .out0(new_n209));
  nanp02aa1n03x5               g114(.a(new_n206), .b(new_n209), .o1(\s[20] ));
  nor042aa1n06x5               g115(.a(new_n187), .b(new_n183), .o1(new_n211));
  nona23aa1n09x5               g116(.a(new_n204), .b(new_n198), .c(new_n197), .d(new_n203), .out0(new_n212));
  nano23aa1n09x5               g117(.a(new_n212), .b(new_n192), .c(new_n189), .d(new_n193), .out0(new_n213));
  inv040aa1n03x5               g118(.a(new_n213), .o1(new_n214));
  oai012aa1d24x5               g119(.a(new_n204), .b(new_n203), .c(new_n197), .o1(new_n215));
  oai012aa1n12x5               g120(.a(new_n215), .b(new_n212), .c(new_n196), .o1(new_n216));
  oabi12aa1n06x5               g121(.a(new_n216), .b(new_n211), .c(new_n214), .out0(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[21] ), .b(\b[20] ), .out0(new_n220));
  xorc02aa1n02x5               g125(.a(\a[22] ), .b(\b[21] ), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n222), .b(new_n219), .c(new_n217), .d(new_n220), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n220), .b(new_n216), .c(new_n179), .d(new_n213), .o1(new_n224));
  nona22aa1n03x5               g129(.a(new_n224), .b(new_n222), .c(new_n219), .out0(new_n225));
  nanp02aa1n02x5               g130(.a(new_n223), .b(new_n225), .o1(\s[22] ));
  nano23aa1n09x5               g131(.a(new_n197), .b(new_n203), .c(new_n204), .d(new_n198), .out0(new_n227));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv040aa1d32x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  nand23aa1n09x5               g135(.a(new_n194), .b(new_n227), .c(new_n230), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n215), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n230), .b(new_n232), .c(new_n227), .d(new_n207), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\b[21] ), .o1(new_n234));
  oao003aa1n02x5               g139(.a(new_n229), .b(new_n234), .c(new_n219), .carry(new_n235));
  inv000aa1n02x5               g140(.a(new_n235), .o1(new_n236));
  nanp02aa1n02x5               g141(.a(new_n233), .b(new_n236), .o1(new_n237));
  oabi12aa1n06x5               g142(.a(new_n237), .b(new_n211), .c(new_n231), .out0(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  xorc02aa1n06x5               g145(.a(\a[23] ), .b(\b[22] ), .out0(new_n241));
  norp02aa1n03x5               g146(.a(\b[23] ), .b(\a[24] ), .o1(new_n242));
  nand42aa1n03x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  nanb02aa1n06x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n240), .c(new_n238), .d(new_n241), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n231), .o1(new_n246));
  aoai13aa1n02x5               g151(.a(new_n241), .b(new_n237), .c(new_n179), .d(new_n246), .o1(new_n247));
  nona22aa1n03x5               g152(.a(new_n247), .b(new_n244), .c(new_n240), .out0(new_n248));
  nanp02aa1n02x5               g153(.a(new_n245), .b(new_n248), .o1(\s[24] ));
  norb02aa1n02x7               g154(.a(new_n241), .b(new_n244), .out0(new_n250));
  nano22aa1n02x4               g155(.a(new_n214), .b(new_n250), .c(new_n230), .out0(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  inv030aa1n02x5               g157(.a(new_n250), .o1(new_n253));
  oai012aa1n02x5               g158(.a(new_n243), .b(new_n242), .c(new_n240), .o1(new_n254));
  aoai13aa1n12x5               g159(.a(new_n254), .b(new_n253), .c(new_n233), .d(new_n236), .o1(new_n255));
  oabi12aa1n06x5               g160(.a(new_n255), .b(new_n211), .c(new_n252), .out0(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  tech160nm_fixorc02aa1n04x5   g163(.a(\a[25] ), .b(\b[24] ), .out0(new_n259));
  nor002aa1n02x5               g164(.a(\b[25] ), .b(\a[26] ), .o1(new_n260));
  nand42aa1n03x5               g165(.a(\b[25] ), .b(\a[26] ), .o1(new_n261));
  norb02aa1n03x4               g166(.a(new_n261), .b(new_n260), .out0(new_n262));
  inv040aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n03x5               g168(.a(new_n263), .b(new_n258), .c(new_n256), .d(new_n259), .o1(new_n264));
  aoai13aa1n02x5               g169(.a(new_n259), .b(new_n255), .c(new_n179), .d(new_n251), .o1(new_n265));
  nona22aa1n03x5               g170(.a(new_n265), .b(new_n263), .c(new_n258), .out0(new_n266));
  nanp02aa1n02x5               g171(.a(new_n264), .b(new_n266), .o1(\s[26] ));
  norb02aa1n12x5               g172(.a(new_n259), .b(new_n263), .out0(new_n268));
  nano22aa1d15x5               g173(.a(new_n231), .b(new_n250), .c(new_n268), .out0(new_n269));
  oai012aa1n18x5               g174(.a(new_n269), .b(new_n187), .c(new_n183), .o1(new_n270));
  oai012aa1n02x5               g175(.a(new_n261), .b(new_n260), .c(new_n258), .o1(new_n271));
  aobi12aa1n12x5               g176(.a(new_n271), .b(new_n255), .c(new_n268), .out0(new_n272));
  xorc02aa1n02x5               g177(.a(\a[27] ), .b(\b[26] ), .out0(new_n273));
  xnbna2aa1n03x5               g178(.a(new_n273), .b(new_n272), .c(new_n270), .out0(\s[27] ));
  nanp02aa1n06x5               g179(.a(new_n272), .b(new_n270), .o1(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  norp02aa1n02x5               g181(.a(\b[27] ), .b(\a[28] ), .o1(new_n277));
  nand42aa1n03x5               g182(.a(\b[27] ), .b(\a[28] ), .o1(new_n278));
  norb02aa1n03x5               g183(.a(new_n278), .b(new_n277), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n276), .c(new_n275), .d(new_n273), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n250), .b(new_n235), .c(new_n216), .d(new_n230), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n268), .o1(new_n283));
  aoai13aa1n04x5               g188(.a(new_n271), .b(new_n283), .c(new_n282), .d(new_n254), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n273), .b(new_n284), .c(new_n179), .d(new_n269), .o1(new_n285));
  nona22aa1n02x5               g190(.a(new_n285), .b(new_n280), .c(new_n276), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n281), .b(new_n286), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n273), .b(new_n280), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n284), .c(new_n179), .d(new_n269), .o1(new_n289));
  aoi012aa1n02x5               g194(.a(new_n277), .b(new_n276), .c(new_n278), .o1(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  aobi12aa1n06x5               g197(.a(new_n288), .b(new_n272), .c(new_n270), .out0(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n291), .out0(new_n294));
  nor002aa1n02x5               g199(.a(new_n292), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g201(.a(new_n291), .b(new_n273), .c(new_n279), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n284), .c(new_n179), .d(new_n269), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[29] ), .b(\a[30] ), .out0(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n298), .c(new_n299), .o1(new_n301));
  aobi12aa1n06x5               g206(.a(new_n297), .b(new_n272), .c(new_n270), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n299), .c(new_n300), .out0(new_n303));
  nor002aa1n02x5               g208(.a(new_n301), .b(new_n303), .o1(\s[30] ));
  nano23aa1n03x7               g209(.a(new_n300), .b(new_n291), .c(new_n273), .d(new_n279), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n284), .c(new_n179), .d(new_n269), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  aobi12aa1n06x5               g214(.a(new_n305), .b(new_n272), .c(new_n270), .out0(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n307), .c(new_n308), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[31] ));
  xnrb03aa1n02x5               g217(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g218(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g220(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norp02aa1n02x5               g221(.a(\b[4] ), .b(\a[5] ), .o1(new_n317));
  aoib12aa1n02x5               g222(.a(new_n317), .b(new_n107), .c(new_n113), .out0(new_n318));
  xnrb03aa1n02x5               g223(.a(new_n318), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g224(.a(new_n110), .o1(new_n320));
  nanb03aa1n02x5               g225(.a(new_n108), .b(new_n318), .c(new_n109), .out0(new_n321));
  aoi022aa1n02x5               g226(.a(new_n321), .b(new_n109), .c(new_n320), .d(new_n111), .o1(new_n322));
  nanp02aa1n02x5               g227(.a(new_n321), .b(new_n117), .o1(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(\s[7] ));
  xobna2aa1n03x5               g229(.a(new_n114), .b(new_n323), .c(new_n320), .out0(\s[8] ));
  xobna2aa1n03x5               g230(.a(new_n124), .b(new_n136), .c(new_n139), .out0(\s[9] ));
endmodule


