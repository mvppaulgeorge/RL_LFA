// Benchmark "adder" written by ABC on Wed Jul 17 21:35:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n317,
    new_n320, new_n321, new_n323, new_n324, new_n326, new_n327, new_n328,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  tech160nm_fioai012aa1n05x5   g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  nor022aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1d04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n08x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  tech160nm_fiaoi012aa1n03p5x5 g012(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n108));
  oai012aa1n09x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nor022aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand22aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor022aa1n08x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1d18x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  nor043aa1n04x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  tech160nm_fioai012aa1n03p5x5 g022(.a(new_n111), .b(new_n112), .c(new_n110), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[5] ), .o1(new_n119));
  oai022aa1n02x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  oaib12aa1n03x5               g025(.a(new_n120), .b(new_n119), .c(\a[6] ), .out0(new_n121));
  oai012aa1n12x5               g026(.a(new_n118), .b(new_n114), .c(new_n121), .o1(new_n122));
  and002aa1n02x5               g027(.a(\b[8] ), .b(\a[9] ), .o(new_n123));
  norp02aa1n02x5               g028(.a(new_n123), .b(new_n97), .o1(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n125));
  nor042aa1n06x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand42aa1d28x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1n02x7               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  nor042aa1n06x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nand22aa1n12x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nona22aa1n03x5               g037(.a(new_n125), .b(new_n126), .c(new_n97), .out0(new_n133));
  nona23aa1n03x5               g038(.a(new_n133), .b(new_n127), .c(new_n130), .d(new_n132), .out0(new_n134));
  inv040aa1n04x5               g039(.a(new_n130), .o1(new_n135));
  aoi022aa1n02x5               g040(.a(new_n133), .b(new_n127), .c(new_n135), .d(new_n131), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n134), .b(new_n136), .out0(\s[11] ));
  nor042aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n134), .c(new_n135), .out0(\s[12] ));
  nanb03aa1n12x5               g046(.a(new_n138), .b(new_n139), .c(new_n131), .out0(new_n142));
  nano32aa1n02x4               g047(.a(new_n142), .b(new_n124), .c(new_n128), .d(new_n135), .out0(new_n143));
  aoai13aa1n03x5               g048(.a(new_n143), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n144));
  oai112aa1n06x5               g049(.a(new_n135), .b(new_n127), .c(new_n126), .d(new_n97), .o1(new_n145));
  oaoi03aa1n09x5               g050(.a(\a[12] ), .b(\b[11] ), .c(new_n135), .o1(new_n146));
  oabi12aa1n18x5               g051(.a(new_n146), .b(new_n145), .c(new_n142), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n144), .b(new_n148), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1d28x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  aoi012aa1n02x5               g057(.a(new_n151), .b(new_n149), .c(new_n152), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nand42aa1d28x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  aoi012aa1n12x5               g061(.a(new_n155), .b(new_n151), .c(new_n156), .o1(new_n157));
  nano23aa1d15x5               g062(.a(new_n151), .b(new_n155), .c(new_n156), .d(new_n152), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n157), .b(new_n159), .c(new_n144), .d(new_n148), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nand02aa1n03x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nor002aa1n03x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nand02aa1n03x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  aoai13aa1n02x7               g071(.a(new_n166), .b(new_n162), .c(new_n160), .d(new_n163), .o1(new_n167));
  aoi112aa1n02x5               g072(.a(new_n166), .b(new_n162), .c(new_n160), .d(new_n163), .o1(new_n168));
  norb02aa1n03x4               g073(.a(new_n167), .b(new_n168), .out0(\s[16] ));
  nano22aa1n03x7               g074(.a(new_n138), .b(new_n131), .c(new_n139), .out0(new_n170));
  nona32aa1n03x5               g075(.a(new_n128), .b(new_n123), .c(new_n130), .d(new_n97), .out0(new_n171));
  nona23aa1d16x5               g076(.a(new_n165), .b(new_n163), .c(new_n162), .d(new_n164), .out0(new_n172));
  nano23aa1d12x5               g077(.a(new_n171), .b(new_n172), .c(new_n158), .d(new_n170), .out0(new_n173));
  aoai13aa1n06x5               g078(.a(new_n173), .b(new_n122), .c(new_n109), .d(new_n117), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n157), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n172), .o1(new_n176));
  aoai13aa1n12x5               g081(.a(new_n176), .b(new_n175), .c(new_n147), .d(new_n158), .o1(new_n177));
  tech160nm_fiaoi012aa1n05x5   g082(.a(new_n164), .b(new_n162), .c(new_n165), .o1(new_n178));
  nanp03aa1d12x5               g083(.a(new_n174), .b(new_n177), .c(new_n178), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n03x5               g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  inv040aa1n02x5               g090(.a(new_n122), .o1(new_n186));
  aob012aa1d15x5               g091(.a(new_n186), .b(new_n109), .c(new_n117), .out0(new_n187));
  oai012aa1n02x5               g092(.a(new_n127), .b(\b[10] ), .c(\a[11] ), .o1(new_n188));
  oab012aa1n02x4               g093(.a(new_n188), .b(new_n97), .c(new_n126), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n158), .b(new_n146), .c(new_n189), .d(new_n170), .o1(new_n190));
  aoai13aa1n06x5               g095(.a(new_n178), .b(new_n172), .c(new_n190), .d(new_n157), .o1(new_n191));
  xroi22aa1d06x4               g096(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n191), .c(new_n187), .d(new_n173), .o1(new_n193));
  oaih22aa1d12x5               g098(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n194));
  oaib12aa1n18x5               g099(.a(new_n194), .b(new_n181), .c(\b[17] ), .out0(new_n195));
  nor002aa1d24x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nand02aa1d08x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanb02aa1d24x5               g102(.a(new_n196), .b(new_n197), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n193), .c(new_n195), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g106(.a(new_n196), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n195), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n199), .b(new_n203), .c(new_n179), .d(new_n192), .o1(new_n204));
  nor002aa1d24x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand02aa1n04x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  tech160nm_fiaoi012aa1n02p5x5 g112(.a(new_n207), .b(new_n204), .c(new_n202), .o1(new_n208));
  aoi012aa1n02x5               g113(.a(new_n198), .b(new_n193), .c(new_n195), .o1(new_n209));
  nano22aa1n02x4               g114(.a(new_n209), .b(new_n202), .c(new_n207), .out0(new_n210));
  norp02aa1n03x5               g115(.a(new_n208), .b(new_n210), .o1(\s[20] ));
  nona23aa1d18x5               g116(.a(new_n206), .b(new_n197), .c(new_n196), .d(new_n205), .out0(new_n212));
  inv000aa1n06x5               g117(.a(new_n212), .o1(new_n213));
  nand02aa1d06x5               g118(.a(new_n192), .b(new_n213), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n191), .c(new_n187), .d(new_n173), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n205), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(new_n196), .b(new_n206), .o1(new_n218));
  nor003aa1n03x5               g123(.a(new_n195), .b(new_n198), .c(new_n207), .o1(new_n219));
  nano22aa1n03x7               g124(.a(new_n219), .b(new_n217), .c(new_n218), .out0(new_n220));
  xnrc02aa1n12x5               g125(.a(\b[20] ), .b(\a[21] ), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n216), .c(new_n220), .out0(\s[21] ));
  orn002aa1n02x5               g128(.a(\a[21] ), .b(\b[20] ), .o(new_n224));
  oai112aa1n06x5               g129(.a(new_n218), .b(new_n217), .c(new_n212), .d(new_n195), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n222), .b(new_n225), .c(new_n179), .d(new_n215), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[21] ), .b(\a[22] ), .out0(new_n227));
  tech160nm_fiaoi012aa1n02p5x5 g132(.a(new_n227), .b(new_n226), .c(new_n224), .o1(new_n228));
  aoi012aa1n02x5               g133(.a(new_n221), .b(new_n216), .c(new_n220), .o1(new_n229));
  nano22aa1n02x4               g134(.a(new_n229), .b(new_n224), .c(new_n227), .out0(new_n230));
  nor002aa1n02x5               g135(.a(new_n228), .b(new_n230), .o1(\s[22] ));
  nor042aa1n02x5               g136(.a(new_n227), .b(new_n221), .o1(new_n232));
  and003aa1n02x5               g137(.a(new_n192), .b(new_n213), .c(new_n232), .o(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n191), .c(new_n187), .d(new_n173), .o1(new_n234));
  tech160nm_fioaoi03aa1n03p5x5 g139(.a(\a[22] ), .b(\b[21] ), .c(new_n224), .o1(new_n235));
  tech160nm_fiaoi012aa1n04x5   g140(.a(new_n235), .b(new_n225), .c(new_n232), .o1(new_n236));
  xorc02aa1n12x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  xnbna2aa1n03x5               g142(.a(new_n237), .b(new_n234), .c(new_n236), .out0(\s[23] ));
  inv000aa1d42x5               g143(.a(\a[23] ), .o1(new_n239));
  nanb02aa1n02x5               g144(.a(\b[22] ), .b(new_n239), .out0(new_n240));
  inv020aa1n02x5               g145(.a(new_n236), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n237), .b(new_n241), .c(new_n179), .d(new_n233), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[23] ), .b(\a[24] ), .out0(new_n243));
  tech160nm_fiaoi012aa1n02p5x5 g148(.a(new_n243), .b(new_n242), .c(new_n240), .o1(new_n244));
  aobi12aa1n02x5               g149(.a(new_n237), .b(new_n234), .c(new_n236), .out0(new_n245));
  nano22aa1n02x4               g150(.a(new_n245), .b(new_n240), .c(new_n243), .out0(new_n246));
  norp02aa1n03x5               g151(.a(new_n244), .b(new_n246), .o1(\s[24] ));
  norb02aa1n02x7               g152(.a(new_n237), .b(new_n243), .out0(new_n248));
  nano22aa1n02x4               g153(.a(new_n214), .b(new_n248), .c(new_n232), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n191), .c(new_n187), .d(new_n173), .o1(new_n250));
  norp02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n252));
  nanb03aa1n02x5               g157(.a(new_n243), .b(new_n235), .c(new_n237), .out0(new_n253));
  nona22aa1n02x4               g158(.a(new_n253), .b(new_n252), .c(new_n251), .out0(new_n254));
  aoi013aa1n02x5               g159(.a(new_n254), .b(new_n225), .c(new_n232), .d(new_n248), .o1(new_n255));
  xnrc02aa1n12x5               g160(.a(\b[24] ), .b(\a[25] ), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  xnbna2aa1n03x5               g162(.a(new_n257), .b(new_n250), .c(new_n255), .out0(\s[25] ));
  nor042aa1n03x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  inv020aa1n02x5               g165(.a(new_n255), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n257), .b(new_n261), .c(new_n179), .d(new_n249), .o1(new_n262));
  xnrc02aa1n02x5               g167(.a(\b[25] ), .b(\a[26] ), .out0(new_n263));
  tech160nm_fiaoi012aa1n02p5x5 g168(.a(new_n263), .b(new_n262), .c(new_n260), .o1(new_n264));
  tech160nm_fiaoi012aa1n03p5x5 g169(.a(new_n256), .b(new_n250), .c(new_n255), .o1(new_n265));
  nano22aa1n03x7               g170(.a(new_n265), .b(new_n260), .c(new_n263), .out0(new_n266));
  nor002aa1n02x5               g171(.a(new_n264), .b(new_n266), .o1(\s[26] ));
  norp02aa1n02x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  and002aa1n02x5               g173(.a(\b[26] ), .b(\a[27] ), .o(new_n269));
  norp02aa1n02x5               g174(.a(new_n269), .b(new_n268), .o1(new_n270));
  nor042aa1n02x5               g175(.a(new_n263), .b(new_n256), .o1(new_n271));
  inv000aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  nano23aa1n06x5               g177(.a(new_n214), .b(new_n272), .c(new_n248), .d(new_n232), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n191), .c(new_n187), .d(new_n173), .o1(new_n274));
  nano22aa1n03x7               g179(.a(new_n220), .b(new_n232), .c(new_n248), .out0(new_n275));
  oao003aa1n06x5               g180(.a(\a[26] ), .b(\b[25] ), .c(new_n260), .carry(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  oaoi13aa1n09x5               g182(.a(new_n277), .b(new_n271), .c(new_n275), .d(new_n254), .o1(new_n278));
  xnbna2aa1n06x5               g183(.a(new_n270), .b(new_n274), .c(new_n278), .out0(\s[27] ));
  inv000aa1n06x5               g184(.a(new_n268), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n269), .o1(new_n281));
  nand43aa1n03x5               g186(.a(new_n225), .b(new_n232), .c(new_n248), .o1(new_n282));
  inv000aa1n02x5               g187(.a(new_n254), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n276), .b(new_n272), .c(new_n282), .d(new_n283), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n281), .b(new_n284), .c(new_n179), .d(new_n273), .o1(new_n285));
  xnrc02aa1n02x5               g190(.a(\b[27] ), .b(\a[28] ), .out0(new_n286));
  tech160nm_fiaoi012aa1n02p5x5 g191(.a(new_n286), .b(new_n285), .c(new_n280), .o1(new_n287));
  aoi012aa1n06x5               g192(.a(new_n269), .b(new_n274), .c(new_n278), .o1(new_n288));
  nano22aa1n03x5               g193(.a(new_n288), .b(new_n280), .c(new_n286), .out0(new_n289));
  norp02aa1n03x5               g194(.a(new_n287), .b(new_n289), .o1(\s[28] ));
  nano22aa1n02x4               g195(.a(new_n286), .b(new_n281), .c(new_n280), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n284), .c(new_n179), .d(new_n273), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[28] ), .b(\a[29] ), .out0(new_n294));
  tech160nm_fiaoi012aa1n02p5x5 g199(.a(new_n294), .b(new_n292), .c(new_n293), .o1(new_n295));
  aobi12aa1n06x5               g200(.a(new_n291), .b(new_n274), .c(new_n278), .out0(new_n296));
  nano22aa1n02x4               g201(.a(new_n296), .b(new_n293), .c(new_n294), .out0(new_n297));
  norp02aa1n03x5               g202(.a(new_n295), .b(new_n297), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g204(.a(new_n270), .b(new_n294), .c(new_n286), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n284), .c(new_n179), .d(new_n273), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[29] ), .b(\b[28] ), .c(new_n293), .carry(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[29] ), .b(\a[30] ), .out0(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n301), .c(new_n302), .o1(new_n304));
  aobi12aa1n06x5               g209(.a(new_n300), .b(new_n274), .c(new_n278), .out0(new_n305));
  nano22aa1n02x4               g210(.a(new_n305), .b(new_n302), .c(new_n303), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n304), .b(new_n306), .o1(\s[30] ));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  norb03aa1n02x5               g213(.a(new_n291), .b(new_n303), .c(new_n294), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n284), .c(new_n179), .d(new_n273), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .c(new_n302), .carry(new_n311));
  tech160nm_fiaoi012aa1n02p5x5 g216(.a(new_n308), .b(new_n310), .c(new_n311), .o1(new_n312));
  aobi12aa1n06x5               g217(.a(new_n309), .b(new_n274), .c(new_n278), .out0(new_n313));
  nano22aa1n03x5               g218(.a(new_n313), .b(new_n308), .c(new_n311), .out0(new_n314));
  norp02aa1n03x5               g219(.a(new_n312), .b(new_n314), .o1(\s[31] ));
  xnrb03aa1n02x5               g220(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g221(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g223(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aob012aa1n02x5               g224(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(new_n320));
  tech160nm_fioai012aa1n03p5x5 g225(.a(new_n320), .b(\b[4] ), .c(\a[5] ), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g227(.a(new_n115), .b(new_n321), .out0(new_n323));
  oaib12aa1n06x5               g228(.a(new_n323), .b(\a[6] ), .c(new_n119), .out0(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g230(.a(new_n110), .b(new_n111), .out0(new_n326));
  inv000aa1d42x5               g231(.a(new_n326), .o1(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n112), .c(new_n324), .d(new_n113), .o1(new_n328));
  aoi112aa1n02x5               g233(.a(new_n327), .b(new_n112), .c(new_n324), .d(new_n113), .o1(new_n329));
  norb02aa1n02x7               g234(.a(new_n328), .b(new_n329), .out0(\s[8] ));
  xorb03aa1n02x5               g235(.a(new_n187), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


