// Benchmark "adder" written by ABC on Wed Jul 17 17:06:05 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n320, new_n323, new_n325, new_n326, new_n327,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1n09x5               g002(.a(new_n97), .o1(new_n98));
  norp02aa1n12x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand02aa1d06x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  tech160nm_fiaoi012aa1n03p5x5 g006(.a(new_n99), .b(new_n101), .c(new_n100), .o1(new_n102));
  and002aa1n24x5               g007(.a(\b[5] ), .b(\a[6] ), .o(new_n103));
  nor042aa1d18x5               g008(.a(\b[4] ), .b(\a[5] ), .o1(new_n104));
  oab012aa1n04x5               g009(.a(new_n104), .b(\a[6] ), .c(\b[5] ), .out0(new_n105));
  nand02aa1n04x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  nona23aa1d18x5               g011(.a(new_n106), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n107));
  oai013aa1n09x5               g012(.a(new_n102), .b(new_n107), .c(new_n103), .d(new_n105), .o1(new_n108));
  nand42aa1n02x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  nand22aa1n12x5               g014(.a(\b[0] ), .b(\a[1] ), .o1(new_n110));
  nor042aa1n09x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n109), .b(new_n111), .c(new_n110), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  nand02aa1d06x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nor022aa1n16x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  nanp02aa1n04x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nona23aa1n12x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  tech160nm_fioai012aa1n03p5x5 g022(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n118));
  oaih12aa1n12x5               g023(.a(new_n118), .b(new_n117), .c(new_n112), .o1(new_n119));
  tech160nm_fixnrc02aa1n04x5   g024(.a(\b[5] ), .b(\a[6] ), .out0(new_n120));
  nanp02aa1n04x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nanb02aa1n02x5               g026(.a(new_n104), .b(new_n121), .out0(new_n122));
  nor043aa1d12x5               g027(.a(new_n107), .b(new_n120), .c(new_n122), .o1(new_n123));
  nand42aa1n08x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n97), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n108), .c(new_n123), .d(new_n119), .o1(new_n126));
  nor002aa1n16x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n08x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  aobi12aa1n06x5               g035(.a(new_n129), .b(new_n126), .c(new_n98), .out0(new_n131));
  nanp02aa1n24x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n132), .b(new_n133), .out0(new_n134));
  tech160nm_fioaoi03aa1n02p5x5 g039(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n135));
  oai012aa1n06x5               g040(.a(new_n134), .b(new_n131), .c(new_n135), .o1(new_n136));
  nanb02aa1d24x5               g041(.a(new_n133), .b(new_n132), .out0(new_n137));
  tech160nm_fioai012aa1n05x5   g042(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n138));
  nano22aa1n02x4               g043(.a(new_n131), .b(new_n137), .c(new_n138), .out0(new_n139));
  norb02aa1n02x5               g044(.a(new_n136), .b(new_n139), .out0(\s[11] ));
  nor042aa1n09x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand02aa1d28x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  nona22aa1n02x5               g048(.a(new_n136), .b(new_n143), .c(new_n133), .out0(new_n144));
  inv000aa1d42x5               g049(.a(new_n133), .o1(new_n145));
  nanb02aa1d36x5               g050(.a(new_n141), .b(new_n142), .out0(new_n146));
  tech160nm_fiaoi012aa1n03p5x5 g051(.a(new_n146), .b(new_n136), .c(new_n145), .o1(new_n147));
  norb02aa1n03x4               g052(.a(new_n144), .b(new_n147), .out0(\s[12] ));
  nano23aa1d18x5               g053(.a(new_n97), .b(new_n127), .c(new_n128), .d(new_n124), .out0(new_n149));
  nona22aa1n09x5               g054(.a(new_n149), .b(new_n146), .c(new_n137), .out0(new_n150));
  inv040aa1n02x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n108), .c(new_n123), .d(new_n119), .o1(new_n152));
  aoi012aa1n02x7               g057(.a(new_n141), .b(new_n133), .c(new_n142), .o1(new_n153));
  oai013aa1d12x5               g058(.a(new_n153), .b(new_n138), .c(new_n137), .d(new_n146), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  nand42aa1n20x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nor042aa1n02x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  norb02aa1n06x5               g062(.a(new_n156), .b(new_n157), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n152), .c(new_n155), .out0(\s[13] ));
  inv030aa1d32x5               g064(.a(\a[13] ), .o1(new_n160));
  inv000aa1d42x5               g065(.a(\b[12] ), .o1(new_n161));
  nor003aa1n02x5               g066(.a(new_n107), .b(new_n105), .c(new_n103), .o1(new_n162));
  norb02aa1n03x4               g067(.a(new_n102), .b(new_n162), .out0(new_n163));
  nanp02aa1n03x5               g068(.a(new_n119), .b(new_n123), .o1(new_n164));
  aoai13aa1n02x5               g069(.a(new_n155), .b(new_n150), .c(new_n163), .d(new_n164), .o1(new_n165));
  oaoi03aa1n02x5               g070(.a(new_n160), .b(new_n161), .c(new_n165), .o1(new_n166));
  norp02aa1n24x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nanp02aa1n12x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  norb02aa1n06x4               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnrc02aa1n02x5               g074(.a(new_n166), .b(new_n169), .out0(\s[14] ));
  nona23aa1n02x4               g075(.a(new_n156), .b(new_n168), .c(new_n167), .d(new_n157), .out0(new_n171));
  aoai13aa1n02x7               g076(.a(new_n168), .b(new_n167), .c(new_n160), .d(new_n161), .o1(new_n172));
  aoai13aa1n04x5               g077(.a(new_n172), .b(new_n171), .c(new_n152), .d(new_n155), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n03x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nand22aa1n12x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  nor042aa1d18x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand22aa1n04x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  norb02aa1n03x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  aoi112aa1n02x5               g085(.a(new_n180), .b(new_n175), .c(new_n173), .d(new_n177), .o1(new_n181));
  aoai13aa1n03x5               g086(.a(new_n180), .b(new_n175), .c(new_n173), .d(new_n176), .o1(new_n182));
  norb02aa1n02x7               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano23aa1n06x5               g088(.a(new_n178), .b(new_n175), .c(new_n179), .d(new_n176), .out0(new_n184));
  nand23aa1n09x5               g089(.a(new_n184), .b(new_n158), .c(new_n169), .o1(new_n185));
  nor042aa1n06x5               g090(.a(new_n185), .b(new_n150), .o1(new_n186));
  aoai13aa1n12x5               g091(.a(new_n186), .b(new_n108), .c(new_n123), .d(new_n119), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n178), .o1(new_n188));
  aoi112aa1n06x5               g093(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n189));
  inv000aa1n02x5               g094(.a(new_n189), .o1(new_n190));
  nanb03aa1n02x5               g095(.a(new_n172), .b(new_n180), .c(new_n177), .out0(new_n191));
  nand03aa1n02x5               g096(.a(new_n135), .b(new_n134), .c(new_n143), .o1(new_n192));
  tech160nm_fiaoi012aa1n02p5x5 g097(.a(new_n185), .b(new_n192), .c(new_n153), .o1(new_n193));
  nano32aa1n03x7               g098(.a(new_n193), .b(new_n191), .c(new_n190), .d(new_n188), .out0(new_n194));
  nanp02aa1n09x5               g099(.a(new_n194), .b(new_n187), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g101(.a(\a[18] ), .o1(new_n197));
  inv000aa1d42x5               g102(.a(\a[17] ), .o1(new_n198));
  inv000aa1d42x5               g103(.a(\b[16] ), .o1(new_n199));
  oaoi03aa1n03x5               g104(.a(new_n198), .b(new_n199), .c(new_n195), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n197), .out0(\s[18] ));
  xroi22aa1d06x4               g106(.a(new_n198), .b(\b[16] ), .c(new_n197), .d(\b[17] ), .out0(new_n202));
  nanp02aa1n02x5               g107(.a(new_n199), .b(new_n198), .o1(new_n203));
  oaoi03aa1n09x5               g108(.a(\a[18] ), .b(\b[17] ), .c(new_n203), .o1(new_n204));
  nand22aa1n03x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nor042aa1n06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n204), .c(new_n195), .d(new_n202), .o1(new_n208));
  aoi112aa1n02x5               g113(.a(new_n207), .b(new_n204), .c(new_n195), .d(new_n202), .o1(new_n209));
  norb02aa1n02x7               g114(.a(new_n208), .b(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand22aa1n06x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  nona22aa1n02x5               g119(.a(new_n208), .b(new_n214), .c(new_n206), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n214), .o1(new_n216));
  oaoi13aa1n06x5               g121(.a(new_n216), .b(new_n208), .c(\a[19] ), .d(\b[18] ), .o1(new_n217));
  norb02aa1n03x4               g122(.a(new_n215), .b(new_n217), .out0(\s[20] ));
  nano23aa1n06x5               g123(.a(new_n212), .b(new_n206), .c(new_n213), .d(new_n205), .out0(new_n219));
  nanp02aa1n02x5               g124(.a(new_n202), .b(new_n219), .o1(new_n220));
  oai022aa1n03x5               g125(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n221));
  oaib12aa1n09x5               g126(.a(new_n221), .b(new_n197), .c(\b[17] ), .out0(new_n222));
  nona23aa1n09x5               g127(.a(new_n205), .b(new_n213), .c(new_n212), .d(new_n206), .out0(new_n223));
  aoi012aa1n06x5               g128(.a(new_n212), .b(new_n206), .c(new_n213), .o1(new_n224));
  oai012aa1n18x5               g129(.a(new_n224), .b(new_n223), .c(new_n222), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoai13aa1n04x5               g131(.a(new_n226), .b(new_n220), .c(new_n194), .d(new_n187), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  xorc02aa1n02x5               g134(.a(\a[21] ), .b(\b[20] ), .out0(new_n230));
  xorc02aa1n02x5               g135(.a(\a[22] ), .b(\b[21] ), .out0(new_n231));
  aoi112aa1n02x5               g136(.a(new_n229), .b(new_n231), .c(new_n227), .d(new_n230), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n231), .b(new_n229), .c(new_n227), .d(new_n230), .o1(new_n233));
  norb02aa1n02x7               g138(.a(new_n233), .b(new_n232), .out0(\s[22] ));
  inv000aa1d42x5               g139(.a(\a[21] ), .o1(new_n235));
  inv040aa1d32x5               g140(.a(\a[22] ), .o1(new_n236));
  xroi22aa1d06x4               g141(.a(new_n235), .b(\b[20] ), .c(new_n236), .d(\b[21] ), .out0(new_n237));
  nand03aa1n02x5               g142(.a(new_n237), .b(new_n202), .c(new_n219), .o1(new_n238));
  inv000aa1d42x5               g143(.a(\b[21] ), .o1(new_n239));
  oaoi03aa1n12x5               g144(.a(new_n236), .b(new_n239), .c(new_n229), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  tech160nm_fiaoi012aa1n03p5x5 g146(.a(new_n241), .b(new_n225), .c(new_n237), .o1(new_n242));
  aoai13aa1n04x5               g147(.a(new_n242), .b(new_n238), .c(new_n194), .d(new_n187), .o1(new_n243));
  xorb03aa1n02x5               g148(.a(new_n243), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n04x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  and002aa1n12x5               g150(.a(\b[22] ), .b(\a[23] ), .o(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[24] ), .b(\b[23] ), .out0(new_n248));
  aoi112aa1n03x4               g153(.a(new_n245), .b(new_n248), .c(new_n243), .d(new_n247), .o1(new_n249));
  aoai13aa1n03x5               g154(.a(new_n248), .b(new_n245), .c(new_n243), .d(new_n247), .o1(new_n250));
  norb02aa1n02x7               g155(.a(new_n250), .b(new_n249), .out0(\s[24] ));
  nano22aa1n03x7               g156(.a(new_n245), .b(new_n248), .c(new_n247), .out0(new_n252));
  inv030aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  nor002aa1n02x5               g158(.a(new_n238), .b(new_n253), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n224), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n237), .b(new_n255), .c(new_n219), .d(new_n204), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n245), .o1(new_n257));
  oao003aa1n02x5               g162(.a(\a[24] ), .b(\b[23] ), .c(new_n257), .carry(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n253), .c(new_n256), .d(new_n240), .o1(new_n259));
  tech160nm_fixorc02aa1n05x5   g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n259), .c(new_n195), .d(new_n254), .o1(new_n261));
  aoi112aa1n02x5               g166(.a(new_n260), .b(new_n259), .c(new_n195), .d(new_n254), .o1(new_n262));
  norb02aa1n02x7               g167(.a(new_n261), .b(new_n262), .out0(\s[25] ));
  nor042aa1n03x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  tech160nm_fixorc02aa1n04x5   g169(.a(\a[26] ), .b(\b[25] ), .out0(new_n265));
  nona22aa1n02x5               g170(.a(new_n261), .b(new_n265), .c(new_n264), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n264), .o1(new_n267));
  aobi12aa1n06x5               g172(.a(new_n265), .b(new_n261), .c(new_n267), .out0(new_n268));
  norb02aa1n03x4               g173(.a(new_n266), .b(new_n268), .out0(\s[26] ));
  nanp02aa1n06x5               g174(.a(new_n163), .b(new_n164), .o1(new_n270));
  nano22aa1n02x4               g175(.a(new_n172), .b(new_n177), .c(new_n180), .out0(new_n271));
  nanb02aa1n06x5               g176(.a(new_n185), .b(new_n154), .out0(new_n272));
  nona32aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n189), .d(new_n178), .out0(new_n273));
  and002aa1n06x5               g178(.a(new_n265), .b(new_n260), .o(new_n274));
  nano22aa1n03x7               g179(.a(new_n238), .b(new_n252), .c(new_n274), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n273), .c(new_n270), .d(new_n186), .o1(new_n276));
  oao003aa1n02x5               g181(.a(\a[26] ), .b(\b[25] ), .c(new_n267), .carry(new_n277));
  aobi12aa1n06x5               g182(.a(new_n277), .b(new_n259), .c(new_n274), .out0(new_n278));
  nor042aa1n03x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  norb02aa1n02x5               g185(.a(new_n280), .b(new_n279), .out0(new_n281));
  xnbna2aa1n03x5               g186(.a(new_n281), .b(new_n278), .c(new_n276), .out0(\s[27] ));
  inv000aa1n06x5               g187(.a(new_n279), .o1(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[27] ), .b(\a[28] ), .out0(new_n284));
  aobi12aa1n02x7               g189(.a(new_n280), .b(new_n278), .c(new_n276), .out0(new_n285));
  nano22aa1n02x4               g190(.a(new_n285), .b(new_n283), .c(new_n284), .out0(new_n286));
  aobi12aa1n06x5               g191(.a(new_n275), .b(new_n194), .c(new_n187), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n252), .b(new_n241), .c(new_n225), .d(new_n237), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n274), .o1(new_n289));
  aoai13aa1n04x5               g194(.a(new_n277), .b(new_n289), .c(new_n288), .d(new_n258), .o1(new_n290));
  oaih12aa1n02x5               g195(.a(new_n280), .b(new_n290), .c(new_n287), .o1(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n284), .b(new_n291), .c(new_n283), .o1(new_n292));
  nor002aa1n02x5               g197(.a(new_n292), .b(new_n286), .o1(\s[28] ));
  nano22aa1n02x4               g198(.a(new_n284), .b(new_n283), .c(new_n280), .out0(new_n294));
  oaih12aa1n02x5               g199(.a(new_n294), .b(new_n290), .c(new_n287), .o1(new_n295));
  oao003aa1n03x5               g200(.a(\a[28] ), .b(\b[27] ), .c(new_n283), .carry(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[28] ), .b(\a[29] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n295), .c(new_n296), .o1(new_n298));
  aobi12aa1n02x7               g203(.a(new_n294), .b(new_n278), .c(new_n276), .out0(new_n299));
  nano22aa1n02x4               g204(.a(new_n299), .b(new_n296), .c(new_n297), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n298), .b(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g206(.a(new_n110), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g207(.a(new_n281), .b(new_n297), .c(new_n284), .out0(new_n303));
  oaih12aa1n02x5               g208(.a(new_n303), .b(new_n290), .c(new_n287), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .out0(new_n306));
  tech160nm_fiaoi012aa1n02p5x5 g211(.a(new_n306), .b(new_n304), .c(new_n305), .o1(new_n307));
  aobi12aa1n02x7               g212(.a(new_n303), .b(new_n278), .c(new_n276), .out0(new_n308));
  nano22aa1n02x4               g213(.a(new_n308), .b(new_n305), .c(new_n306), .out0(new_n309));
  norp02aa1n03x5               g214(.a(new_n307), .b(new_n309), .o1(\s[30] ));
  xnrc02aa1n02x5               g215(.a(\b[30] ), .b(\a[31] ), .out0(new_n311));
  norb03aa1n02x5               g216(.a(new_n294), .b(new_n306), .c(new_n297), .out0(new_n312));
  aobi12aa1n02x7               g217(.a(new_n312), .b(new_n278), .c(new_n276), .out0(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n314));
  nano22aa1n02x4               g219(.a(new_n313), .b(new_n311), .c(new_n314), .out0(new_n315));
  oaih12aa1n02x5               g220(.a(new_n312), .b(new_n290), .c(new_n287), .o1(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n311), .b(new_n316), .c(new_n314), .o1(new_n317));
  norp02aa1n03x5               g222(.a(new_n317), .b(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g223(.a(new_n112), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g224(.a(\a[3] ), .b(\b[2] ), .c(new_n112), .o1(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g226(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioai012aa1n05x5   g227(.a(new_n121), .b(new_n119), .c(new_n104), .o1(new_n323));
  xnrb03aa1n02x5               g228(.a(new_n323), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g229(.a(new_n103), .o1(new_n325));
  nanb02aa1n02x5               g230(.a(new_n101), .b(new_n106), .out0(new_n326));
  nanb02aa1n02x5               g231(.a(new_n120), .b(new_n323), .out0(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n326), .b(new_n327), .c(new_n325), .out0(\s[7] ));
  aoi013aa1n03x5               g233(.a(new_n101), .b(new_n327), .c(new_n106), .d(new_n325), .o1(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g235(.a(new_n125), .b(new_n163), .c(new_n164), .out0(\s[9] ));
endmodule


