// Benchmark "adder" written by ABC on Wed Jul 17 16:53:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n329, new_n331, new_n333, new_n334,
    new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  nor002aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor022aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n02x4               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  oai012aa1n02x7               g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oaih12aa1n06x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1n12x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor022aa1n06x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  nand22aa1n04x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor042aa1n04x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanb02aa1n06x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  tech160nm_fixorc02aa1n02p5x5 g022(.a(\a[5] ), .b(\b[4] ), .out0(new_n118));
  norb03aa1n09x5               g023(.a(new_n118), .b(new_n114), .c(new_n117), .out0(new_n119));
  inv000aa1d42x5               g024(.a(new_n110), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n111), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n112), .o1(new_n122));
  norp02aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  aoai13aa1n06x5               g028(.a(new_n113), .b(new_n116), .c(new_n123), .d(new_n115), .o1(new_n124));
  aoai13aa1n06x5               g029(.a(new_n120), .b(new_n121), .c(new_n124), .d(new_n122), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoai13aa1n02x5               g031(.a(new_n126), .b(new_n125), .c(new_n119), .d(new_n109), .o1(new_n127));
  xobna2aa1n03x5               g032(.a(new_n97), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  nand42aa1n04x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nor002aa1d32x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanb02aa1n12x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  oai022aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n132));
  nanb02aa1n02x5               g037(.a(new_n132), .b(new_n127), .out0(new_n133));
  aob012aa1n02x5               g038(.a(new_n133), .b(\b[9] ), .c(\a[10] ), .out0(new_n134));
  inv040aa1n04x5               g039(.a(new_n130), .o1(new_n135));
  aoi022aa1d18x5               g040(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n136));
  nand02aa1d16x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  aoi022aa1n02x5               g043(.a(new_n134), .b(new_n131), .c(new_n133), .d(new_n138), .o1(\s[11] ));
  inv020aa1n02x5               g044(.a(new_n102), .o1(new_n140));
  nano23aa1n03x7               g045(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n141));
  aobi12aa1n06x5               g046(.a(new_n108), .b(new_n141), .c(new_n140), .out0(new_n142));
  nanb02aa1n02x5               g047(.a(new_n110), .b(new_n111), .out0(new_n143));
  norb02aa1n02x5               g048(.a(new_n113), .b(new_n112), .out0(new_n144));
  nona23aa1n03x5               g049(.a(new_n118), .b(new_n144), .c(new_n143), .d(new_n117), .out0(new_n145));
  nanp02aa1n02x5               g050(.a(new_n124), .b(new_n122), .o1(new_n146));
  aoi012aa1n02x7               g051(.a(new_n110), .b(new_n146), .c(new_n111), .o1(new_n147));
  tech160nm_fioai012aa1n03p5x5 g052(.a(new_n147), .b(new_n142), .c(new_n145), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n138), .b(new_n132), .c(new_n148), .d(new_n126), .o1(new_n149));
  nor042aa1n02x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand02aa1n06x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  norb02aa1n06x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n149), .c(new_n135), .out0(\s[12] ));
  nona23aa1d24x5               g058(.a(new_n152), .b(new_n126), .c(new_n97), .d(new_n131), .out0(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n125), .c(new_n119), .d(new_n109), .o1(new_n156));
  oaoi03aa1n03x5               g061(.a(\a[12] ), .b(\b[11] ), .c(new_n135), .o1(new_n157));
  nanb03aa1n12x5               g062(.a(new_n150), .b(new_n132), .c(new_n151), .out0(new_n158));
  oabi12aa1n18x5               g063(.a(new_n157), .b(new_n158), .c(new_n137), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(new_n156), .b(new_n160), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanp02aa1n04x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n163), .b(new_n161), .c(new_n164), .o1(new_n165));
  xnrb03aa1n02x5               g070(.a(new_n165), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand22aa1n09x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nona23aa1d18x5               g073(.a(new_n168), .b(new_n164), .c(new_n163), .d(new_n167), .out0(new_n169));
  inv030aa1n02x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n159), .c(new_n148), .d(new_n155), .o1(new_n171));
  aoi012aa1n02x5               g076(.a(new_n167), .b(new_n163), .c(new_n168), .o1(new_n172));
  nor042aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand02aa1n06x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nanb02aa1n06x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  xobna2aa1n03x5               g080(.a(new_n175), .b(new_n171), .c(new_n172), .out0(\s[15] ));
  aoai13aa1n04x5               g081(.a(new_n172), .b(new_n169), .c(new_n156), .d(new_n160), .o1(new_n177));
  nor002aa1n03x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n03x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n173), .c(new_n177), .d(new_n174), .o1(new_n181));
  aoi112aa1n02x5               g086(.a(new_n173), .b(new_n180), .c(new_n177), .d(new_n174), .o1(new_n182));
  nanb02aa1n02x5               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano23aa1n02x5               g088(.a(new_n173), .b(new_n178), .c(new_n179), .d(new_n174), .out0(new_n184));
  nano22aa1n12x5               g089(.a(new_n154), .b(new_n170), .c(new_n184), .out0(new_n185));
  aoai13aa1n12x5               g090(.a(new_n185), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n186));
  norp03aa1n06x5               g091(.a(new_n169), .b(new_n175), .c(new_n180), .o1(new_n187));
  aoai13aa1n02x5               g092(.a(new_n174), .b(new_n167), .c(new_n163), .d(new_n168), .o1(new_n188));
  aboi22aa1n03x5               g093(.a(new_n173), .b(new_n188), .c(\a[16] ), .d(\b[15] ), .out0(new_n189));
  aoi112aa1n09x5               g094(.a(new_n178), .b(new_n189), .c(new_n159), .d(new_n187), .o1(new_n190));
  nor042aa1d18x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  nand42aa1n08x5               g096(.a(\b[16] ), .b(\a[17] ), .o1(new_n192));
  norb02aa1n02x5               g097(.a(new_n192), .b(new_n191), .out0(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n193), .b(new_n186), .c(new_n190), .out0(\s[17] ));
  inv000aa1d42x5               g099(.a(\a[18] ), .o1(new_n195));
  nand02aa1d08x5               g100(.a(new_n186), .b(new_n190), .o1(new_n196));
  tech160nm_fiaoi012aa1n05x5   g101(.a(new_n191), .b(new_n196), .c(new_n193), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[17] ), .c(new_n195), .out0(\s[18] ));
  nanp02aa1n03x5               g103(.a(new_n159), .b(new_n187), .o1(new_n199));
  nona22aa1n03x5               g104(.a(new_n199), .b(new_n189), .c(new_n178), .out0(new_n200));
  nor042aa1d18x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand42aa1n16x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nano23aa1d15x5               g107(.a(new_n191), .b(new_n201), .c(new_n202), .d(new_n192), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n200), .c(new_n148), .d(new_n185), .o1(new_n204));
  oa0012aa1n02x5               g109(.a(new_n202), .b(new_n201), .c(new_n191), .o(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  nor042aa1n09x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nanp02aa1n04x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n09x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n204), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g116(.a(new_n204), .b(new_n206), .o1(new_n212));
  nor042aa1n04x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand22aa1n12x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1n06x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  aoai13aa1n02x5               g120(.a(new_n215), .b(new_n207), .c(new_n212), .d(new_n208), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n209), .b(new_n205), .c(new_n196), .d(new_n203), .o1(new_n217));
  nona22aa1n02x5               g122(.a(new_n217), .b(new_n215), .c(new_n207), .out0(new_n218));
  nanp02aa1n03x5               g123(.a(new_n216), .b(new_n218), .o1(\s[20] ));
  nanb03aa1d18x5               g124(.a(new_n215), .b(new_n203), .c(new_n209), .out0(new_n220));
  nanb03aa1n09x5               g125(.a(new_n213), .b(new_n214), .c(new_n208), .out0(new_n221));
  orn002aa1n02x7               g126(.a(\a[19] ), .b(\b[18] ), .o(new_n222));
  oai112aa1n06x5               g127(.a(new_n222), .b(new_n202), .c(new_n201), .d(new_n191), .o1(new_n223));
  tech160nm_fiaoi012aa1n05x5   g128(.a(new_n213), .b(new_n207), .c(new_n214), .o1(new_n224));
  oai012aa1n12x5               g129(.a(new_n224), .b(new_n223), .c(new_n221), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  aoai13aa1n04x5               g131(.a(new_n226), .b(new_n220), .c(new_n186), .d(new_n190), .o1(new_n227));
  nor042aa1n06x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  nand42aa1n04x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n220), .o1(new_n231));
  aoi112aa1n02x5               g136(.a(new_n230), .b(new_n225), .c(new_n196), .d(new_n231), .o1(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n227), .c(new_n230), .o1(\s[21] ));
  nor042aa1n04x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  nand02aa1n06x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n235), .b(new_n234), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n228), .c(new_n227), .d(new_n230), .o1(new_n238));
  nand42aa1n02x5               g143(.a(new_n227), .b(new_n230), .o1(new_n239));
  nona22aa1n02x4               g144(.a(new_n239), .b(new_n237), .c(new_n228), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[22] ));
  nano23aa1n06x5               g146(.a(new_n228), .b(new_n234), .c(new_n235), .d(new_n229), .out0(new_n242));
  nanb02aa1n02x5               g147(.a(new_n220), .b(new_n242), .out0(new_n243));
  nano22aa1n03x7               g148(.a(new_n213), .b(new_n208), .c(new_n214), .out0(new_n244));
  oaih12aa1n02x5               g149(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .o1(new_n245));
  oab012aa1n03x5               g150(.a(new_n245), .b(new_n191), .c(new_n201), .out0(new_n246));
  inv020aa1n03x5               g151(.a(new_n224), .o1(new_n247));
  aoai13aa1n06x5               g152(.a(new_n242), .b(new_n247), .c(new_n246), .d(new_n244), .o1(new_n248));
  oa0012aa1n02x5               g153(.a(new_n235), .b(new_n234), .c(new_n228), .o(new_n249));
  inv020aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  nanp02aa1n02x5               g155(.a(new_n248), .b(new_n250), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n252), .b(new_n243), .c(new_n186), .d(new_n190), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  tech160nm_fixnrc02aa1n05x5   g161(.a(\b[23] ), .b(\a[24] ), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n255), .c(new_n253), .d(new_n256), .o1(new_n258));
  nand42aa1n02x5               g163(.a(new_n253), .b(new_n256), .o1(new_n259));
  nona22aa1n02x4               g164(.a(new_n259), .b(new_n257), .c(new_n255), .out0(new_n260));
  nanp02aa1n03x5               g165(.a(new_n260), .b(new_n258), .o1(\s[24] ));
  norb02aa1n06x4               g166(.a(new_n256), .b(new_n257), .out0(new_n262));
  nanb03aa1n03x5               g167(.a(new_n220), .b(new_n262), .c(new_n242), .out0(new_n263));
  inv020aa1n04x5               g168(.a(new_n262), .o1(new_n264));
  orn002aa1n02x5               g169(.a(\a[23] ), .b(\b[22] ), .o(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n265), .carry(new_n266));
  aoai13aa1n12x5               g171(.a(new_n266), .b(new_n264), .c(new_n248), .d(new_n250), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n04x5               g173(.a(new_n268), .b(new_n263), .c(new_n186), .d(new_n190), .o1(new_n269));
  xorb03aa1n02x5               g174(.a(new_n269), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  tech160nm_fixnrc02aa1n05x5   g177(.a(\b[25] ), .b(\a[26] ), .out0(new_n273));
  aoai13aa1n03x5               g178(.a(new_n273), .b(new_n271), .c(new_n269), .d(new_n272), .o1(new_n274));
  nand42aa1n02x5               g179(.a(new_n269), .b(new_n272), .o1(new_n275));
  nona22aa1n02x4               g180(.a(new_n275), .b(new_n273), .c(new_n271), .out0(new_n276));
  nanp02aa1n03x5               g181(.a(new_n276), .b(new_n274), .o1(\s[26] ));
  norb02aa1n03x4               g182(.a(new_n272), .b(new_n273), .out0(new_n278));
  inv000aa1n02x5               g183(.a(new_n278), .o1(new_n279));
  nano23aa1d12x5               g184(.a(new_n279), .b(new_n220), .c(new_n262), .d(new_n242), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n200), .c(new_n148), .d(new_n185), .o1(new_n281));
  nanp02aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .o1(new_n282));
  oai022aa1n02x5               g187(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n283));
  aoi022aa1n12x5               g188(.a(new_n267), .b(new_n278), .c(new_n282), .d(new_n283), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n284), .c(new_n281), .out0(\s[27] ));
  nanp02aa1n03x5               g191(.a(new_n284), .b(new_n281), .o1(new_n287));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  xnrc02aa1n12x5               g193(.a(\b[27] ), .b(\a[28] ), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n288), .c(new_n287), .d(new_n285), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n262), .b(new_n249), .c(new_n225), .d(new_n242), .o1(new_n291));
  nanp02aa1n02x5               g196(.a(new_n283), .b(new_n282), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n292), .b(new_n279), .c(new_n291), .d(new_n266), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n285), .b(new_n293), .c(new_n196), .d(new_n280), .o1(new_n294));
  nona22aa1n02x5               g199(.a(new_n294), .b(new_n289), .c(new_n288), .out0(new_n295));
  nanp02aa1n03x5               g200(.a(new_n290), .b(new_n295), .o1(\s[28] ));
  norb02aa1n03x5               g201(.a(new_n285), .b(new_n289), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n293), .c(new_n196), .d(new_n280), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n297), .o1(new_n299));
  orn002aa1n02x5               g204(.a(\a[27] ), .b(\b[26] ), .o(new_n300));
  oao003aa1n03x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n300), .carry(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n299), .c(new_n284), .d(new_n281), .o1(new_n302));
  tech160nm_fixorc02aa1n02p5x5 g207(.a(\a[29] ), .b(\b[28] ), .out0(new_n303));
  norb02aa1n02x5               g208(.a(new_n301), .b(new_n303), .out0(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n298), .d(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g211(.a(new_n289), .b(new_n285), .c(new_n303), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n293), .c(new_n196), .d(new_n280), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n307), .o1(new_n309));
  oaoi03aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .o1(new_n310));
  inv000aa1n03x5               g215(.a(new_n310), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n309), .c(new_n284), .d(new_n281), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .out0(new_n313));
  and002aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .o(new_n314));
  oabi12aa1n02x5               g219(.a(new_n313), .b(\a[29] ), .c(\b[28] ), .out0(new_n315));
  oab012aa1n02x4               g220(.a(new_n315), .b(new_n301), .c(new_n314), .out0(new_n316));
  aoi022aa1n02x7               g221(.a(new_n312), .b(new_n313), .c(new_n308), .d(new_n316), .o1(\s[30] ));
  nand03aa1n02x5               g222(.a(new_n297), .b(new_n303), .c(new_n313), .o1(new_n318));
  nanb02aa1n03x5               g223(.a(new_n318), .b(new_n287), .out0(new_n319));
  xorc02aa1n02x5               g224(.a(\a[31] ), .b(\b[30] ), .out0(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n320), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n321), .b(new_n318), .c(new_n284), .d(new_n281), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n319), .b(new_n322), .c(new_n323), .d(new_n320), .o1(\s[31] ));
  xnrb03aa1n02x5               g229(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  norb02aa1n02x5               g230(.a(new_n104), .b(new_n103), .out0(new_n326));
  aoi112aa1n02x5               g231(.a(new_n105), .b(new_n326), .c(new_n140), .d(new_n106), .o1(new_n327));
  aoib12aa1n02x5               g232(.a(new_n327), .b(new_n109), .c(new_n103), .out0(\s[4] ));
  nanp02aa1n02x5               g233(.a(new_n141), .b(new_n140), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n118), .b(new_n329), .c(new_n108), .out0(\s[5] ));
  oaoi03aa1n02x5               g235(.a(\a[5] ), .b(\b[4] ), .c(new_n142), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g237(.a(new_n144), .b(new_n116), .c(new_n331), .d(new_n115), .o1(new_n333));
  aoi112aa1n02x5               g238(.a(new_n116), .b(new_n144), .c(new_n331), .d(new_n115), .o1(new_n334));
  norb02aa1n02x5               g239(.a(new_n333), .b(new_n334), .out0(\s[7] ));
  xobna2aa1n03x5               g240(.a(new_n143), .b(new_n333), .c(new_n122), .out0(\s[8] ));
  aoi112aa1n02x5               g241(.a(new_n125), .b(new_n126), .c(new_n119), .d(new_n109), .o1(new_n337));
  aoi012aa1n02x5               g242(.a(new_n337), .b(new_n148), .c(new_n126), .o1(\s[9] ));
endmodule


