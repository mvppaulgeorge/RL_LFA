// Benchmark "adder" written by ABC on Wed Jul 17 17:21:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n184, new_n185, new_n186, new_n187, new_n188, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n303,
    new_n306, new_n307, new_n308, new_n310, new_n312;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[4] ), .o1(new_n97));
  inv040aa1d28x5               g002(.a(\b[3] ), .o1(new_n98));
  aoi112aa1n03x5               g003(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n99));
  aoi012aa1n02x7               g004(.a(new_n99), .b(new_n97), .c(new_n98), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  nor002aa1n08x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oai012aa1n12x5               g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  inv000aa1d42x5               g009(.a(\a[3] ), .o1(new_n105));
  obai22aa1d24x5               g010(.a(\b[2] ), .b(new_n105), .c(\b[3] ), .d(\a[4] ), .out0(new_n106));
  oai022aa1n04x7               g011(.a(new_n97), .b(new_n98), .c(\a[3] ), .d(\b[2] ), .o1(new_n107));
  oai013aa1n09x5               g012(.a(new_n100), .b(new_n104), .c(new_n107), .d(new_n106), .o1(new_n108));
  aoi022aa1n06x5               g013(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n109));
  oai122aa1n06x5               g014(.a(new_n109), .b(\a[6] ), .c(\b[5] ), .d(\a[5] ), .e(\b[4] ), .o1(new_n110));
  nanp02aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  orn002aa1n24x5               g016(.a(\a[8] ), .b(\b[7] ), .o(new_n112));
  nand42aa1n10x5               g017(.a(new_n112), .b(new_n111), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\a[6] ), .o1(new_n114));
  obai22aa1d24x5               g019(.a(\b[5] ), .b(new_n114), .c(\b[6] ), .d(\a[7] ), .out0(new_n115));
  nor043aa1d12x5               g020(.a(new_n110), .b(new_n113), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[7] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\b[6] ), .o1(new_n118));
  norp02aa1n02x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  aoai13aa1n04x5               g024(.a(new_n111), .b(new_n119), .c(new_n118), .d(new_n117), .o1(new_n120));
  oaih22aa1d12x5               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  oaib12aa1n06x5               g026(.a(new_n121), .b(new_n118), .c(\a[7] ), .out0(new_n122));
  oai013aa1d12x5               g027(.a(new_n120), .b(new_n122), .c(new_n113), .d(new_n115), .o1(new_n123));
  aoi012aa1n06x5               g028(.a(new_n123), .b(new_n108), .c(new_n116), .o1(new_n124));
  tech160nm_fioaoi03aa1n03p5x5 g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  xorb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n04x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand22aa1n12x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n03x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nanp02aa1n03x5               g034(.a(new_n125), .b(new_n129), .o1(new_n130));
  nor002aa1n03x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  tech160nm_fiaoi012aa1n04x5   g036(.a(new_n127), .b(new_n131), .c(new_n128), .o1(new_n132));
  nand22aa1n06x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n03x4               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n130), .c(new_n132), .out0(\s[11] ));
  nor042aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand02aa1d06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(new_n139));
  inv020aa1n03x5               g044(.a(new_n132), .o1(new_n140));
  nona22aa1n03x5               g045(.a(new_n130), .b(new_n140), .c(new_n134), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n139), .b(new_n141), .c(new_n133), .out0(\s[12] ));
  tech160nm_fixorc02aa1n05x5   g047(.a(\a[9] ), .b(\b[8] ), .out0(new_n143));
  nano32aa1n03x7               g048(.a(new_n139), .b(new_n143), .c(new_n135), .d(new_n129), .out0(new_n144));
  aoai13aa1n03x5               g049(.a(new_n144), .b(new_n123), .c(new_n108), .d(new_n116), .o1(new_n145));
  nano23aa1n06x5               g050(.a(new_n137), .b(new_n134), .c(new_n138), .d(new_n133), .out0(new_n146));
  oa0012aa1n03x5               g051(.a(new_n138), .b(new_n137), .c(new_n134), .o(new_n147));
  aoi012aa1n06x5               g052(.a(new_n147), .b(new_n146), .c(new_n140), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n145), .b(new_n148), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nand42aa1d28x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nor002aa1d32x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  aoi012aa1n02x5               g057(.a(new_n152), .b(new_n149), .c(new_n151), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d24x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nand02aa1d24x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nano23aa1d15x5               g061(.a(new_n155), .b(new_n152), .c(new_n156), .d(new_n151), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoi012aa1n02x5               g063(.a(new_n155), .b(new_n152), .c(new_n156), .o1(new_n159));
  aoai13aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n145), .d(new_n148), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  orn002aa1n02x5               g066(.a(\a[15] ), .b(\b[14] ), .o(new_n162));
  xorc02aa1n12x5               g067(.a(\a[15] ), .b(\b[14] ), .out0(new_n163));
  nanp02aa1n03x5               g068(.a(new_n160), .b(new_n163), .o1(new_n164));
  xorc02aa1n12x5               g069(.a(\a[16] ), .b(\b[15] ), .out0(new_n165));
  xnbna2aa1n03x5               g070(.a(new_n165), .b(new_n164), .c(new_n162), .out0(\s[16] ));
  nand23aa1d12x5               g071(.a(new_n157), .b(new_n163), .c(new_n165), .o1(new_n167));
  nano32aa1d12x5               g072(.a(new_n167), .b(new_n146), .c(new_n143), .d(new_n129), .out0(new_n168));
  oao003aa1n02x5               g073(.a(\a[16] ), .b(\b[15] ), .c(new_n162), .carry(new_n169));
  nanp02aa1n02x5               g074(.a(new_n146), .b(new_n140), .o1(new_n170));
  inv000aa1n02x5               g075(.a(new_n147), .o1(new_n171));
  tech160nm_fiaoi012aa1n04x5   g076(.a(new_n167), .b(new_n170), .c(new_n171), .o1(new_n172));
  nanb03aa1n03x5               g077(.a(new_n159), .b(new_n165), .c(new_n163), .out0(new_n173));
  nano22aa1n06x5               g078(.a(new_n172), .b(new_n173), .c(new_n169), .out0(new_n174));
  oaib12aa1n02x5               g079(.a(new_n174), .b(new_n124), .c(new_n168), .out0(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nand42aa1n04x5               g081(.a(\b[16] ), .b(\a[17] ), .o1(new_n177));
  aoai13aa1n06x5               g082(.a(new_n168), .b(new_n123), .c(new_n108), .d(new_n116), .o1(new_n178));
  oai112aa1n03x5               g083(.a(new_n178), .b(new_n174), .c(\b[16] ), .d(\a[17] ), .o1(new_n179));
  nor042aa1n06x5               g084(.a(\b[17] ), .b(\a[18] ), .o1(new_n180));
  nand22aa1n09x5               g085(.a(\b[17] ), .b(\a[18] ), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  xnbna2aa1n03x5               g087(.a(new_n182), .b(new_n179), .c(new_n177), .out0(\s[18] ));
  nor042aa1d18x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  nano23aa1d15x5               g089(.a(new_n184), .b(new_n180), .c(new_n181), .d(new_n177), .out0(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  aoi012aa1d24x5               g091(.a(new_n180), .b(new_n184), .c(new_n181), .o1(new_n187));
  aoai13aa1n04x5               g092(.a(new_n187), .b(new_n186), .c(new_n178), .d(new_n174), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g094(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand22aa1n04x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nor002aa1d32x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nor002aa1d24x5               g097(.a(\b[19] ), .b(\a[20] ), .o1(new_n193));
  nand02aa1d12x5               g098(.a(\b[19] ), .b(\a[20] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  aoai13aa1n03x5               g100(.a(new_n195), .b(new_n192), .c(new_n188), .d(new_n191), .o1(new_n196));
  aoi112aa1n03x4               g101(.a(new_n195), .b(new_n192), .c(new_n188), .d(new_n191), .o1(new_n197));
  nanb02aa1n03x5               g102(.a(new_n197), .b(new_n196), .out0(\s[20] ));
  nano23aa1n09x5               g103(.a(new_n193), .b(new_n192), .c(new_n194), .d(new_n191), .out0(new_n199));
  nand02aa1n02x5               g104(.a(new_n199), .b(new_n185), .o1(new_n200));
  nona23aa1d18x5               g105(.a(new_n191), .b(new_n194), .c(new_n193), .d(new_n192), .out0(new_n201));
  tech160nm_fioai012aa1n03p5x5 g106(.a(new_n194), .b(new_n193), .c(new_n192), .o1(new_n202));
  oai012aa1n18x5               g107(.a(new_n202), .b(new_n201), .c(new_n187), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n04x5               g109(.a(new_n204), .b(new_n200), .c(new_n178), .d(new_n174), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g111(.a(\b[20] ), .b(\a[21] ), .o1(new_n207));
  xnrc02aa1n12x5               g112(.a(\b[20] ), .b(\a[21] ), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  tech160nm_fixnrc02aa1n05x5   g114(.a(\b[21] ), .b(\a[22] ), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n205), .d(new_n209), .o1(new_n211));
  aoi112aa1n03x4               g116(.a(new_n207), .b(new_n210), .c(new_n205), .d(new_n209), .o1(new_n212));
  nanb02aa1n03x5               g117(.a(new_n212), .b(new_n211), .out0(\s[22] ));
  norp03aa1n06x5               g118(.a(new_n122), .b(new_n113), .c(new_n115), .o1(new_n214));
  norb02aa1n06x4               g119(.a(new_n120), .b(new_n214), .out0(new_n215));
  aob012aa1n06x5               g120(.a(new_n215), .b(new_n108), .c(new_n116), .out0(new_n216));
  oai112aa1n03x5               g121(.a(new_n169), .b(new_n173), .c(new_n148), .d(new_n167), .o1(new_n217));
  norp02aa1n06x5               g122(.a(new_n210), .b(new_n208), .o1(new_n218));
  and003aa1n03x5               g123(.a(new_n218), .b(new_n199), .c(new_n185), .o(new_n219));
  aoai13aa1n06x5               g124(.a(new_n219), .b(new_n217), .c(new_n216), .d(new_n168), .o1(new_n220));
  inv030aa1n02x5               g125(.a(new_n187), .o1(new_n221));
  inv040aa1n02x5               g126(.a(new_n202), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n218), .b(new_n222), .c(new_n199), .d(new_n221), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\a[22] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\b[21] ), .o1(new_n225));
  oao003aa1n02x5               g130(.a(new_n224), .b(new_n225), .c(new_n207), .carry(new_n226));
  inv000aa1n02x5               g131(.a(new_n226), .o1(new_n227));
  nand22aa1n04x5               g132(.a(new_n223), .b(new_n227), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  nor002aa1n04x5               g134(.a(\b[22] ), .b(\a[23] ), .o1(new_n230));
  nand42aa1n03x5               g135(.a(\b[22] ), .b(\a[23] ), .o1(new_n231));
  nanb02aa1n12x5               g136(.a(new_n230), .b(new_n231), .out0(new_n232));
  xobna2aa1n03x5               g137(.a(new_n232), .b(new_n220), .c(new_n229), .out0(\s[23] ));
  xnrc02aa1n02x5               g138(.a(\b[23] ), .b(\a[24] ), .out0(new_n234));
  nona22aa1n03x5               g139(.a(new_n220), .b(new_n228), .c(new_n230), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n234), .b(new_n235), .c(new_n231), .out0(\s[24] ));
  nor002aa1n02x5               g141(.a(new_n234), .b(new_n232), .o1(new_n237));
  nanb03aa1n02x5               g142(.a(new_n200), .b(new_n237), .c(new_n218), .out0(new_n238));
  inv000aa1n02x5               g143(.a(new_n237), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\a[24] ), .o1(new_n240));
  inv000aa1d42x5               g145(.a(\b[23] ), .o1(new_n241));
  oao003aa1n02x5               g146(.a(new_n240), .b(new_n241), .c(new_n230), .carry(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n239), .c(new_n223), .d(new_n227), .o1(new_n244));
  inv040aa1n03x5               g149(.a(new_n244), .o1(new_n245));
  aoai13aa1n04x5               g150(.a(new_n245), .b(new_n238), .c(new_n178), .d(new_n174), .o1(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g152(.a(\b[24] ), .b(\a[25] ), .o1(new_n248));
  xorc02aa1n03x5               g153(.a(\a[25] ), .b(\b[24] ), .out0(new_n249));
  nor002aa1n02x5               g154(.a(\b[25] ), .b(\a[26] ), .o1(new_n250));
  nanp02aa1n02x5               g155(.a(\b[25] ), .b(\a[26] ), .o1(new_n251));
  nanb02aa1n06x5               g156(.a(new_n250), .b(new_n251), .out0(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n248), .c(new_n246), .d(new_n249), .o1(new_n253));
  aoi112aa1n03x4               g158(.a(new_n248), .b(new_n252), .c(new_n246), .d(new_n249), .o1(new_n254));
  nanb02aa1n03x5               g159(.a(new_n254), .b(new_n253), .out0(\s[26] ));
  norb02aa1n09x5               g160(.a(new_n249), .b(new_n252), .out0(new_n256));
  nano32aa1n03x7               g161(.a(new_n200), .b(new_n256), .c(new_n218), .d(new_n237), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n217), .c(new_n216), .d(new_n168), .o1(new_n258));
  oai012aa1n02x5               g163(.a(new_n251), .b(new_n250), .c(new_n248), .o1(new_n259));
  aobi12aa1n06x5               g164(.a(new_n259), .b(new_n244), .c(new_n256), .out0(new_n260));
  norp02aa1n02x5               g165(.a(\b[26] ), .b(\a[27] ), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(\b[26] ), .b(\a[27] ), .o1(new_n262));
  norb02aa1n02x5               g167(.a(new_n262), .b(new_n261), .out0(new_n263));
  xnbna2aa1n03x5               g168(.a(new_n263), .b(new_n260), .c(new_n258), .out0(\s[27] ));
  norp02aa1n02x5               g169(.a(\b[27] ), .b(\a[28] ), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(\b[27] ), .b(\a[28] ), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n266), .b(new_n265), .out0(new_n267));
  oai112aa1n03x5               g172(.a(new_n260), .b(new_n258), .c(\b[26] ), .d(\a[27] ), .o1(new_n268));
  aoi012aa1n02x5               g173(.a(new_n267), .b(new_n268), .c(new_n262), .o1(new_n269));
  aobi12aa1n06x5               g174(.a(new_n257), .b(new_n178), .c(new_n174), .out0(new_n270));
  aoai13aa1n02x7               g175(.a(new_n237), .b(new_n226), .c(new_n203), .d(new_n218), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n256), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n259), .b(new_n272), .c(new_n271), .d(new_n243), .o1(new_n273));
  norp03aa1n03x5               g178(.a(new_n273), .b(new_n270), .c(new_n261), .o1(new_n274));
  nano22aa1n03x7               g179(.a(new_n274), .b(new_n262), .c(new_n267), .out0(new_n275));
  nor002aa1n02x5               g180(.a(new_n269), .b(new_n275), .o1(\s[28] ));
  nano23aa1n02x4               g181(.a(new_n261), .b(new_n265), .c(new_n266), .d(new_n262), .out0(new_n277));
  oaih12aa1n02x5               g182(.a(new_n277), .b(new_n273), .c(new_n270), .o1(new_n278));
  aoi012aa1n02x5               g183(.a(new_n265), .b(new_n261), .c(new_n266), .o1(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[28] ), .b(\a[29] ), .out0(new_n280));
  tech160nm_fiaoi012aa1n03p5x5 g185(.a(new_n280), .b(new_n278), .c(new_n279), .o1(new_n281));
  aobi12aa1n02x7               g186(.a(new_n277), .b(new_n260), .c(new_n258), .out0(new_n282));
  nano22aa1n02x4               g187(.a(new_n282), .b(new_n279), .c(new_n280), .out0(new_n283));
  norp02aa1n03x5               g188(.a(new_n281), .b(new_n283), .o1(\s[29] ));
  xorb03aa1n02x5               g189(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g190(.a(new_n280), .b(new_n263), .c(new_n267), .out0(new_n286));
  oaih12aa1n02x5               g191(.a(new_n286), .b(new_n273), .c(new_n270), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[29] ), .b(\b[28] ), .c(new_n279), .carry(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[29] ), .b(\a[30] ), .out0(new_n289));
  tech160nm_fiaoi012aa1n03p5x5 g194(.a(new_n289), .b(new_n287), .c(new_n288), .o1(new_n290));
  aobi12aa1n02x7               g195(.a(new_n286), .b(new_n260), .c(new_n258), .out0(new_n291));
  nano22aa1n02x4               g196(.a(new_n291), .b(new_n288), .c(new_n289), .out0(new_n292));
  norp02aa1n03x5               g197(.a(new_n290), .b(new_n292), .o1(\s[30] ));
  xnrc02aa1n02x5               g198(.a(\b[30] ), .b(\a[31] ), .out0(new_n294));
  nano23aa1n02x4               g199(.a(new_n289), .b(new_n280), .c(new_n267), .d(new_n263), .out0(new_n295));
  oaih12aa1n02x5               g200(.a(new_n295), .b(new_n273), .c(new_n270), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[30] ), .b(\b[29] ), .c(new_n288), .carry(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n294), .b(new_n296), .c(new_n297), .o1(new_n298));
  aobi12aa1n06x5               g203(.a(new_n295), .b(new_n260), .c(new_n258), .out0(new_n299));
  nano22aa1n02x4               g204(.a(new_n299), .b(new_n294), .c(new_n297), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n298), .b(new_n300), .o1(\s[31] ));
  xorb03aa1n02x5               g206(.a(new_n104), .b(\b[2] ), .c(new_n105), .out0(\s[3] ));
  oaoi03aa1n02x5               g207(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n303));
  xorb03aa1n02x5               g208(.a(new_n303), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g209(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g210(.a(\a[5] ), .o1(new_n306));
  inv000aa1d42x5               g211(.a(\b[4] ), .o1(new_n307));
  oaoi03aa1n02x5               g212(.a(new_n306), .b(new_n307), .c(new_n108), .o1(new_n308));
  xorb03aa1n02x5               g213(.a(new_n308), .b(\b[5] ), .c(new_n114), .out0(\s[6] ));
  oao003aa1n03x5               g214(.a(\a[6] ), .b(\b[5] ), .c(new_n308), .carry(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[6] ), .c(new_n117), .out0(\s[7] ));
  oaoi03aa1n02x5               g216(.a(\a[7] ), .b(\b[6] ), .c(new_n310), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrc02aa1n02x5               g218(.a(new_n124), .b(new_n143), .out0(\s[9] ));
endmodule


