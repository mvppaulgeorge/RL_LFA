// Benchmark "adder" written by ABC on Thu Jul 18 02:02:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n355, new_n357, new_n358, new_n359,
    new_n362, new_n364, new_n366, new_n367, new_n368, new_n370;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  norp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1d28x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nona22aa1n02x4               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  oai012aa1n18x5               g007(.a(new_n100), .b(\b[3] ), .c(\a[4] ), .o1(new_n103));
  and002aa1n24x5               g008(.a(\b[2] ), .b(\a[3] ), .o(new_n104));
  nanp02aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  oai012aa1n02x5               g010(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .o1(new_n106));
  nor003aa1n02x5               g011(.a(new_n106), .b(new_n103), .c(new_n104), .o1(new_n107));
  orn002aa1n02x5               g012(.a(\a[3] ), .b(\b[2] ), .o(new_n108));
  oaoi03aa1n02x5               g013(.a(\a[4] ), .b(\b[3] ), .c(new_n108), .o1(new_n109));
  norp02aa1n12x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor002aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  nor002aa1n03x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand22aa1n02x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  norb02aa1n03x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nor042aa1n09x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  norb02aa1n09x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  nano22aa1n03x5               g025(.a(new_n114), .b(new_n117), .c(new_n120), .out0(new_n121));
  aoai13aa1n06x5               g026(.a(new_n121), .b(new_n109), .c(new_n102), .d(new_n107), .o1(new_n122));
  nano23aa1n06x5               g027(.a(new_n115), .b(new_n118), .c(new_n119), .d(new_n116), .out0(new_n123));
  inv000aa1d42x5               g028(.a(new_n110), .o1(new_n124));
  aob012aa1n02x5               g029(.a(new_n124), .b(new_n112), .c(new_n111), .out0(new_n125));
  inv000aa1d42x5               g030(.a(new_n118), .o1(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[8] ), .b(\b[7] ), .c(new_n126), .o1(new_n127));
  aoi012aa1n12x5               g032(.a(new_n127), .b(new_n123), .c(new_n125), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n98), .b(new_n130), .c(new_n122), .d(new_n128), .o1(new_n131));
  nor022aa1n12x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norb02aa1n09x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  nanp03aa1n02x5               g039(.a(new_n100), .b(\a[1] ), .c(\b[0] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n103), .o1(new_n136));
  nor002aa1n02x5               g041(.a(new_n106), .b(new_n104), .o1(new_n137));
  oai112aa1n04x5               g042(.a(new_n137), .b(new_n136), .c(new_n135), .d(new_n99), .o1(new_n138));
  inv000aa1n02x5               g043(.a(new_n109), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n110), .b(new_n111), .out0(new_n140));
  nanb02aa1n02x5               g045(.a(new_n112), .b(new_n113), .out0(new_n141));
  nona22aa1n09x5               g046(.a(new_n123), .b(new_n141), .c(new_n140), .out0(new_n142));
  aoai13aa1n12x5               g047(.a(new_n128), .b(new_n142), .c(new_n138), .d(new_n139), .o1(new_n143));
  aoi112aa1n02x5               g048(.a(new_n134), .b(new_n97), .c(new_n143), .d(new_n129), .o1(new_n144));
  aoi012aa1n02x5               g049(.a(new_n144), .b(new_n131), .c(new_n134), .o1(\s[10] ));
  inv000aa1d42x5               g050(.a(new_n132), .o1(new_n146));
  aoai13aa1n06x5               g051(.a(new_n134), .b(new_n97), .c(new_n143), .d(new_n129), .o1(new_n147));
  nor002aa1n16x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nanp02aa1n04x5               g053(.a(\b[10] ), .b(\a[11] ), .o1(new_n149));
  norb02aa1n09x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n147), .c(new_n146), .out0(\s[11] ));
  aoai13aa1n02x5               g056(.a(new_n150), .b(new_n132), .c(new_n131), .d(new_n133), .o1(new_n152));
  nor042aa1n04x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  nanp02aa1n04x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  aoib12aa1n02x5               g060(.a(new_n148), .b(new_n154), .c(new_n153), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n148), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n150), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n157), .b(new_n158), .c(new_n147), .d(new_n146), .o1(new_n159));
  aoi022aa1n02x5               g064(.a(new_n159), .b(new_n155), .c(new_n152), .d(new_n156), .o1(\s[12] ));
  nona23aa1d18x5               g065(.a(new_n154), .b(new_n149), .c(new_n148), .d(new_n153), .out0(new_n161));
  nano22aa1n12x5               g066(.a(new_n161), .b(new_n129), .c(new_n134), .out0(new_n162));
  nanp02aa1n02x5               g067(.a(new_n143), .b(new_n162), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n162), .o1(new_n164));
  tech160nm_fiaoi012aa1n05x5   g069(.a(new_n132), .b(new_n97), .c(new_n133), .o1(new_n165));
  tech160nm_fioai012aa1n03p5x5 g070(.a(new_n154), .b(new_n153), .c(new_n148), .o1(new_n166));
  oai012aa1d24x5               g071(.a(new_n166), .b(new_n161), .c(new_n165), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n164), .c(new_n122), .d(new_n128), .o1(new_n169));
  nor002aa1n02x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  nanb03aa1n06x5               g077(.a(new_n165), .b(new_n150), .c(new_n155), .out0(new_n173));
  nano22aa1n02x4               g078(.a(new_n172), .b(new_n173), .c(new_n166), .out0(new_n174));
  aoi022aa1n02x5               g079(.a(new_n169), .b(new_n172), .c(new_n163), .d(new_n174), .o1(\s[13] ));
  orn002aa1n02x5               g080(.a(\a[13] ), .b(\b[12] ), .o(new_n176));
  aoai13aa1n02x5               g081(.a(new_n172), .b(new_n167), .c(new_n143), .d(new_n162), .o1(new_n177));
  nor002aa1n02x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  tech160nm_finand02aa1n03p5x5 g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n177), .c(new_n176), .out0(\s[14] ));
  nano23aa1n02x5               g086(.a(new_n170), .b(new_n178), .c(new_n179), .d(new_n171), .out0(new_n182));
  aoai13aa1n03x5               g087(.a(new_n182), .b(new_n167), .c(new_n143), .d(new_n162), .o1(new_n183));
  aoi012aa1n06x5               g088(.a(new_n178), .b(new_n170), .c(new_n179), .o1(new_n184));
  nor042aa1n06x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nanp02aa1n02x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  norb02aa1n02x5               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n183), .c(new_n184), .out0(\s[15] ));
  inv000aa1n02x5               g093(.a(new_n184), .o1(new_n189));
  aoai13aa1n02x5               g094(.a(new_n187), .b(new_n189), .c(new_n169), .d(new_n182), .o1(new_n190));
  nor042aa1n02x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nand42aa1n02x5               g096(.a(\b[15] ), .b(\a[16] ), .o1(new_n192));
  norb02aa1n02x5               g097(.a(new_n192), .b(new_n191), .out0(new_n193));
  aoib12aa1n02x5               g098(.a(new_n185), .b(new_n192), .c(new_n191), .out0(new_n194));
  inv000aa1d42x5               g099(.a(new_n185), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n187), .o1(new_n196));
  aoai13aa1n03x5               g101(.a(new_n195), .b(new_n196), .c(new_n183), .d(new_n184), .o1(new_n197));
  aoi022aa1n02x5               g102(.a(new_n197), .b(new_n193), .c(new_n190), .d(new_n194), .o1(\s[16] ));
  nona23aa1n06x5               g103(.a(new_n192), .b(new_n186), .c(new_n185), .d(new_n191), .out0(new_n199));
  nano22aa1n03x7               g104(.a(new_n199), .b(new_n172), .c(new_n180), .out0(new_n200));
  nand02aa1d04x5               g105(.a(new_n162), .b(new_n200), .o1(new_n201));
  oai012aa1n02x5               g106(.a(new_n192), .b(new_n191), .c(new_n185), .o1(new_n202));
  tech160nm_fioai012aa1n04x5   g107(.a(new_n202), .b(new_n199), .c(new_n184), .o1(new_n203));
  aoi012aa1n09x5               g108(.a(new_n203), .b(new_n167), .c(new_n200), .o1(new_n204));
  aoai13aa1n12x5               g109(.a(new_n204), .b(new_n201), .c(new_n122), .d(new_n128), .o1(new_n205));
  xorc02aa1n02x5               g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  oai112aa1n02x5               g111(.a(new_n202), .b(new_n206), .c(new_n199), .d(new_n184), .o1(new_n207));
  aoi012aa1n02x5               g112(.a(new_n207), .b(new_n167), .c(new_n200), .o1(new_n208));
  aoai13aa1n02x5               g113(.a(new_n208), .b(new_n201), .c(new_n122), .d(new_n128), .o1(new_n209));
  oaib12aa1n02x5               g114(.a(new_n209), .b(new_n206), .c(new_n205), .out0(\s[17] ));
  inv000aa1d42x5               g115(.a(\a[17] ), .o1(new_n211));
  oaib12aa1n06x5               g116(.a(new_n205), .b(new_n211), .c(\b[16] ), .out0(new_n212));
  oaib12aa1n06x5               g117(.a(new_n212), .b(\b[16] ), .c(new_n211), .out0(new_n213));
  xorc02aa1n02x5               g118(.a(\a[18] ), .b(\b[17] ), .out0(new_n214));
  oabi12aa1n02x5               g119(.a(new_n214), .b(\a[17] ), .c(\b[16] ), .out0(new_n215));
  aboi22aa1n03x5               g120(.a(new_n215), .b(new_n212), .c(new_n213), .d(new_n214), .out0(\s[18] ));
  nano23aa1n02x4               g121(.a(new_n148), .b(new_n153), .c(new_n154), .d(new_n149), .out0(new_n217));
  nano23aa1n02x5               g122(.a(new_n185), .b(new_n191), .c(new_n192), .d(new_n186), .out0(new_n218));
  nanp02aa1n02x5               g123(.a(new_n218), .b(new_n182), .o1(new_n219));
  nano32aa1n06x5               g124(.a(new_n219), .b(new_n217), .c(new_n134), .d(new_n129), .out0(new_n220));
  aobi12aa1n06x5               g125(.a(new_n202), .b(new_n218), .c(new_n189), .out0(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n219), .c(new_n173), .d(new_n166), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\a[18] ), .o1(new_n223));
  xroi22aa1d04x5               g128(.a(new_n211), .b(\b[16] ), .c(new_n223), .d(\b[17] ), .out0(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n222), .c(new_n143), .d(new_n220), .o1(new_n225));
  nor042aa1n02x5               g130(.a(\b[17] ), .b(\a[18] ), .o1(new_n226));
  aoi112aa1n06x5               g131(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n227));
  norp02aa1n09x5               g132(.a(new_n227), .b(new_n226), .o1(new_n228));
  tech160nm_fixorc02aa1n04x5   g133(.a(\a[19] ), .b(\b[18] ), .out0(new_n229));
  xnbna2aa1n03x5               g134(.a(new_n229), .b(new_n225), .c(new_n228), .out0(\s[19] ));
  xnrc02aa1n02x5               g135(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g136(.a(new_n228), .o1(new_n232));
  aoai13aa1n04x5               g137(.a(new_n229), .b(new_n232), .c(new_n205), .d(new_n224), .o1(new_n233));
  xorc02aa1n02x5               g138(.a(\a[20] ), .b(\b[19] ), .out0(new_n234));
  orn002aa1n02x5               g139(.a(\a[19] ), .b(\b[18] ), .o(new_n235));
  norb02aa1n02x5               g140(.a(new_n235), .b(new_n234), .out0(new_n236));
  tech160nm_fixnrc02aa1n04x5   g141(.a(\b[18] ), .b(\a[19] ), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n235), .b(new_n237), .c(new_n225), .d(new_n228), .o1(new_n238));
  aoi022aa1n02x5               g143(.a(new_n238), .b(new_n234), .c(new_n233), .d(new_n236), .o1(\s[20] ));
  tech160nm_fixnrc02aa1n04x5   g144(.a(\b[19] ), .b(\a[20] ), .out0(new_n240));
  nano32aa1n02x4               g145(.a(new_n240), .b(new_n229), .c(new_n214), .d(new_n206), .out0(new_n241));
  aoai13aa1n03x5               g146(.a(new_n241), .b(new_n222), .c(new_n143), .d(new_n220), .o1(new_n242));
  oao003aa1n02x5               g147(.a(\a[20] ), .b(\b[19] ), .c(new_n235), .carry(new_n243));
  oai013aa1d12x5               g148(.a(new_n243), .b(new_n228), .c(new_n237), .d(new_n240), .o1(new_n244));
  nor042aa1n06x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  nand02aa1n03x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  norb02aa1n02x5               g151(.a(new_n246), .b(new_n245), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n244), .c(new_n205), .d(new_n241), .o1(new_n248));
  oai112aa1n04x5               g153(.a(new_n229), .b(new_n234), .c(new_n227), .d(new_n226), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n247), .o1(new_n250));
  and003aa1n02x5               g155(.a(new_n249), .b(new_n250), .c(new_n243), .o(new_n251));
  aobi12aa1n02x7               g156(.a(new_n248), .b(new_n251), .c(new_n242), .out0(\s[21] ));
  nor042aa1n02x5               g157(.a(\b[21] ), .b(\a[22] ), .o1(new_n253));
  nand02aa1n03x5               g158(.a(\b[21] ), .b(\a[22] ), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  aoib12aa1n02x5               g160(.a(new_n245), .b(new_n254), .c(new_n253), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n244), .o1(new_n257));
  inv020aa1n04x5               g162(.a(new_n245), .o1(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n250), .c(new_n242), .d(new_n257), .o1(new_n259));
  aoi022aa1n03x5               g164(.a(new_n259), .b(new_n255), .c(new_n248), .d(new_n256), .o1(\s[22] ));
  nor002aa1n02x5               g165(.a(new_n240), .b(new_n237), .o1(new_n261));
  nano23aa1d15x5               g166(.a(new_n245), .b(new_n253), .c(new_n254), .d(new_n246), .out0(new_n262));
  and003aa1n02x5               g167(.a(new_n224), .b(new_n261), .c(new_n262), .o(new_n263));
  aoai13aa1n02x7               g168(.a(new_n263), .b(new_n222), .c(new_n143), .d(new_n220), .o1(new_n264));
  oaoi03aa1n09x5               g169(.a(\a[22] ), .b(\b[21] ), .c(new_n258), .o1(new_n265));
  aoi012aa1d18x5               g170(.a(new_n265), .b(new_n244), .c(new_n262), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  nor042aa1n09x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .o1(new_n269));
  norb02aa1n02x5               g174(.a(new_n269), .b(new_n268), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n267), .c(new_n205), .d(new_n263), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(new_n270), .b(new_n265), .c(new_n244), .d(new_n262), .o1(new_n272));
  aobi12aa1n02x7               g177(.a(new_n271), .b(new_n272), .c(new_n264), .out0(\s[23] ));
  nor042aa1n02x5               g178(.a(\b[23] ), .b(\a[24] ), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(\b[23] ), .b(\a[24] ), .o1(new_n275));
  norb02aa1n02x5               g180(.a(new_n275), .b(new_n274), .out0(new_n276));
  aoib12aa1n02x5               g181(.a(new_n268), .b(new_n275), .c(new_n274), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n268), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n270), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n278), .b(new_n279), .c(new_n264), .d(new_n266), .o1(new_n280));
  aoi022aa1n03x5               g185(.a(new_n280), .b(new_n276), .c(new_n271), .d(new_n277), .o1(\s[24] ));
  nano23aa1n06x5               g186(.a(new_n268), .b(new_n274), .c(new_n275), .d(new_n269), .out0(new_n282));
  nand22aa1n09x5               g187(.a(new_n282), .b(new_n262), .o1(new_n283));
  nano22aa1n02x4               g188(.a(new_n283), .b(new_n224), .c(new_n261), .out0(new_n284));
  oaoi03aa1n02x5               g189(.a(\a[24] ), .b(\b[23] ), .c(new_n278), .o1(new_n285));
  aoi012aa1n12x5               g190(.a(new_n285), .b(new_n282), .c(new_n265), .o1(new_n286));
  aoai13aa1n12x5               g191(.a(new_n286), .b(new_n283), .c(new_n249), .d(new_n243), .o1(new_n287));
  xorc02aa1n12x5               g192(.a(\a[25] ), .b(\b[24] ), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n287), .c(new_n205), .d(new_n284), .o1(new_n289));
  aoai13aa1n02x7               g194(.a(new_n284), .b(new_n222), .c(new_n143), .d(new_n220), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n283), .o1(new_n291));
  nand02aa1d04x5               g196(.a(new_n244), .b(new_n291), .o1(new_n292));
  aoi112aa1n02x5               g197(.a(new_n285), .b(new_n288), .c(new_n282), .d(new_n265), .o1(new_n293));
  and003aa1n02x5               g198(.a(new_n290), .b(new_n293), .c(new_n292), .o(new_n294));
  norb02aa1n03x4               g199(.a(new_n289), .b(new_n294), .out0(\s[25] ));
  xorc02aa1n02x5               g200(.a(\a[26] ), .b(\b[25] ), .out0(new_n296));
  norp02aa1n02x5               g201(.a(\b[24] ), .b(\a[25] ), .o1(new_n297));
  norp02aa1n02x5               g202(.a(new_n296), .b(new_n297), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n287), .o1(new_n299));
  inv000aa1n02x5               g204(.a(new_n297), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n288), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n300), .b(new_n301), .c(new_n290), .d(new_n299), .o1(new_n302));
  aoi022aa1n02x5               g207(.a(new_n302), .b(new_n296), .c(new_n289), .d(new_n298), .o1(\s[26] ));
  nand02aa1d06x5               g208(.a(new_n296), .b(new_n288), .o1(new_n304));
  nano23aa1n06x5               g209(.a(new_n304), .b(new_n283), .c(new_n224), .d(new_n261), .out0(new_n305));
  aoai13aa1n06x5               g210(.a(new_n305), .b(new_n222), .c(new_n143), .d(new_n220), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n304), .o1(new_n307));
  oaoi03aa1n12x5               g212(.a(\a[26] ), .b(\b[25] ), .c(new_n300), .o1(new_n308));
  aoi012aa1n12x5               g213(.a(new_n308), .b(new_n287), .c(new_n307), .o1(new_n309));
  nor042aa1n03x5               g214(.a(\b[26] ), .b(\a[27] ), .o1(new_n310));
  and002aa1n06x5               g215(.a(\b[26] ), .b(\a[27] ), .o(new_n311));
  nor042aa1n04x5               g216(.a(new_n311), .b(new_n310), .o1(new_n312));
  norb02aa1n02x5               g217(.a(new_n312), .b(new_n308), .out0(new_n313));
  oai112aa1n02x5               g218(.a(new_n306), .b(new_n313), .c(new_n304), .d(new_n299), .o1(new_n314));
  aoai13aa1n02x5               g219(.a(new_n314), .b(new_n312), .c(new_n306), .d(new_n309), .o1(\s[27] ));
  inv000aa1d42x5               g220(.a(new_n308), .o1(new_n316));
  aoai13aa1n06x5               g221(.a(new_n316), .b(new_n304), .c(new_n292), .d(new_n286), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n311), .o1(new_n318));
  aoai13aa1n02x5               g223(.a(new_n318), .b(new_n317), .c(new_n205), .d(new_n305), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n310), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n311), .c(new_n306), .d(new_n309), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[28] ), .b(\b[27] ), .out0(new_n322));
  norp02aa1n02x5               g227(.a(new_n322), .b(new_n310), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n319), .d(new_n323), .o1(\s[28] ));
  and002aa1n12x5               g229(.a(new_n322), .b(new_n312), .o(new_n325));
  aoai13aa1n02x5               g230(.a(new_n325), .b(new_n317), .c(new_n205), .d(new_n305), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n325), .o1(new_n327));
  oaoi03aa1n12x5               g232(.a(\a[28] ), .b(\b[27] ), .c(new_n320), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n328), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n327), .c(new_n306), .d(new_n309), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[29] ), .b(\b[28] ), .out0(new_n331));
  norp02aa1n02x5               g236(.a(new_n328), .b(new_n331), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n326), .d(new_n332), .o1(\s[29] ));
  xorb03aa1n02x5               g238(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g239(.a(new_n322), .b(new_n331), .c(new_n312), .o(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n317), .c(new_n205), .d(new_n305), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n335), .o1(new_n337));
  inv000aa1d42x5               g242(.a(\b[28] ), .o1(new_n338));
  oaib12aa1n02x5               g243(.a(new_n328), .b(new_n338), .c(\a[29] ), .out0(new_n339));
  oa0012aa1n02x5               g244(.a(new_n339), .b(\b[28] ), .c(\a[29] ), .o(new_n340));
  aoai13aa1n03x5               g245(.a(new_n340), .b(new_n337), .c(new_n306), .d(new_n309), .o1(new_n341));
  xorc02aa1n02x5               g246(.a(\a[30] ), .b(\b[29] ), .out0(new_n342));
  oabi12aa1n02x5               g247(.a(new_n342), .b(\a[29] ), .c(\b[28] ), .out0(new_n343));
  norb02aa1n02x5               g248(.a(new_n339), .b(new_n343), .out0(new_n344));
  aoi022aa1n03x5               g249(.a(new_n341), .b(new_n342), .c(new_n336), .d(new_n344), .o1(\s[30] ));
  nanp03aa1n02x5               g250(.a(new_n325), .b(new_n331), .c(new_n342), .o1(new_n346));
  inv000aa1n02x5               g251(.a(new_n346), .o1(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n317), .c(new_n205), .d(new_n305), .o1(new_n348));
  xorc02aa1n02x5               g253(.a(\a[31] ), .b(\b[30] ), .out0(new_n349));
  oai122aa1n02x7               g254(.a(new_n339), .b(\a[30] ), .c(\b[29] ), .d(\a[29] ), .e(\b[28] ), .o1(new_n350));
  aob012aa1n02x5               g255(.a(new_n350), .b(\b[29] ), .c(\a[30] ), .out0(new_n351));
  norb02aa1n02x5               g256(.a(new_n351), .b(new_n349), .out0(new_n352));
  aoai13aa1n03x5               g257(.a(new_n351), .b(new_n346), .c(new_n306), .d(new_n309), .o1(new_n353));
  aoi022aa1n03x5               g258(.a(new_n353), .b(new_n349), .c(new_n348), .d(new_n352), .o1(\s[31] ));
  xorc02aa1n02x5               g259(.a(\a[3] ), .b(\b[2] ), .out0(new_n355));
  xobna2aa1n03x5               g260(.a(new_n355), .b(new_n102), .c(new_n100), .out0(\s[3] ));
  inv000aa1d42x5               g261(.a(new_n104), .o1(new_n357));
  aob012aa1n02x5               g262(.a(new_n355), .b(new_n102), .c(new_n100), .out0(new_n358));
  xnrc02aa1n02x5               g263(.a(\b[3] ), .b(\a[4] ), .out0(new_n359));
  xnbna2aa1n03x5               g264(.a(new_n359), .b(new_n358), .c(new_n357), .out0(\s[4] ));
  xobna2aa1n03x5               g265(.a(new_n141), .b(new_n138), .c(new_n139), .out0(\s[5] ));
  nona22aa1n02x4               g266(.a(new_n138), .b(new_n109), .c(new_n141), .out0(new_n362));
  xnbna2aa1n03x5               g267(.a(new_n140), .b(new_n362), .c(new_n113), .out0(\s[6] ));
  nanb03aa1n02x5               g268(.a(new_n140), .b(new_n362), .c(new_n113), .out0(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n120), .b(new_n364), .c(new_n124), .out0(\s[7] ));
  aob012aa1n02x5               g270(.a(new_n120), .b(new_n364), .c(new_n124), .out0(new_n366));
  nanp02aa1n02x5               g271(.a(new_n366), .b(new_n126), .o1(new_n367));
  aoib12aa1n02x5               g272(.a(new_n118), .b(new_n116), .c(new_n115), .out0(new_n368));
  aoi022aa1n02x5               g273(.a(new_n367), .b(new_n117), .c(new_n366), .d(new_n368), .o1(\s[8] ));
  aoi112aa1n02x5               g274(.a(new_n129), .b(new_n127), .c(new_n123), .d(new_n125), .o1(new_n370));
  aoi022aa1n02x5               g275(.a(new_n143), .b(new_n129), .c(new_n122), .d(new_n370), .o1(\s[9] ));
endmodule


