// Benchmark "adder" written by ABC on Wed Jul 17 15:25:46 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n329, new_n330, new_n331, new_n332, new_n334,
    new_n335, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1d18x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv040aa1n08x5               g003(.a(new_n98), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand42aa1n06x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  tech160nm_fiaoi012aa1n03p5x5 g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor022aa1n06x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  tech160nm_finand02aa1n03p5x5 g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n03x5               g012(.a(new_n104), .b(new_n107), .c(new_n106), .d(new_n105), .out0(new_n108));
  inv000aa1d42x5               g013(.a(\a[3] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  aoai13aa1n02x7               g015(.a(new_n104), .b(new_n105), .c(new_n110), .d(new_n109), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n111), .b(new_n108), .c(new_n103), .o1(new_n112));
  nand42aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n03x7               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  tech160nm_fixorc02aa1n04x5   g022(.a(\a[5] ), .b(\b[4] ), .out0(new_n118));
  norp02aa1n02x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nand42aa1n16x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  norb02aa1n02x5               g025(.a(new_n120), .b(new_n119), .out0(new_n121));
  and003aa1n06x5               g026(.a(new_n117), .b(new_n121), .c(new_n118), .o(new_n122));
  inv000aa1d42x5               g027(.a(\a[8] ), .o1(new_n123));
  oaih22aa1d12x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  aoi022aa1d24x5               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  aoai13aa1n02x5               g030(.a(new_n113), .b(new_n115), .c(new_n124), .d(new_n125), .o1(new_n126));
  oaib12aa1n03x5               g031(.a(new_n126), .b(\b[7] ), .c(new_n123), .out0(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n03x5               g033(.a(new_n128), .b(new_n127), .c(new_n122), .d(new_n112), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g035(.a(new_n97), .o1(new_n131));
  oaoi03aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  aoai13aa1n06x5               g038(.a(new_n133), .b(new_n131), .c(new_n129), .d(new_n99), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n02x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  nor042aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand02aa1n03x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  aoai13aa1n03x5               g046(.a(new_n141), .b(new_n136), .c(new_n134), .d(new_n138), .o1(new_n142));
  nanp02aa1n02x5               g047(.a(new_n134), .b(new_n138), .o1(new_n143));
  nona22aa1n02x4               g048(.a(new_n143), .b(new_n141), .c(new_n136), .out0(new_n144));
  nanp02aa1n02x5               g049(.a(new_n144), .b(new_n142), .o1(\s[12] ));
  nano23aa1n06x5               g050(.a(new_n136), .b(new_n139), .c(new_n140), .d(new_n137), .out0(new_n146));
  and003aa1n02x5               g051(.a(new_n146), .b(new_n128), .c(new_n97), .o(new_n147));
  aoai13aa1n06x5               g052(.a(new_n147), .b(new_n127), .c(new_n122), .d(new_n112), .o1(new_n148));
  oai022aa1n02x5               g053(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n149));
  aoi022aa1n06x5               g054(.a(new_n146), .b(new_n132), .c(new_n140), .d(new_n149), .o1(new_n150));
  nor002aa1n10x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1d28x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n148), .c(new_n150), .out0(\s[13] ));
  nanp02aa1n02x5               g059(.a(new_n148), .b(new_n150), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n151), .b(new_n155), .c(new_n153), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand42aa1n16x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nano23aa1d15x5               g064(.a(new_n151), .b(new_n158), .c(new_n159), .d(new_n152), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n158), .b(new_n151), .c(new_n159), .o1(new_n162));
  aoai13aa1n04x5               g067(.a(new_n162), .b(new_n161), .c(new_n148), .d(new_n150), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanp02aa1n02x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  tech160nm_fixnrc02aa1n03p5x5 g071(.a(\b[15] ), .b(\a[16] ), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n168));
  nanb02aa1n03x5               g073(.a(new_n165), .b(new_n166), .out0(new_n169));
  nanb02aa1n02x5               g074(.a(new_n169), .b(new_n163), .out0(new_n170));
  nona22aa1n02x4               g075(.a(new_n170), .b(new_n167), .c(new_n165), .out0(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n168), .o1(\s[16] ));
  nona22aa1n12x5               g077(.a(new_n160), .b(new_n167), .c(new_n169), .out0(new_n173));
  nano32aa1d12x5               g078(.a(new_n173), .b(new_n146), .c(new_n128), .d(new_n97), .out0(new_n174));
  aoai13aa1n12x5               g079(.a(new_n174), .b(new_n127), .c(new_n122), .d(new_n112), .o1(new_n175));
  nor042aa1n04x5               g080(.a(new_n150), .b(new_n173), .o1(new_n176));
  inv000aa1d42x5               g081(.a(\a[16] ), .o1(new_n177));
  inv000aa1d42x5               g082(.a(\b[15] ), .o1(new_n178));
  aoai13aa1n03x5               g083(.a(new_n166), .b(new_n158), .c(new_n151), .d(new_n159), .o1(new_n179));
  tech160nm_fioai012aa1n03p5x5 g084(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .o1(new_n180));
  tech160nm_fioaoi03aa1n03p5x5 g085(.a(new_n177), .b(new_n178), .c(new_n180), .o1(new_n181));
  norb02aa1d21x5               g086(.a(new_n181), .b(new_n176), .out0(new_n182));
  xorc02aa1n02x5               g087(.a(\a[17] ), .b(\b[16] ), .out0(new_n183));
  xnbna2aa1n03x5               g088(.a(new_n183), .b(new_n175), .c(new_n182), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[18] ), .o1(new_n185));
  nanp02aa1n06x5               g090(.a(new_n175), .b(new_n182), .o1(new_n186));
  nor042aa1n03x5               g091(.a(\b[16] ), .b(\a[17] ), .o1(new_n187));
  tech160nm_fiaoi012aa1n05x5   g092(.a(new_n187), .b(new_n186), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  xroi22aa1d06x4               g095(.a(new_n190), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  aob012aa1n03x5               g097(.a(new_n187), .b(\b[17] ), .c(\a[18] ), .out0(new_n193));
  oaib12aa1n18x5               g098(.a(new_n193), .b(\b[17] ), .c(new_n185), .out0(new_n194));
  inv000aa1d42x5               g099(.a(new_n194), .o1(new_n195));
  aoai13aa1n04x5               g100(.a(new_n195), .b(new_n192), .c(new_n175), .d(new_n182), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanp02aa1n04x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  norb02aa1n09x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  nor042aa1d18x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nand02aa1d28x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  norb02aa1d27x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  aoai13aa1n03x5               g110(.a(new_n205), .b(new_n199), .c(new_n196), .d(new_n201), .o1(new_n206));
  nand02aa1n02x5               g111(.a(new_n196), .b(new_n201), .o1(new_n207));
  nona22aa1n02x5               g112(.a(new_n207), .b(new_n205), .c(new_n199), .out0(new_n208));
  nanp02aa1n03x5               g113(.a(new_n208), .b(new_n206), .o1(\s[20] ));
  nano23aa1n03x7               g114(.a(new_n199), .b(new_n202), .c(new_n203), .d(new_n200), .out0(new_n210));
  nanp02aa1n02x5               g115(.a(new_n191), .b(new_n210), .o1(new_n211));
  tech160nm_fioai012aa1n05x5   g116(.a(new_n203), .b(new_n202), .c(new_n199), .o1(new_n212));
  inv000aa1n02x5               g117(.a(new_n212), .o1(new_n213));
  aoi012aa1n02x5               g118(.a(new_n213), .b(new_n210), .c(new_n194), .o1(new_n214));
  aoai13aa1n04x5               g119(.a(new_n214), .b(new_n211), .c(new_n175), .d(new_n182), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n04x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  tech160nm_fixorc02aa1n04x5   g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[21] ), .b(\a[22] ), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n215), .d(new_n218), .o1(new_n220));
  nand02aa1n02x5               g125(.a(new_n215), .b(new_n218), .o1(new_n221));
  nona22aa1n02x5               g126(.a(new_n221), .b(new_n219), .c(new_n217), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n222), .b(new_n220), .o1(\s[22] ));
  xnrc02aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .out0(new_n224));
  norp02aa1n02x5               g129(.a(new_n219), .b(new_n224), .o1(new_n225));
  nand23aa1n06x5               g130(.a(new_n191), .b(new_n225), .c(new_n210), .o1(new_n226));
  nor042aa1n02x5               g131(.a(\b[17] ), .b(\a[18] ), .o1(new_n227));
  aoi112aa1n09x5               g132(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n228));
  oai112aa1n06x5               g133(.a(new_n201), .b(new_n204), .c(new_n228), .d(new_n227), .o1(new_n229));
  nanb02aa1n03x5               g134(.a(new_n219), .b(new_n218), .out0(new_n230));
  inv000aa1d42x5               g135(.a(\a[22] ), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\b[21] ), .o1(new_n232));
  oaoi03aa1n03x5               g137(.a(new_n231), .b(new_n232), .c(new_n217), .o1(new_n233));
  aoai13aa1n12x5               g138(.a(new_n233), .b(new_n230), .c(new_n229), .d(new_n212), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n226), .c(new_n175), .d(new_n182), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  tech160nm_fixorc02aa1n02p5x5 g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xnrc02aa1n02x5               g144(.a(\b[23] ), .b(\a[24] ), .out0(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n238), .c(new_n236), .d(new_n239), .o1(new_n241));
  nand02aa1n02x5               g146(.a(new_n236), .b(new_n239), .o1(new_n242));
  nona22aa1n02x5               g147(.a(new_n242), .b(new_n240), .c(new_n238), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n243), .b(new_n241), .o1(\s[24] ));
  norb02aa1n02x5               g149(.a(new_n239), .b(new_n240), .out0(new_n245));
  nanb02aa1n02x5               g150(.a(new_n226), .b(new_n245), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n225), .b(new_n213), .c(new_n210), .d(new_n194), .o1(new_n247));
  inv000aa1n02x5               g152(.a(new_n245), .o1(new_n248));
  inv000aa1d42x5               g153(.a(\a[24] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\b[23] ), .o1(new_n250));
  oao003aa1n06x5               g155(.a(new_n249), .b(new_n250), .c(new_n238), .carry(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n248), .c(new_n247), .d(new_n233), .o1(new_n253));
  inv030aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  aoai13aa1n04x5               g159(.a(new_n254), .b(new_n246), .c(new_n175), .d(new_n182), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n02x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  nor002aa1n02x5               g163(.a(\b[25] ), .b(\a[26] ), .o1(new_n259));
  nand42aa1n03x5               g164(.a(\b[25] ), .b(\a[26] ), .o1(new_n260));
  norb02aa1n09x5               g165(.a(new_n260), .b(new_n259), .out0(new_n261));
  inv040aa1n03x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n263));
  nand02aa1n02x5               g168(.a(new_n255), .b(new_n258), .o1(new_n264));
  nona22aa1n02x5               g169(.a(new_n264), .b(new_n262), .c(new_n257), .out0(new_n265));
  nanp02aa1n03x5               g170(.a(new_n265), .b(new_n263), .o1(\s[26] ));
  orn002aa1n02x5               g171(.a(\a[2] ), .b(\b[1] ), .o(new_n267));
  aob012aa1n02x5               g172(.a(new_n267), .b(new_n101), .c(new_n102), .out0(new_n268));
  norb02aa1n02x5               g173(.a(new_n104), .b(new_n105), .out0(new_n269));
  norb02aa1n02x5               g174(.a(new_n107), .b(new_n106), .out0(new_n270));
  nanp03aa1n02x5               g175(.a(new_n268), .b(new_n269), .c(new_n270), .o1(new_n271));
  nanp03aa1n02x5               g176(.a(new_n117), .b(new_n118), .c(new_n121), .o1(new_n272));
  inv000aa1d42x5               g177(.a(\b[7] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n115), .o1(new_n274));
  norp02aa1n02x5               g179(.a(\b[4] ), .b(\a[5] ), .o1(new_n275));
  oai012aa1n02x5               g180(.a(new_n125), .b(new_n119), .c(new_n275), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(new_n276), .b(new_n274), .o1(new_n277));
  oaoi03aa1n02x5               g182(.a(new_n123), .b(new_n273), .c(new_n277), .o1(new_n278));
  aoai13aa1n02x5               g183(.a(new_n278), .b(new_n272), .c(new_n271), .d(new_n111), .o1(new_n279));
  oai012aa1n02x5               g184(.a(new_n181), .b(new_n150), .c(new_n173), .o1(new_n280));
  norb02aa1n02x5               g185(.a(new_n258), .b(new_n262), .out0(new_n281));
  nano22aa1n03x7               g186(.a(new_n226), .b(new_n281), .c(new_n245), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n280), .c(new_n279), .d(new_n174), .o1(new_n283));
  oai012aa1n02x5               g188(.a(new_n260), .b(new_n259), .c(new_n257), .o1(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n253), .c(new_n281), .out0(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n283), .out0(\s[27] ));
  aoai13aa1n04x5               g192(.a(new_n281), .b(new_n251), .c(new_n234), .d(new_n245), .o1(new_n288));
  nand43aa1n02x5               g193(.a(new_n283), .b(new_n288), .c(new_n284), .o1(new_n289));
  norp02aa1n02x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  norp02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .o1(new_n291));
  nanp02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .o1(new_n292));
  nanb02aa1n06x5               g197(.a(new_n291), .b(new_n292), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n289), .d(new_n286), .o1(new_n294));
  aobi12aa1n06x5               g199(.a(new_n282), .b(new_n175), .c(new_n182), .out0(new_n295));
  nand02aa1d04x5               g200(.a(new_n288), .b(new_n284), .o1(new_n296));
  oaih12aa1n02x5               g201(.a(new_n286), .b(new_n296), .c(new_n295), .o1(new_n297));
  nona22aa1n02x5               g202(.a(new_n297), .b(new_n293), .c(new_n290), .out0(new_n298));
  nanp02aa1n03x5               g203(.a(new_n294), .b(new_n298), .o1(\s[28] ));
  norb02aa1n03x5               g204(.a(new_n286), .b(new_n293), .out0(new_n300));
  oaih12aa1n02x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n300), .o1(new_n302));
  aoi012aa1n02x5               g207(.a(new_n291), .b(new_n290), .c(new_n292), .o1(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n302), .c(new_n285), .d(new_n283), .o1(new_n304));
  tech160nm_fixorc02aa1n05x5   g209(.a(\a[29] ), .b(\b[28] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n303), .b(new_n305), .out0(new_n306));
  aoi022aa1n03x5               g211(.a(new_n304), .b(new_n305), .c(new_n301), .d(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g213(.a(new_n293), .b(new_n286), .c(new_n305), .out0(new_n309));
  oaih12aa1n02x5               g214(.a(new_n309), .b(new_n296), .c(new_n295), .o1(new_n310));
  inv000aa1n02x5               g215(.a(new_n309), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n312));
  aoai13aa1n02x7               g217(.a(new_n312), .b(new_n311), .c(new_n285), .d(new_n283), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  norb02aa1n02x5               g219(.a(new_n312), .b(new_n314), .out0(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n310), .d(new_n315), .o1(\s[30] ));
  nanp03aa1n02x5               g221(.a(new_n300), .b(new_n305), .c(new_n314), .o1(new_n317));
  oabi12aa1n03x5               g222(.a(new_n317), .b(new_n296), .c(new_n295), .out0(new_n318));
  xorc02aa1n02x5               g223(.a(\a[31] ), .b(\b[30] ), .out0(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n312), .carry(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(new_n321));
  aoai13aa1n02x7               g226(.a(new_n320), .b(new_n317), .c(new_n285), .d(new_n283), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n322), .b(new_n319), .c(new_n318), .d(new_n321), .o1(\s[31] ));
  xorb03aa1n02x5               g228(.a(new_n103), .b(\b[2] ), .c(new_n109), .out0(\s[3] ));
  aoi112aa1n02x5               g229(.a(new_n106), .b(new_n269), .c(new_n268), .d(new_n107), .o1(new_n325));
  aoib12aa1n02x5               g230(.a(new_n325), .b(new_n112), .c(new_n105), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n112), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g232(.a(new_n275), .b(new_n112), .c(new_n118), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n120), .o1(new_n329));
  norp02aa1n02x5               g234(.a(new_n124), .b(new_n329), .o1(new_n330));
  aobi12aa1n12x5               g235(.a(new_n330), .b(new_n112), .c(new_n118), .out0(new_n331));
  inv000aa1d42x5               g236(.a(new_n331), .o1(new_n332));
  oai012aa1n02x5               g237(.a(new_n332), .b(new_n328), .c(new_n121), .o1(\s[6] ));
  nanb02aa1n02x5               g238(.a(new_n115), .b(new_n116), .out0(new_n334));
  nano32aa1n03x7               g239(.a(new_n331), .b(new_n120), .c(new_n116), .d(new_n274), .out0(new_n335));
  oaoi13aa1n02x5               g240(.a(new_n335), .b(new_n334), .c(new_n329), .d(new_n331), .o1(\s[7] ));
  norp02aa1n02x5               g241(.a(new_n335), .b(new_n115), .o1(new_n337));
  xorb03aa1n02x5               g242(.a(new_n337), .b(\b[7] ), .c(new_n123), .out0(\s[8] ));
  xorb03aa1n02x5               g243(.a(new_n279), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


