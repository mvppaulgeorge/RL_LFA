// Benchmark "adder" written by ABC on Wed Jul 17 23:16:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n316, new_n318, new_n320;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n03x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor042aa1n03x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  norp02aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor022aa1n04x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  tech160nm_finand02aa1n03p5x5 g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nand42aa1n03x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nano23aa1n03x7               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  nor022aa1n04x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nand02aa1d04x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor042aa1n06x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  aoi012aa1n02x5               g014(.a(new_n107), .b(new_n109), .c(new_n108), .o1(new_n110));
  inv020aa1n02x5               g015(.a(new_n110), .o1(new_n111));
  ao0012aa1n03x5               g016(.a(new_n102), .b(new_n104), .c(new_n103), .o(new_n112));
  tech160nm_fiaoi012aa1n03p5x5 g017(.a(new_n112), .b(new_n106), .c(new_n111), .o1(new_n113));
  nor042aa1n04x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nand42aa1n02x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  nor022aa1n04x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  nano23aa1n02x4               g022(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n118));
  and002aa1n02x5               g023(.a(\b[1] ), .b(\a[2] ), .o(new_n119));
  nanp02aa1n02x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  nor002aa1n02x5               g025(.a(\b[1] ), .b(\a[2] ), .o1(new_n121));
  oab012aa1n03x5               g026(.a(new_n119), .b(new_n121), .c(new_n120), .out0(new_n122));
  nanp02aa1n03x5               g027(.a(new_n118), .b(new_n122), .o1(new_n123));
  tech160nm_fiaoi012aa1n04x5   g028(.a(new_n114), .b(new_n116), .c(new_n115), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  nano23aa1n02x4               g030(.a(new_n107), .b(new_n109), .c(new_n125), .d(new_n108), .out0(new_n126));
  nanp02aa1n02x5               g031(.a(new_n126), .b(new_n106), .o1(new_n127));
  aoai13aa1n06x5               g032(.a(new_n113), .b(new_n127), .c(new_n123), .d(new_n124), .o1(new_n128));
  aob012aa1n06x5               g033(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n99), .b(new_n129), .c(new_n101), .out0(\s[10] ));
  aoi013aa1n06x4               g035(.a(new_n98), .b(new_n129), .c(new_n101), .d(new_n99), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1n03x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n06x4               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  nor042aa1n04x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1n10x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n12x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n133), .c(new_n131), .d(new_n135), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(new_n131), .b(new_n135), .o1(new_n141));
  nona22aa1n02x4               g046(.a(new_n141), .b(new_n139), .c(new_n133), .out0(new_n142));
  nanp02aa1n02x5               g047(.a(new_n142), .b(new_n140), .o1(\s[12] ));
  aoi112aa1n02x5               g048(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n144));
  oai112aa1n03x5               g049(.a(new_n138), .b(new_n135), .c(new_n144), .d(new_n97), .o1(new_n145));
  aoi012aa1n02x5               g050(.a(new_n136), .b(new_n133), .c(new_n137), .o1(new_n146));
  and002aa1n02x5               g051(.a(new_n145), .b(new_n146), .o(new_n147));
  nona23aa1n03x5               g052(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n148));
  oabi12aa1n03x5               g053(.a(new_n112), .b(new_n148), .c(new_n110), .out0(new_n149));
  nona23aa1n02x5               g054(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n150));
  oabi12aa1n02x5               g055(.a(new_n119), .b(new_n120), .c(new_n121), .out0(new_n151));
  oaih12aa1n06x5               g056(.a(new_n124), .b(new_n150), .c(new_n151), .o1(new_n152));
  nona23aa1n02x4               g057(.a(new_n125), .b(new_n108), .c(new_n107), .d(new_n109), .out0(new_n153));
  nor042aa1n02x5               g058(.a(new_n153), .b(new_n148), .o1(new_n154));
  xorc02aa1n02x5               g059(.a(\a[9] ), .b(\b[8] ), .out0(new_n155));
  nano32aa1n02x4               g060(.a(new_n139), .b(new_n155), .c(new_n99), .d(new_n135), .out0(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n149), .c(new_n152), .d(new_n154), .o1(new_n157));
  tech160nm_fixorc02aa1n03p5x5 g062(.a(\a[13] ), .b(\b[12] ), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n157), .c(new_n147), .out0(\s[13] ));
  inv000aa1d42x5               g064(.a(\a[14] ), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(new_n157), .b(new_n147), .o1(new_n161));
  nor042aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  aoi012aa1n02x5               g067(.a(new_n162), .b(new_n161), .c(new_n158), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[13] ), .c(new_n160), .out0(\s[14] ));
  xorc02aa1n02x5               g069(.a(\a[14] ), .b(\b[13] ), .out0(new_n165));
  and002aa1n02x5               g070(.a(new_n165), .b(new_n158), .o(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  inv000aa1d42x5               g072(.a(\b[13] ), .o1(new_n168));
  oao003aa1n12x5               g073(.a(new_n160), .b(new_n168), .c(new_n162), .carry(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n167), .c(new_n157), .d(new_n147), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1d28x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nor002aa1n03x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand42aa1n08x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n173), .c(new_n171), .d(new_n174), .o1(new_n178));
  aoi112aa1n02x5               g083(.a(new_n177), .b(new_n173), .c(new_n171), .d(new_n174), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  nano23aa1n06x5               g085(.a(new_n173), .b(new_n175), .c(new_n176), .d(new_n174), .out0(new_n181));
  tech160nm_fiao0012aa1n02p5x5 g086(.a(new_n175), .b(new_n173), .c(new_n176), .o(new_n182));
  tech160nm_fiaoi012aa1n03p5x5 g087(.a(new_n182), .b(new_n181), .c(new_n169), .o1(new_n183));
  nanp03aa1n06x5               g088(.a(new_n181), .b(new_n158), .c(new_n165), .o1(new_n184));
  aoai13aa1n06x5               g089(.a(new_n183), .b(new_n184), .c(new_n146), .d(new_n145), .o1(new_n185));
  inv040aa1n06x5               g090(.a(new_n185), .o1(new_n186));
  nano23aa1n02x4               g091(.a(new_n133), .b(new_n136), .c(new_n137), .d(new_n134), .out0(new_n187));
  nano32aa1n03x7               g092(.a(new_n184), .b(new_n155), .c(new_n187), .d(new_n99), .out0(new_n188));
  aoai13aa1n12x5               g093(.a(new_n188), .b(new_n149), .c(new_n154), .d(new_n152), .o1(new_n189));
  nanp02aa1n06x5               g094(.a(new_n189), .b(new_n186), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g096(.a(\a[18] ), .o1(new_n192));
  inv040aa1d30x5               g097(.a(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[16] ), .o1(new_n194));
  oaoi03aa1n03x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d06x4               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  nor042aa1n02x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  aoi112aa1n09x5               g104(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n200));
  nor002aa1n04x5               g105(.a(new_n200), .b(new_n199), .o1(new_n201));
  aoai13aa1n04x5               g106(.a(new_n201), .b(new_n198), .c(new_n189), .d(new_n186), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n16x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand02aa1d06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nor002aa1d24x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nand42aa1d28x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n15x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n205), .c(new_n202), .d(new_n206), .o1(new_n211));
  norb02aa1n03x5               g116(.a(new_n206), .b(new_n205), .out0(new_n212));
  nand02aa1n02x5               g117(.a(new_n202), .b(new_n212), .o1(new_n213));
  nona22aa1n03x5               g118(.a(new_n213), .b(new_n210), .c(new_n205), .out0(new_n214));
  nanp02aa1n03x5               g119(.a(new_n214), .b(new_n211), .o1(\s[20] ));
  nona23aa1n09x5               g120(.a(new_n208), .b(new_n206), .c(new_n205), .d(new_n207), .out0(new_n216));
  aoi012aa1n06x5               g121(.a(new_n207), .b(new_n205), .c(new_n208), .o1(new_n217));
  oai012aa1n12x5               g122(.a(new_n217), .b(new_n216), .c(new_n201), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  nanb02aa1n06x5               g124(.a(new_n216), .b(new_n197), .out0(new_n220));
  aoai13aa1n04x5               g125(.a(new_n219), .b(new_n220), .c(new_n189), .d(new_n186), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n16x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  xorc02aa1n12x5               g128(.a(\a[21] ), .b(\b[20] ), .out0(new_n224));
  xnrc02aa1n12x5               g129(.a(\b[21] ), .b(\a[22] ), .out0(new_n225));
  aoai13aa1n03x5               g130(.a(new_n225), .b(new_n223), .c(new_n221), .d(new_n224), .o1(new_n226));
  nand02aa1n02x5               g131(.a(new_n221), .b(new_n224), .o1(new_n227));
  nona22aa1n02x5               g132(.a(new_n227), .b(new_n225), .c(new_n223), .out0(new_n228));
  nanp02aa1n03x5               g133(.a(new_n228), .b(new_n226), .o1(\s[22] ));
  oai112aa1n06x5               g134(.a(new_n212), .b(new_n209), .c(new_n200), .d(new_n199), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(new_n225), .b(new_n224), .out0(new_n231));
  inv000aa1d42x5               g136(.a(\a[22] ), .o1(new_n232));
  inv040aa1d28x5               g137(.a(\b[21] ), .o1(new_n233));
  oaoi03aa1n12x5               g138(.a(new_n232), .b(new_n233), .c(new_n223), .o1(new_n234));
  aoai13aa1n12x5               g139(.a(new_n234), .b(new_n231), .c(new_n230), .d(new_n217), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  nona23aa1n08x5               g141(.a(new_n197), .b(new_n224), .c(new_n225), .d(new_n216), .out0(new_n237));
  aoai13aa1n04x5               g142(.a(new_n236), .b(new_n237), .c(new_n189), .d(new_n186), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  xorc02aa1n02x5               g145(.a(\a[23] ), .b(\b[22] ), .out0(new_n241));
  xorc02aa1n12x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n240), .c(new_n238), .d(new_n241), .o1(new_n244));
  nand02aa1n02x5               g149(.a(new_n238), .b(new_n241), .o1(new_n245));
  nona22aa1n02x5               g150(.a(new_n245), .b(new_n243), .c(new_n240), .out0(new_n246));
  nanp02aa1n03x5               g151(.a(new_n246), .b(new_n244), .o1(\s[24] ));
  norb02aa1n02x5               g152(.a(new_n224), .b(new_n225), .out0(new_n248));
  and002aa1n02x5               g153(.a(new_n242), .b(new_n241), .o(new_n249));
  nano22aa1n03x7               g154(.a(new_n220), .b(new_n249), .c(new_n248), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n185), .c(new_n128), .d(new_n188), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n234), .o1(new_n252));
  aoai13aa1n02x7               g157(.a(new_n249), .b(new_n252), .c(new_n218), .d(new_n248), .o1(new_n253));
  inv000aa1d42x5               g158(.a(\a[24] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\b[23] ), .o1(new_n255));
  tech160nm_fioaoi03aa1n03p5x5 g160(.a(new_n254), .b(new_n255), .c(new_n240), .o1(new_n256));
  nanp02aa1n03x5               g161(.a(new_n253), .b(new_n256), .o1(new_n257));
  nanb02aa1n03x5               g162(.a(new_n257), .b(new_n251), .out0(new_n258));
  xorb03aa1n02x5               g163(.a(new_n258), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g164(.a(\b[24] ), .b(\a[25] ), .o1(new_n260));
  xorc02aa1n02x5               g165(.a(\a[25] ), .b(\b[24] ), .out0(new_n261));
  xorc02aa1n12x5               g166(.a(\a[26] ), .b(\b[25] ), .out0(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n03x5               g168(.a(new_n263), .b(new_n260), .c(new_n258), .d(new_n261), .o1(new_n264));
  aoai13aa1n03x5               g169(.a(new_n261), .b(new_n257), .c(new_n190), .d(new_n250), .o1(new_n265));
  nona22aa1n02x5               g170(.a(new_n265), .b(new_n263), .c(new_n260), .out0(new_n266));
  nanp02aa1n03x5               g171(.a(new_n264), .b(new_n266), .o1(\s[26] ));
  inv000aa1d42x5               g172(.a(new_n256), .o1(new_n268));
  and002aa1n06x5               g173(.a(new_n262), .b(new_n261), .o(new_n269));
  aoai13aa1n04x5               g174(.a(new_n269), .b(new_n268), .c(new_n235), .d(new_n249), .o1(new_n270));
  aoi112aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n271));
  oab012aa1n02x4               g176(.a(new_n271), .b(\a[26] ), .c(\b[25] ), .out0(new_n272));
  nano22aa1n03x7               g177(.a(new_n237), .b(new_n249), .c(new_n269), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n185), .c(new_n128), .d(new_n188), .o1(new_n274));
  nand43aa1n03x5               g179(.a(new_n274), .b(new_n270), .c(new_n272), .o1(new_n275));
  xorb03aa1n03x5               g180(.a(new_n275), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[27] ), .b(\a[28] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n269), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n272), .b(new_n281), .c(new_n253), .d(new_n256), .o1(new_n282));
  aobi12aa1n06x5               g187(.a(new_n273), .b(new_n189), .c(new_n186), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n278), .b(new_n282), .c(new_n283), .o1(new_n284));
  nona22aa1n02x5               g189(.a(new_n284), .b(new_n279), .c(new_n277), .out0(new_n285));
  nanp02aa1n03x5               g190(.a(new_n280), .b(new_n285), .o1(\s[28] ));
  norb02aa1n02x5               g191(.a(new_n278), .b(new_n279), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n282), .c(new_n283), .o1(new_n288));
  aob012aa1n03x5               g193(.a(new_n277), .b(\b[27] ), .c(\a[28] ), .out0(new_n289));
  oa0012aa1n12x5               g194(.a(new_n289), .b(\b[27] ), .c(\a[28] ), .o(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[28] ), .b(\a[29] ), .out0(new_n292));
  nona22aa1n02x5               g197(.a(new_n288), .b(new_n291), .c(new_n292), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n292), .b(new_n291), .c(new_n275), .d(new_n287), .o1(new_n294));
  nanp02aa1n03x5               g199(.a(new_n294), .b(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g201(.a(new_n278), .b(new_n292), .c(new_n279), .out0(new_n297));
  oaoi03aa1n09x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .o1(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[29] ), .b(\a[30] ), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n275), .d(new_n297), .o1(new_n300));
  oaih12aa1n02x5               g205(.a(new_n297), .b(new_n282), .c(new_n283), .o1(new_n301));
  nona22aa1n02x5               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  nanp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[30] ));
  nanb02aa1n02x5               g208(.a(new_n299), .b(new_n298), .out0(new_n304));
  oai012aa1n02x5               g209(.a(new_n304), .b(\b[29] ), .c(\a[30] ), .o1(new_n305));
  norb02aa1n02x5               g210(.a(new_n297), .b(new_n299), .out0(new_n306));
  oaih12aa1n02x5               g211(.a(new_n306), .b(new_n282), .c(new_n283), .o1(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  nona22aa1n02x5               g213(.a(new_n307), .b(new_n308), .c(new_n305), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n308), .b(new_n305), .c(new_n275), .d(new_n306), .o1(new_n310));
  nanp02aa1n03x5               g215(.a(new_n310), .b(new_n309), .o1(\s[31] ));
  xorb03aa1n02x5               g216(.a(new_n122), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi012aa1n02x5               g217(.a(new_n116), .b(new_n122), .c(new_n117), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g219(.a(new_n152), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g220(.a(new_n109), .b(new_n152), .c(new_n125), .o1(new_n316));
  xnrb03aa1n02x5               g221(.a(new_n316), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g222(.a(new_n110), .b(new_n153), .c(new_n123), .d(new_n124), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g224(.a(new_n104), .b(new_n318), .c(new_n105), .o1(new_n320));
  xnrb03aa1n02x5               g225(.a(new_n320), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g226(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


