// Benchmark "adder" written by ABC on Thu Jul 18 11:35:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n319,
    new_n321, new_n322, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor002aa1d24x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand42aa1n10x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nand42aa1n10x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nona23aa1n12x5               g007(.a(new_n102), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n103));
  nor002aa1d32x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nand02aa1n16x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  nand02aa1n06x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nona23aa1d24x5               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  nor042aa1n12x5               g013(.a(new_n108), .b(new_n103), .o1(new_n109));
  inv040aa1d32x5               g014(.a(\a[4] ), .o1(new_n110));
  inv000aa1d48x5               g015(.a(\b[3] ), .o1(new_n111));
  nand42aa1n08x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nand42aa1n04x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  nand02aa1n06x5               g018(.a(new_n112), .b(new_n113), .o1(new_n114));
  xnrc02aa1n12x5               g019(.a(\b[2] ), .b(\a[3] ), .out0(new_n115));
  nand42aa1n04x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand02aa1d16x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  nor042aa1n12x5               g022(.a(\b[1] ), .b(\a[2] ), .o1(new_n118));
  oaih12aa1n12x5               g023(.a(new_n116), .b(new_n118), .c(new_n117), .o1(new_n119));
  aoi112aa1n06x5               g024(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n120));
  norb02aa1n09x5               g025(.a(new_n112), .b(new_n120), .out0(new_n121));
  oai013aa1d12x5               g026(.a(new_n121), .b(new_n115), .c(new_n119), .d(new_n114), .o1(new_n122));
  aoi112aa1n02x7               g027(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n123));
  nano23aa1n09x5               g028(.a(new_n99), .b(new_n101), .c(new_n102), .d(new_n100), .out0(new_n124));
  oa0012aa1n12x5               g029(.a(new_n105), .b(new_n106), .c(new_n104), .o(new_n125));
  nanp02aa1n02x5               g030(.a(new_n124), .b(new_n125), .o1(new_n126));
  nona22aa1n02x4               g031(.a(new_n126), .b(new_n123), .c(new_n99), .out0(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n127), .c(new_n109), .d(new_n122), .o1(new_n129));
  nor042aa1n12x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  and002aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .o(new_n131));
  nor042aa1n03x5               g036(.a(new_n131), .b(new_n130), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  inv000aa1n06x5               g038(.a(new_n131), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand22aa1n12x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  nona22aa1n02x4               g042(.a(new_n129), .b(new_n130), .c(new_n97), .out0(new_n138));
  xobna2aa1n03x5               g043(.a(new_n137), .b(new_n138), .c(new_n134), .out0(\s[11] ));
  aoi013aa1n02x4               g044(.a(new_n135), .b(new_n138), .c(new_n137), .d(new_n134), .o1(new_n140));
  xnrb03aa1n03x5               g045(.a(new_n140), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nand02aa1d04x5               g046(.a(new_n122), .b(new_n109), .o1(new_n142));
  aoi112aa1n06x5               g047(.a(new_n123), .b(new_n99), .c(new_n124), .d(new_n125), .o1(new_n143));
  nor002aa1d32x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand22aa1n12x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nano23aa1n06x5               g050(.a(new_n135), .b(new_n144), .c(new_n145), .d(new_n136), .out0(new_n146));
  nanp03aa1n03x5               g051(.a(new_n146), .b(new_n128), .c(new_n132), .o1(new_n147));
  nona23aa1n09x5               g052(.a(new_n145), .b(new_n136), .c(new_n135), .d(new_n144), .out0(new_n148));
  oai012aa1n18x5               g053(.a(new_n134), .b(new_n130), .c(new_n97), .o1(new_n149));
  ao0012aa1n03x7               g054(.a(new_n144), .b(new_n135), .c(new_n145), .o(new_n150));
  oabi12aa1n18x5               g055(.a(new_n150), .b(new_n148), .c(new_n149), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n06x5               g057(.a(new_n152), .b(new_n147), .c(new_n142), .d(new_n143), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g059(.a(\a[14] ), .o1(new_n155));
  nor002aa1n02x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  xnrc02aa1n12x5               g061(.a(\b[12] ), .b(\a[13] ), .out0(new_n157));
  aoib12aa1n02x5               g062(.a(new_n156), .b(new_n153), .c(new_n157), .out0(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(new_n155), .out0(\s[14] ));
  nor042aa1n09x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nanp02aa1n02x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  inv000aa1d42x5               g067(.a(\b[13] ), .o1(new_n163));
  oaoi03aa1n02x5               g068(.a(new_n155), .b(new_n163), .c(new_n156), .o1(new_n164));
  inv000aa1n03x5               g069(.a(new_n164), .o1(new_n165));
  xnrc02aa1n12x5               g070(.a(\b[13] ), .b(\a[14] ), .out0(new_n166));
  nor042aa1n09x5               g071(.a(new_n166), .b(new_n157), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n162), .b(new_n165), .c(new_n153), .d(new_n167), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n165), .b(new_n162), .c(new_n153), .d(new_n167), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(\s[15] ));
  inv030aa1d32x5               g075(.a(new_n160), .o1(new_n171));
  xnrc02aa1n12x5               g076(.a(\b[15] ), .b(\a[16] ), .out0(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n168), .c(new_n171), .out0(\s[16] ));
  nano22aa1n12x5               g079(.a(new_n172), .b(new_n171), .c(new_n161), .out0(new_n175));
  nano22aa1n03x5               g080(.a(new_n147), .b(new_n167), .c(new_n175), .out0(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n127), .c(new_n109), .d(new_n122), .o1(new_n177));
  aoai13aa1n12x5               g082(.a(new_n175), .b(new_n165), .c(new_n151), .d(new_n167), .o1(new_n178));
  oao003aa1n02x5               g083(.a(\a[16] ), .b(\b[15] ), .c(new_n171), .carry(new_n179));
  nanp03aa1d12x5               g084(.a(new_n177), .b(new_n178), .c(new_n179), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g086(.a(\a[18] ), .o1(new_n182));
  inv040aa1n16x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  oaoi03aa1n03x5               g089(.a(new_n183), .b(new_n184), .c(new_n180), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(new_n182), .out0(\s[18] ));
  nano22aa1n03x7               g091(.a(new_n148), .b(new_n128), .c(new_n132), .out0(new_n187));
  nand23aa1n03x5               g092(.a(new_n187), .b(new_n167), .c(new_n175), .o1(new_n188));
  aoi012aa1d18x5               g093(.a(new_n188), .b(new_n142), .c(new_n143), .o1(new_n189));
  inv000aa1n02x5               g094(.a(new_n175), .o1(new_n190));
  oab012aa1n02x5               g095(.a(new_n131), .b(new_n97), .c(new_n130), .out0(new_n191));
  aoai13aa1n03x5               g096(.a(new_n167), .b(new_n150), .c(new_n146), .d(new_n191), .o1(new_n192));
  aoai13aa1n06x5               g097(.a(new_n179), .b(new_n190), .c(new_n192), .d(new_n164), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n183), .b(\b[16] ), .c(new_n182), .d(\b[17] ), .out0(new_n194));
  tech160nm_fioai012aa1n05x5   g099(.a(new_n194), .b(new_n193), .c(new_n189), .o1(new_n195));
  oaih22aa1d12x5               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oaib12aa1n18x5               g101(.a(new_n196), .b(new_n182), .c(\b[17] ), .out0(new_n197));
  nor002aa1d32x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand02aa1d12x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g108(.a(new_n198), .o1(new_n204));
  aoi012aa1n03x5               g109(.a(new_n200), .b(new_n195), .c(new_n197), .o1(new_n205));
  nor002aa1d32x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nand02aa1d28x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nanb02aa1n02x5               g112(.a(new_n206), .b(new_n207), .out0(new_n208));
  nano22aa1n02x4               g113(.a(new_n205), .b(new_n204), .c(new_n208), .out0(new_n209));
  nanp02aa1n02x5               g114(.a(new_n184), .b(new_n183), .o1(new_n210));
  oaoi03aa1n06x5               g115(.a(\a[18] ), .b(\b[17] ), .c(new_n210), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n201), .b(new_n211), .c(new_n180), .d(new_n194), .o1(new_n212));
  aoi012aa1n03x5               g117(.a(new_n208), .b(new_n212), .c(new_n204), .o1(new_n213));
  nor002aa1n02x5               g118(.a(new_n213), .b(new_n209), .o1(\s[20] ));
  nano23aa1n09x5               g119(.a(new_n198), .b(new_n206), .c(new_n207), .d(new_n199), .out0(new_n215));
  nand02aa1d04x5               g120(.a(new_n194), .b(new_n215), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  tech160nm_fioai012aa1n05x5   g122(.a(new_n217), .b(new_n193), .c(new_n189), .o1(new_n218));
  nona23aa1d18x5               g123(.a(new_n207), .b(new_n199), .c(new_n198), .d(new_n206), .out0(new_n219));
  aoi012aa1n12x5               g124(.a(new_n206), .b(new_n198), .c(new_n207), .o1(new_n220));
  oai012aa1d24x5               g125(.a(new_n220), .b(new_n219), .c(new_n197), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  nor002aa1d32x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nand42aa1n03x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n218), .c(new_n222), .out0(\s[21] ));
  inv000aa1d42x5               g131(.a(new_n223), .o1(new_n227));
  aobi12aa1n06x5               g132(.a(new_n225), .b(new_n218), .c(new_n222), .out0(new_n228));
  xnrc02aa1n12x5               g133(.a(\b[21] ), .b(\a[22] ), .out0(new_n229));
  nano22aa1n03x7               g134(.a(new_n228), .b(new_n227), .c(new_n229), .out0(new_n230));
  aoai13aa1n06x5               g135(.a(new_n225), .b(new_n221), .c(new_n180), .d(new_n217), .o1(new_n231));
  tech160nm_fiaoi012aa1n05x5   g136(.a(new_n229), .b(new_n231), .c(new_n227), .o1(new_n232));
  nor002aa1n02x5               g137(.a(new_n232), .b(new_n230), .o1(\s[22] ));
  nano22aa1n09x5               g138(.a(new_n229), .b(new_n227), .c(new_n224), .out0(new_n234));
  and003aa1n02x5               g139(.a(new_n194), .b(new_n234), .c(new_n215), .o(new_n235));
  tech160nm_fioai012aa1n05x5   g140(.a(new_n235), .b(new_n193), .c(new_n189), .o1(new_n236));
  oao003aa1n09x5               g141(.a(\a[22] ), .b(\b[21] ), .c(new_n227), .carry(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(new_n221), .c(new_n234), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[22] ), .b(\a[23] ), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  xnbna2aa1n03x5               g146(.a(new_n241), .b(new_n236), .c(new_n239), .out0(\s[23] ));
  nor042aa1n06x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  tech160nm_fiaoi012aa1n02p5x5 g149(.a(new_n240), .b(new_n236), .c(new_n239), .o1(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[23] ), .b(\a[24] ), .out0(new_n246));
  nano22aa1n03x5               g151(.a(new_n245), .b(new_n244), .c(new_n246), .out0(new_n247));
  inv000aa1n03x5               g152(.a(new_n239), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n241), .b(new_n248), .c(new_n180), .d(new_n235), .o1(new_n249));
  aoi012aa1n03x5               g154(.a(new_n246), .b(new_n249), .c(new_n244), .o1(new_n250));
  nor002aa1n02x5               g155(.a(new_n250), .b(new_n247), .o1(\s[24] ));
  nor042aa1n02x5               g156(.a(new_n246), .b(new_n240), .o1(new_n252));
  nano22aa1n03x7               g157(.a(new_n216), .b(new_n234), .c(new_n252), .out0(new_n253));
  tech160nm_fioai012aa1n05x5   g158(.a(new_n253), .b(new_n193), .c(new_n189), .o1(new_n254));
  inv000aa1n03x5               g159(.a(new_n220), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n234), .b(new_n255), .c(new_n215), .d(new_n211), .o1(new_n256));
  inv030aa1n02x5               g161(.a(new_n252), .o1(new_n257));
  oao003aa1n06x5               g162(.a(\a[24] ), .b(\b[23] ), .c(new_n244), .carry(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n257), .c(new_n256), .d(new_n237), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[24] ), .b(\a[25] ), .out0(new_n260));
  aoib12aa1n06x5               g165(.a(new_n260), .b(new_n254), .c(new_n259), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n260), .o1(new_n262));
  aoi112aa1n02x7               g167(.a(new_n262), .b(new_n259), .c(new_n180), .d(new_n253), .o1(new_n263));
  norp02aa1n03x5               g168(.a(new_n261), .b(new_n263), .o1(\s[25] ));
  nor042aa1n03x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  xnrc02aa1n12x5               g171(.a(\b[25] ), .b(\a[26] ), .out0(new_n267));
  nano22aa1n03x7               g172(.a(new_n261), .b(new_n266), .c(new_n267), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n262), .b(new_n259), .c(new_n180), .d(new_n253), .o1(new_n269));
  aoi012aa1n03x5               g174(.a(new_n267), .b(new_n269), .c(new_n266), .o1(new_n270));
  nor002aa1n02x5               g175(.a(new_n270), .b(new_n268), .o1(\s[26] ));
  nor042aa1n09x5               g176(.a(new_n267), .b(new_n260), .o1(new_n272));
  nano32aa1n09x5               g177(.a(new_n216), .b(new_n272), .c(new_n234), .d(new_n252), .out0(new_n273));
  oai012aa1n09x5               g178(.a(new_n273), .b(new_n193), .c(new_n189), .o1(new_n274));
  oao003aa1n03x5               g179(.a(\a[26] ), .b(\b[25] ), .c(new_n266), .carry(new_n275));
  aobi12aa1n06x5               g180(.a(new_n275), .b(new_n259), .c(new_n272), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n274), .c(new_n276), .out0(\s[27] ));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  inv040aa1n03x5               g184(.a(new_n279), .o1(new_n280));
  aobi12aa1n02x5               g185(.a(new_n277), .b(new_n274), .c(new_n276), .out0(new_n281));
  xnrc02aa1n02x5               g186(.a(\b[27] ), .b(\a[28] ), .out0(new_n282));
  nano22aa1n03x5               g187(.a(new_n281), .b(new_n280), .c(new_n282), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n252), .b(new_n238), .c(new_n221), .d(new_n234), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n272), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n275), .b(new_n285), .c(new_n284), .d(new_n258), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n277), .b(new_n286), .c(new_n180), .d(new_n273), .o1(new_n287));
  aoi012aa1n03x5               g192(.a(new_n282), .b(new_n287), .c(new_n280), .o1(new_n288));
  nor002aa1n02x5               g193(.a(new_n288), .b(new_n283), .o1(\s[28] ));
  norb02aa1n02x5               g194(.a(new_n277), .b(new_n282), .out0(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n286), .c(new_n180), .d(new_n273), .o1(new_n291));
  oao003aa1n02x5               g196(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  aoi012aa1n03x5               g198(.a(new_n293), .b(new_n291), .c(new_n292), .o1(new_n294));
  aobi12aa1n03x5               g199(.a(new_n290), .b(new_n274), .c(new_n276), .out0(new_n295));
  nano22aa1n02x5               g200(.a(new_n295), .b(new_n292), .c(new_n293), .out0(new_n296));
  nor002aa1n02x5               g201(.a(new_n294), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g202(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g203(.a(new_n277), .b(new_n293), .c(new_n282), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n286), .c(new_n180), .d(new_n273), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[29] ), .b(\b[28] ), .c(new_n292), .carry(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[29] ), .b(\a[30] ), .out0(new_n302));
  aoi012aa1n03x5               g207(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n303));
  aobi12aa1n02x5               g208(.a(new_n299), .b(new_n274), .c(new_n276), .out0(new_n304));
  nano22aa1n02x4               g209(.a(new_n304), .b(new_n301), .c(new_n302), .out0(new_n305));
  nor002aa1n02x5               g210(.a(new_n303), .b(new_n305), .o1(\s[30] ));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n299), .b(new_n302), .out0(new_n308));
  aobi12aa1n02x5               g213(.a(new_n308), .b(new_n274), .c(new_n276), .out0(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n301), .carry(new_n310));
  nano22aa1n03x5               g215(.a(new_n309), .b(new_n307), .c(new_n310), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n308), .b(new_n286), .c(new_n180), .d(new_n273), .o1(new_n312));
  aoi012aa1n03x5               g217(.a(new_n307), .b(new_n312), .c(new_n310), .o1(new_n313));
  nor002aa1n02x5               g218(.a(new_n313), .b(new_n311), .o1(\s[31] ));
  xnrb03aa1n02x5               g219(.a(new_n119), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g220(.a(\a[3] ), .b(\b[2] ), .c(new_n119), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g222(.a(new_n122), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g223(.a(new_n106), .b(new_n122), .c(new_n107), .o1(new_n319));
  xnrb03aa1n02x5               g224(.a(new_n319), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g225(.a(new_n108), .o1(new_n321));
  tech160nm_fiao0012aa1n02p5x5 g226(.a(new_n125), .b(new_n122), .c(new_n321), .o(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g228(.a(new_n101), .b(new_n322), .c(new_n102), .o1(new_n324));
  xnrb03aa1n02x5               g229(.a(new_n324), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g230(.a(new_n128), .b(new_n142), .c(new_n143), .out0(\s[9] ));
endmodule


