// Benchmark "adder" written by ABC on Thu Jul 18 15:29:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n151, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[3] ), .b(\a[4] ), .o1(new_n97));
  nanp02aa1n06x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  tech160nm_fiaoi012aa1n03p5x5 g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[1] ), .o1(new_n102));
  nand22aa1n03x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  tech160nm_fioaoi03aa1n04x5   g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n105), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n106));
  oai012aa1n06x5               g011(.a(new_n100), .b(new_n106), .c(new_n104), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor022aa1n04x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nor002aa1n04x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nona23aa1n02x4               g016(.a(new_n108), .b(new_n111), .c(new_n110), .d(new_n109), .out0(new_n112));
  xorc02aa1n12x5               g017(.a(\a[8] ), .b(\b[7] ), .out0(new_n113));
  norp02aa1n24x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanb02aa1n03x5               g020(.a(new_n114), .b(new_n115), .out0(new_n116));
  norb03aa1n03x5               g021(.a(new_n113), .b(new_n112), .c(new_n116), .out0(new_n117));
  nano22aa1n03x7               g022(.a(new_n114), .b(new_n108), .c(new_n115), .out0(new_n118));
  oai022aa1n02x5               g023(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n119));
  nand43aa1n03x5               g024(.a(new_n118), .b(new_n113), .c(new_n119), .o1(new_n120));
  inv000aa1n02x5               g025(.a(new_n114), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[8] ), .b(\b[7] ), .c(new_n121), .o1(new_n122));
  nanb02aa1n03x5               g027(.a(new_n122), .b(new_n120), .out0(new_n123));
  tech160nm_fiaoi012aa1n05x5   g028(.a(new_n123), .b(new_n117), .c(new_n107), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  xorb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand02aa1d08x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nor042aa1n06x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  nand02aa1n03x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nona23aa1n09x5               g035(.a(new_n130), .b(new_n128), .c(new_n127), .d(new_n129), .out0(new_n131));
  oai012aa1d24x5               g036(.a(new_n128), .b(new_n129), .c(new_n127), .o1(new_n132));
  nor002aa1n10x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1n08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  oaoi13aa1n03x5               g040(.a(new_n135), .b(new_n132), .c(new_n124), .d(new_n131), .o1(new_n136));
  oai112aa1n02x5               g041(.a(new_n132), .b(new_n135), .c(new_n124), .d(new_n131), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(\s[11] ));
  norp02aa1n03x5               g043(.a(new_n136), .b(new_n133), .o1(new_n139));
  xnrb03aa1n02x5               g044(.a(new_n139), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norp02aa1n12x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand22aa1n12x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nona23aa1n12x5               g047(.a(new_n142), .b(new_n134), .c(new_n133), .d(new_n141), .out0(new_n143));
  norp02aa1n02x5               g048(.a(new_n143), .b(new_n131), .o1(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n123), .c(new_n107), .d(new_n117), .o1(new_n145));
  ao0012aa1n03x7               g050(.a(new_n141), .b(new_n133), .c(new_n142), .o(new_n146));
  oabi12aa1n18x5               g051(.a(new_n146), .b(new_n143), .c(new_n132), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  xnrc02aa1n12x5               g053(.a(\b[12] ), .b(\a[13] ), .out0(new_n149));
  xobna2aa1n03x5               g054(.a(new_n149), .b(new_n145), .c(new_n148), .out0(\s[13] ));
  orn002aa1n24x5               g055(.a(\a[13] ), .b(\b[12] ), .o(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n149), .c(new_n145), .d(new_n148), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nanp02aa1n04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nanb02aa1n06x5               g060(.a(new_n154), .b(new_n155), .out0(new_n156));
  nor042aa1n09x5               g061(.a(new_n149), .b(new_n156), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  oaoi03aa1n09x5               g063(.a(\a[14] ), .b(\b[13] ), .c(new_n151), .o1(new_n159));
  inv000aa1n02x5               g064(.a(new_n159), .o1(new_n160));
  aoai13aa1n04x5               g065(.a(new_n160), .b(new_n158), .c(new_n145), .d(new_n148), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nand42aa1d28x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nor042aa1n04x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nand42aa1n16x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n163), .c(new_n161), .d(new_n164), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n163), .b(new_n168), .c(new_n161), .d(new_n164), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nano23aa1n02x4               g076(.a(new_n127), .b(new_n129), .c(new_n130), .d(new_n128), .out0(new_n172));
  nano23aa1n02x5               g077(.a(new_n133), .b(new_n141), .c(new_n142), .d(new_n134), .out0(new_n173));
  nano23aa1d15x5               g078(.a(new_n163), .b(new_n165), .c(new_n166), .d(new_n164), .out0(new_n174));
  nano32aa1n03x7               g079(.a(new_n158), .b(new_n174), .c(new_n172), .d(new_n173), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n123), .c(new_n107), .d(new_n117), .o1(new_n176));
  aoai13aa1n12x5               g081(.a(new_n174), .b(new_n159), .c(new_n147), .d(new_n157), .o1(new_n177));
  aoi012aa1n02x5               g082(.a(new_n165), .b(new_n163), .c(new_n166), .o1(new_n178));
  nanp03aa1d12x5               g083(.a(new_n176), .b(new_n177), .c(new_n178), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  tech160nm_fioaoi03aa1n03p5x5 g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  oao003aa1n02x5               g090(.a(new_n101), .b(new_n102), .c(new_n103), .carry(new_n186));
  nano23aa1n02x4               g091(.a(new_n97), .b(new_n99), .c(new_n105), .d(new_n98), .out0(new_n187));
  aobi12aa1n03x5               g092(.a(new_n100), .b(new_n187), .c(new_n186), .out0(new_n188));
  nanb02aa1n02x5               g093(.a(new_n109), .b(new_n108), .out0(new_n189));
  norb02aa1n02x5               g094(.a(new_n111), .b(new_n110), .out0(new_n190));
  nona23aa1n09x5               g095(.a(new_n190), .b(new_n113), .c(new_n189), .d(new_n116), .out0(new_n191));
  aoi013aa1n02x4               g096(.a(new_n122), .b(new_n118), .c(new_n113), .d(new_n119), .o1(new_n192));
  nona23aa1n09x5               g097(.a(new_n157), .b(new_n174), .c(new_n143), .d(new_n131), .out0(new_n193));
  oaoi13aa1n09x5               g098(.a(new_n193), .b(new_n192), .c(new_n188), .d(new_n191), .o1(new_n194));
  inv000aa1d42x5               g099(.a(new_n174), .o1(new_n195));
  inv030aa1n04x5               g100(.a(new_n132), .o1(new_n196));
  aoai13aa1n03x5               g101(.a(new_n157), .b(new_n146), .c(new_n173), .d(new_n196), .o1(new_n197));
  aoai13aa1n06x5               g102(.a(new_n178), .b(new_n195), .c(new_n197), .d(new_n160), .o1(new_n198));
  xroi22aa1d06x4               g103(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n199));
  oaih12aa1n02x5               g104(.a(new_n199), .b(new_n198), .c(new_n194), .o1(new_n200));
  oaih22aa1n04x5               g105(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n201));
  oaib12aa1n09x5               g106(.a(new_n201), .b(new_n181), .c(\b[17] ), .out0(new_n202));
  nor002aa1n20x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand02aa1n06x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n200), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g113(.a(new_n203), .o1(new_n209));
  nanp02aa1n02x5               g114(.a(new_n183), .b(new_n182), .o1(new_n210));
  oaoi03aa1n02x5               g115(.a(\a[18] ), .b(\b[17] ), .c(new_n210), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n206), .b(new_n211), .c(new_n179), .d(new_n199), .o1(new_n212));
  nor002aa1n06x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d06x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  aoi012aa1n03x5               g120(.a(new_n215), .b(new_n212), .c(new_n209), .o1(new_n216));
  tech160nm_fiaoi012aa1n02p5x5 g121(.a(new_n205), .b(new_n200), .c(new_n202), .o1(new_n217));
  nano22aa1n03x5               g122(.a(new_n217), .b(new_n209), .c(new_n215), .out0(new_n218));
  norp02aa1n03x5               g123(.a(new_n216), .b(new_n218), .o1(\s[20] ));
  nano23aa1n09x5               g124(.a(new_n203), .b(new_n213), .c(new_n214), .d(new_n204), .out0(new_n220));
  nand02aa1n04x5               g125(.a(new_n199), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  oaih12aa1n02x5               g127(.a(new_n222), .b(new_n198), .c(new_n194), .o1(new_n223));
  nona23aa1d18x5               g128(.a(new_n214), .b(new_n204), .c(new_n203), .d(new_n213), .out0(new_n224));
  aoi012aa1n12x5               g129(.a(new_n213), .b(new_n203), .c(new_n214), .o1(new_n225));
  oai012aa1d24x5               g130(.a(new_n225), .b(new_n224), .c(new_n202), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nor042aa1n09x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  xnbna2aa1n03x5               g135(.a(new_n230), .b(new_n223), .c(new_n227), .out0(\s[21] ));
  inv000aa1d42x5               g136(.a(new_n228), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n230), .b(new_n226), .c(new_n179), .d(new_n222), .o1(new_n233));
  tech160nm_fixnrc02aa1n04x5   g138(.a(\b[21] ), .b(\a[22] ), .out0(new_n234));
  aoi012aa1n03x5               g139(.a(new_n234), .b(new_n233), .c(new_n232), .o1(new_n235));
  aobi12aa1n02x7               g140(.a(new_n230), .b(new_n223), .c(new_n227), .out0(new_n236));
  nano22aa1n02x4               g141(.a(new_n236), .b(new_n232), .c(new_n234), .out0(new_n237));
  norp02aa1n03x5               g142(.a(new_n235), .b(new_n237), .o1(\s[22] ));
  nano22aa1n03x7               g143(.a(new_n234), .b(new_n232), .c(new_n229), .out0(new_n239));
  and003aa1n02x5               g144(.a(new_n199), .b(new_n239), .c(new_n220), .o(new_n240));
  oaih12aa1n02x5               g145(.a(new_n240), .b(new_n198), .c(new_n194), .o1(new_n241));
  oao003aa1n02x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n232), .carry(new_n242));
  inv000aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n243), .b(new_n226), .c(new_n239), .o1(new_n244));
  xnrc02aa1n12x5               g149(.a(\b[22] ), .b(\a[23] ), .out0(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xnbna2aa1n03x5               g151(.a(new_n246), .b(new_n241), .c(new_n244), .out0(\s[23] ));
  nor042aa1n03x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  inv030aa1n02x5               g154(.a(new_n244), .o1(new_n250));
  aoai13aa1n04x5               g155(.a(new_n246), .b(new_n250), .c(new_n179), .d(new_n240), .o1(new_n251));
  xnrc02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .out0(new_n252));
  aoi012aa1n03x5               g157(.a(new_n252), .b(new_n251), .c(new_n249), .o1(new_n253));
  tech160nm_fiaoi012aa1n03p5x5 g158(.a(new_n245), .b(new_n241), .c(new_n244), .o1(new_n254));
  nano22aa1n03x7               g159(.a(new_n254), .b(new_n249), .c(new_n252), .out0(new_n255));
  nor002aa1n02x5               g160(.a(new_n253), .b(new_n255), .o1(\s[24] ));
  nor042aa1n03x5               g161(.a(new_n252), .b(new_n245), .o1(new_n257));
  nano22aa1n03x7               g162(.a(new_n221), .b(new_n239), .c(new_n257), .out0(new_n258));
  oaih12aa1n02x5               g163(.a(new_n258), .b(new_n198), .c(new_n194), .o1(new_n259));
  inv020aa1n04x5               g164(.a(new_n225), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n239), .b(new_n260), .c(new_n220), .d(new_n211), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n257), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .carry(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n261), .d(new_n242), .o1(new_n264));
  xnrc02aa1n12x5               g169(.a(\b[24] ), .b(\a[25] ), .out0(new_n265));
  aoib12aa1n06x5               g170(.a(new_n265), .b(new_n259), .c(new_n264), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n265), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n267), .b(new_n264), .c(new_n179), .d(new_n258), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n266), .b(new_n268), .o1(\s[25] ));
  nor042aa1n03x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoai13aa1n04x5               g176(.a(new_n267), .b(new_n264), .c(new_n179), .d(new_n258), .o1(new_n272));
  xnrc02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .out0(new_n273));
  aoi012aa1n03x5               g178(.a(new_n273), .b(new_n272), .c(new_n271), .o1(new_n274));
  nano22aa1n03x5               g179(.a(new_n266), .b(new_n271), .c(new_n273), .out0(new_n275));
  nor002aa1n02x5               g180(.a(new_n274), .b(new_n275), .o1(\s[26] ));
  nor042aa1n06x5               g181(.a(new_n273), .b(new_n265), .o1(new_n277));
  nano32aa1d12x5               g182(.a(new_n221), .b(new_n277), .c(new_n239), .d(new_n257), .out0(new_n278));
  oai012aa1n06x5               g183(.a(new_n278), .b(new_n198), .c(new_n194), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n280));
  aobi12aa1n06x5               g185(.a(new_n280), .b(new_n264), .c(new_n277), .out0(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n279), .c(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n257), .b(new_n243), .c(new_n226), .d(new_n239), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n277), .o1(new_n287));
  aoai13aa1n12x5               g192(.a(new_n280), .b(new_n287), .c(new_n286), .d(new_n263), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n282), .b(new_n288), .c(new_n179), .d(new_n278), .o1(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[27] ), .b(\a[28] ), .out0(new_n290));
  aoi012aa1n03x5               g195(.a(new_n290), .b(new_n289), .c(new_n285), .o1(new_n291));
  aobi12aa1n03x5               g196(.a(new_n282), .b(new_n279), .c(new_n281), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n285), .c(new_n290), .out0(new_n293));
  nor002aa1n02x5               g198(.a(new_n291), .b(new_n293), .o1(\s[28] ));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  norb02aa1n02x5               g200(.a(new_n282), .b(new_n290), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n288), .c(new_n179), .d(new_n278), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n298));
  aoi012aa1n03x5               g203(.a(new_n295), .b(new_n297), .c(new_n298), .o1(new_n299));
  aobi12aa1n02x7               g204(.a(new_n296), .b(new_n279), .c(new_n281), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n295), .c(new_n298), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g208(.a(\b[29] ), .b(\a[30] ), .out0(new_n304));
  norb03aa1n02x5               g209(.a(new_n282), .b(new_n295), .c(new_n290), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n288), .c(new_n179), .d(new_n278), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n307));
  aoi012aa1n03x5               g212(.a(new_n304), .b(new_n306), .c(new_n307), .o1(new_n308));
  aobi12aa1n02x7               g213(.a(new_n305), .b(new_n279), .c(new_n281), .out0(new_n309));
  nano22aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n307), .out0(new_n310));
  norp02aa1n03x5               g215(.a(new_n308), .b(new_n310), .o1(\s[30] ));
  norb02aa1n02x5               g216(.a(new_n305), .b(new_n304), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n288), .c(new_n179), .d(new_n278), .o1(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  aoi012aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n314), .o1(new_n316));
  aobi12aa1n02x7               g221(.a(new_n312), .b(new_n279), .c(new_n281), .out0(new_n317));
  nano22aa1n03x5               g222(.a(new_n317), .b(new_n314), .c(new_n315), .out0(new_n318));
  norp02aa1n03x5               g223(.a(new_n316), .b(new_n318), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g228(.a(new_n111), .b(new_n107), .c(new_n110), .o1(new_n324));
  xnrb03aa1n02x5               g229(.a(new_n324), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g230(.a(new_n189), .b(new_n324), .out0(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n116), .b(new_n326), .c(new_n108), .out0(\s[7] ));
  nanp02aa1n02x5               g232(.a(new_n326), .b(new_n118), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n113), .b(new_n328), .c(new_n121), .out0(\s[8] ));
  xnrb03aa1n02x5               g234(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


