// Benchmark "adder" written by ABC on Wed Jul 10 16:57:14 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n316, new_n318, new_n320;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  160nm_ficinv00aa1n08x5       g002(.clk(new_n97), .clkout(new_n98));
  and002aa1n02x5               g003(.a(\b[8] ), .b(\a[9] ), .o(new_n99));
  160nm_ficinv00aa1n08x5       g004(.clk(new_n99), .clkout(new_n100));
  and002aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o(new_n101));
  xnrc02aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .out0(new_n102));
  aoi022aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n103));
  oab012aa1n02x4               g008(.a(new_n103), .b(\a[2] ), .c(\b[1] ), .out0(new_n104));
  oa0022aa1n02x5               g009(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n105));
  oaoi13aa1n02x5               g010(.a(new_n101), .b(new_n105), .c(new_n104), .d(new_n102), .o1(new_n106));
  norp02aa1n02x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nona23aa1n02x4               g015(.a(new_n110), .b(new_n108), .c(new_n107), .d(new_n109), .out0(new_n111));
  xorc02aa1n02x5               g016(.a(\a[6] ), .b(\b[5] ), .out0(new_n112));
  xorc02aa1n02x5               g017(.a(\a[5] ), .b(\b[4] ), .out0(new_n113));
  nano22aa1n02x4               g018(.a(new_n111), .b(new_n112), .c(new_n113), .out0(new_n114));
  nanp02aa1n02x5               g019(.a(new_n106), .b(new_n114), .o1(new_n115));
  aoi112aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n116));
  nano23aa1n02x4               g021(.a(new_n107), .b(new_n109), .c(new_n110), .d(new_n108), .out0(new_n117));
  and002aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o(new_n118));
  160nm_ficinv00aa1n08x5       g023(.clk(\a[5] ), .clkout(new_n119));
  160nm_ficinv00aa1n08x5       g024(.clk(\a[6] ), .clkout(new_n120));
  160nm_ficinv00aa1n08x5       g025(.clk(\b[4] ), .clkout(new_n121));
  aboi22aa1n03x5               g026(.a(\b[5] ), .b(new_n120), .c(new_n119), .d(new_n121), .out0(new_n122));
  nona22aa1n02x4               g027(.a(new_n117), .b(new_n118), .c(new_n122), .out0(new_n123));
  nona22aa1n02x4               g028(.a(new_n123), .b(new_n116), .c(new_n107), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  nona22aa1n02x4               g030(.a(new_n115), .b(new_n124), .c(new_n125), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n98), .b(new_n126), .c(new_n100), .out0(\s[10] ));
  nanp02aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  aob012aa1n02x5               g033(.a(new_n97), .b(new_n126), .c(new_n100), .out0(new_n129));
  norp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xobna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n128), .out0(\s[11] ));
  160nm_ficinv00aa1n08x5       g038(.clk(new_n130), .clkout(new_n134));
  nano22aa1n02x4               g039(.a(new_n130), .b(new_n128), .c(new_n131), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n98), .c(new_n126), .d(new_n100), .o1(new_n136));
  xorc02aa1n02x5               g041(.a(\a[12] ), .b(\b[11] ), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n136), .c(new_n134), .out0(\s[12] ));
  xorc02aa1n02x5               g043(.a(\a[13] ), .b(\b[12] ), .out0(new_n139));
  oai022aa1n02x5               g044(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n140));
  nona23aa1n02x4               g045(.a(new_n135), .b(new_n137), .c(new_n140), .d(new_n99), .out0(new_n141));
  160nm_ficinv00aa1n08x5       g046(.clk(new_n141), .clkout(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n124), .c(new_n106), .d(new_n114), .o1(new_n143));
  norp02aa1n02x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  aoi112aa1n02x5               g049(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n145));
  aoi113aa1n02x5               g050(.a(new_n145), .b(new_n144), .c(new_n135), .d(new_n137), .e(new_n140), .o1(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n139), .b(new_n143), .c(new_n146), .out0(\s[13] ));
  orn002aa1n02x5               g052(.a(\a[13] ), .b(\b[12] ), .o(new_n148));
  160nm_ficinv00aa1n08x5       g053(.clk(new_n101), .clkout(new_n149));
  xorc02aa1n02x5               g054(.a(\a[3] ), .b(\b[2] ), .out0(new_n150));
  and002aa1n02x5               g055(.a(\b[0] ), .b(\a[1] ), .o(new_n151));
  oaoi03aa1n02x5               g056(.a(\a[2] ), .b(\b[1] ), .c(new_n151), .o1(new_n152));
  160nm_ficinv00aa1n08x5       g057(.clk(new_n105), .clkout(new_n153));
  aoai13aa1n02x5               g058(.a(new_n149), .b(new_n153), .c(new_n152), .d(new_n150), .o1(new_n154));
  nanp03aa1n02x5               g059(.a(new_n117), .b(new_n112), .c(new_n113), .o1(new_n155));
  160nm_ficinv00aa1n08x5       g060(.clk(new_n118), .clkout(new_n156));
  160nm_ficinv00aa1n08x5       g061(.clk(new_n122), .clkout(new_n157));
  aoi113aa1n02x5               g062(.a(new_n107), .b(new_n116), .c(new_n117), .d(new_n156), .e(new_n157), .o1(new_n158));
  oai012aa1n02x5               g063(.a(new_n158), .b(new_n155), .c(new_n154), .o1(new_n159));
  nanp03aa1n02x5               g064(.a(new_n135), .b(new_n137), .c(new_n140), .o1(new_n160));
  nona22aa1n02x4               g065(.a(new_n160), .b(new_n145), .c(new_n144), .out0(new_n161));
  aoai13aa1n02x5               g066(.a(new_n139), .b(new_n161), .c(new_n159), .d(new_n142), .o1(new_n162));
  xorc02aa1n02x5               g067(.a(\a[14] ), .b(\b[13] ), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n162), .c(new_n148), .out0(\s[14] ));
  and002aa1n02x5               g069(.a(new_n163), .b(new_n139), .o(new_n165));
  160nm_ficinv00aa1n08x5       g070(.clk(new_n165), .clkout(new_n166));
  nanp02aa1n02x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  oai022aa1n02x5               g072(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n168));
  nanp02aa1n02x5               g073(.a(new_n168), .b(new_n167), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n166), .c(new_n143), .d(new_n146), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n02x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n174), .b(new_n175), .out0(new_n176));
  160nm_ficinv00aa1n08x5       g081(.clk(new_n176), .clkout(new_n177));
  aoi112aa1n02x5               g082(.a(new_n177), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n178));
  aoai13aa1n02x5               g083(.a(new_n177), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  nano23aa1n02x4               g085(.a(new_n172), .b(new_n174), .c(new_n175), .d(new_n173), .out0(new_n181));
  nanp03aa1n02x5               g086(.a(new_n181), .b(new_n139), .c(new_n163), .o1(new_n182));
  norp02aa1n02x5               g087(.a(new_n182), .b(new_n141), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n183), .b(new_n124), .c(new_n106), .d(new_n114), .o1(new_n184));
  160nm_ficinv00aa1n08x5       g089(.clk(new_n182), .clkout(new_n185));
  nona23aa1n02x4               g090(.a(new_n175), .b(new_n173), .c(new_n172), .d(new_n174), .out0(new_n186));
  nanp02aa1n02x5               g091(.a(new_n172), .b(new_n175), .o1(new_n187));
  oai122aa1n02x7               g092(.a(new_n187), .b(new_n186), .c(new_n169), .d(\b[15] ), .e(\a[16] ), .o1(new_n188));
  aoi012aa1n02x5               g093(.a(new_n188), .b(new_n161), .c(new_n185), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n184), .b(new_n189), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g096(.clk(\a[18] ), .clkout(new_n192));
  160nm_ficinv00aa1n08x5       g097(.clk(\a[17] ), .clkout(new_n193));
  160nm_ficinv00aa1n08x5       g098(.clk(\b[16] ), .clkout(new_n194));
  oaoi03aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d04x5               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  oai022aa1n02x5               g102(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n198));
  oaib12aa1n02x5               g103(.a(new_n198), .b(new_n192), .c(\b[17] ), .out0(new_n199));
  160nm_ficinv00aa1n08x5       g104(.clk(new_n199), .clkout(new_n200));
  norp02aa1n02x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nanp02aa1n02x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  aoai13aa1n02x5               g108(.a(new_n203), .b(new_n200), .c(new_n190), .d(new_n197), .o1(new_n204));
  aoi112aa1n02x5               g109(.a(new_n203), .b(new_n200), .c(new_n190), .d(new_n197), .o1(new_n205));
  norb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  nona22aa1n02x4               g115(.a(new_n204), .b(new_n210), .c(new_n201), .out0(new_n211));
  orn002aa1n02x5               g116(.a(\a[19] ), .b(\b[18] ), .o(new_n212));
  aobi12aa1n02x5               g117(.a(new_n210), .b(new_n204), .c(new_n212), .out0(new_n213));
  norb02aa1n02x5               g118(.a(new_n211), .b(new_n213), .out0(\s[20] ));
  nano23aa1n02x4               g119(.a(new_n201), .b(new_n208), .c(new_n209), .d(new_n202), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n197), .b(new_n215), .o1(new_n216));
  nona23aa1n02x4               g121(.a(new_n209), .b(new_n202), .c(new_n201), .d(new_n208), .out0(new_n217));
  aoi012aa1n02x5               g122(.a(new_n208), .b(new_n201), .c(new_n209), .o1(new_n218));
  oai012aa1n02x5               g123(.a(new_n218), .b(new_n217), .c(new_n199), .o1(new_n219));
  160nm_ficinv00aa1n08x5       g124(.clk(new_n219), .clkout(new_n220));
  aoai13aa1n02x5               g125(.a(new_n220), .b(new_n216), .c(new_n184), .d(new_n189), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  xorc02aa1n02x5               g128(.a(\a[21] ), .b(\b[20] ), .out0(new_n224));
  xorc02aa1n02x5               g129(.a(\a[22] ), .b(\b[21] ), .out0(new_n225));
  aoi112aa1n02x5               g130(.a(new_n223), .b(new_n225), .c(new_n221), .d(new_n224), .o1(new_n226));
  aoai13aa1n02x5               g131(.a(new_n225), .b(new_n223), .c(new_n221), .d(new_n224), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n227), .b(new_n226), .out0(\s[22] ));
  160nm_ficinv00aa1n08x5       g133(.clk(\a[21] ), .clkout(new_n229));
  160nm_ficinv00aa1n08x5       g134(.clk(\a[22] ), .clkout(new_n230));
  xroi22aa1d04x5               g135(.a(new_n229), .b(\b[20] ), .c(new_n230), .d(\b[21] ), .out0(new_n231));
  nanp03aa1n02x5               g136(.a(new_n231), .b(new_n197), .c(new_n215), .o1(new_n232));
  160nm_ficinv00aa1n08x5       g137(.clk(\b[21] ), .clkout(new_n233));
  oaoi03aa1n02x5               g138(.a(new_n230), .b(new_n233), .c(new_n223), .o1(new_n234));
  160nm_ficinv00aa1n08x5       g139(.clk(new_n234), .clkout(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(new_n219), .c(new_n231), .o1(new_n236));
  aoai13aa1n02x5               g141(.a(new_n236), .b(new_n232), .c(new_n184), .d(new_n189), .o1(new_n237));
  xorb03aa1n02x5               g142(.a(new_n237), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  xorc02aa1n02x5               g144(.a(\a[23] ), .b(\b[22] ), .out0(new_n240));
  xorc02aa1n02x5               g145(.a(\a[24] ), .b(\b[23] ), .out0(new_n241));
  aoi112aa1n02x5               g146(.a(new_n239), .b(new_n241), .c(new_n237), .d(new_n240), .o1(new_n242));
  aoai13aa1n02x5               g147(.a(new_n241), .b(new_n239), .c(new_n237), .d(new_n240), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n243), .b(new_n242), .out0(\s[24] ));
  and002aa1n02x5               g149(.a(new_n241), .b(new_n240), .o(new_n245));
  160nm_ficinv00aa1n08x5       g150(.clk(new_n245), .clkout(new_n246));
  nano32aa1n02x4               g151(.a(new_n246), .b(new_n231), .c(new_n197), .d(new_n215), .out0(new_n247));
  160nm_ficinv00aa1n08x5       g152(.clk(new_n218), .clkout(new_n248));
  aoai13aa1n02x5               g153(.a(new_n231), .b(new_n248), .c(new_n215), .d(new_n200), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n250));
  oab012aa1n02x4               g155(.a(new_n250), .b(\a[24] ), .c(\b[23] ), .out0(new_n251));
  aoai13aa1n02x5               g156(.a(new_n251), .b(new_n246), .c(new_n249), .d(new_n234), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[25] ), .b(\b[24] ), .out0(new_n253));
  aoai13aa1n02x5               g158(.a(new_n253), .b(new_n252), .c(new_n190), .d(new_n247), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n253), .b(new_n252), .c(new_n190), .d(new_n247), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n254), .b(new_n255), .out0(\s[25] ));
  norp02aa1n02x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n02x5               g162(.a(\a[26] ), .b(\b[25] ), .out0(new_n258));
  nona22aa1n02x4               g163(.a(new_n254), .b(new_n258), .c(new_n257), .out0(new_n259));
  160nm_ficinv00aa1n08x5       g164(.clk(new_n257), .clkout(new_n260));
  aobi12aa1n02x5               g165(.a(new_n258), .b(new_n254), .c(new_n260), .out0(new_n261));
  norb02aa1n02x5               g166(.a(new_n259), .b(new_n261), .out0(\s[26] ));
  oabi12aa1n02x5               g167(.a(new_n188), .b(new_n146), .c(new_n182), .out0(new_n263));
  160nm_ficinv00aa1n08x5       g168(.clk(\a[25] ), .clkout(new_n264));
  160nm_ficinv00aa1n08x5       g169(.clk(\a[26] ), .clkout(new_n265));
  xroi22aa1d04x5               g170(.a(new_n264), .b(\b[24] ), .c(new_n265), .d(\b[25] ), .out0(new_n266));
  nano22aa1n02x4               g171(.a(new_n232), .b(new_n245), .c(new_n266), .out0(new_n267));
  aoai13aa1n02x5               g172(.a(new_n267), .b(new_n263), .c(new_n159), .d(new_n183), .o1(new_n268));
  oao003aa1n02x5               g173(.a(\a[26] ), .b(\b[25] ), .c(new_n260), .carry(new_n269));
  aobi12aa1n02x5               g174(.a(new_n269), .b(new_n252), .c(new_n266), .out0(new_n270));
  norp02aa1n02x5               g175(.a(\b[26] ), .b(\a[27] ), .o1(new_n271));
  nanp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  norb02aa1n02x5               g177(.a(new_n272), .b(new_n271), .out0(new_n273));
  xnbna2aa1n03x5               g178(.a(new_n273), .b(new_n270), .c(new_n268), .out0(\s[27] ));
  160nm_ficinv00aa1n08x5       g179(.clk(new_n271), .clkout(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[27] ), .b(\a[28] ), .out0(new_n276));
  160nm_ficinv00aa1n08x5       g181(.clk(new_n267), .clkout(new_n277));
  aoi012aa1n02x5               g182(.a(new_n277), .b(new_n184), .c(new_n189), .o1(new_n278));
  aoai13aa1n02x5               g183(.a(new_n245), .b(new_n235), .c(new_n219), .d(new_n231), .o1(new_n279));
  160nm_ficinv00aa1n08x5       g184(.clk(new_n266), .clkout(new_n280));
  aoai13aa1n02x5               g185(.a(new_n269), .b(new_n280), .c(new_n279), .d(new_n251), .o1(new_n281));
  oai012aa1n02x5               g186(.a(new_n272), .b(new_n281), .c(new_n278), .o1(new_n282));
  aoi012aa1n02x5               g187(.a(new_n276), .b(new_n282), .c(new_n275), .o1(new_n283));
  aobi12aa1n02x5               g188(.a(new_n272), .b(new_n270), .c(new_n268), .out0(new_n284));
  nano22aa1n02x4               g189(.a(new_n284), .b(new_n275), .c(new_n276), .out0(new_n285));
  norp02aa1n02x5               g190(.a(new_n283), .b(new_n285), .o1(\s[28] ));
  nano22aa1n02x4               g191(.a(new_n276), .b(new_n275), .c(new_n272), .out0(new_n287));
  oai012aa1n02x5               g192(.a(new_n287), .b(new_n281), .c(new_n278), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n275), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[28] ), .b(\a[29] ), .out0(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  aobi12aa1n02x5               g196(.a(new_n287), .b(new_n270), .c(new_n268), .out0(new_n292));
  nano22aa1n02x4               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  norp02aa1n02x5               g198(.a(new_n291), .b(new_n293), .o1(\s[29] ));
  xnrb03aa1n02x5               g199(.a(new_n151), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g200(.a(new_n273), .b(new_n290), .c(new_n276), .out0(new_n296));
  oai012aa1n02x5               g201(.a(new_n296), .b(new_n281), .c(new_n278), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[29] ), .b(\a[30] ), .out0(new_n299));
  aoi012aa1n02x5               g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x5               g205(.a(new_n296), .b(new_n270), .c(new_n268), .out0(new_n301));
  nano22aa1n02x4               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n02x5               g207(.a(new_n300), .b(new_n302), .o1(\s[30] ));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  norb03aa1n02x5               g209(.a(new_n287), .b(new_n299), .c(new_n290), .out0(new_n305));
  aobi12aa1n02x5               g210(.a(new_n305), .b(new_n270), .c(new_n268), .out0(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n307));
  nano22aa1n02x4               g212(.a(new_n306), .b(new_n304), .c(new_n307), .out0(new_n308));
  oai012aa1n02x5               g213(.a(new_n305), .b(new_n281), .c(new_n278), .o1(new_n309));
  aoi012aa1n02x5               g214(.a(new_n304), .b(new_n309), .c(new_n307), .o1(new_n310));
  norp02aa1n02x5               g215(.a(new_n310), .b(new_n308), .o1(\s[31] ));
  xnrb03aa1n02x5               g216(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g217(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g219(.a(new_n154), .b(\b[4] ), .c(new_n119), .out0(\s[5] ));
  oaoi03aa1n02x5               g220(.a(new_n119), .b(new_n121), .c(new_n106), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[5] ), .c(new_n120), .out0(\s[6] ));
  oaoi03aa1n02x5               g222(.a(\a[6] ), .b(\b[5] ), .c(new_n316), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g224(.a(new_n109), .b(new_n318), .c(new_n110), .o1(new_n320));
  xnrb03aa1n02x5               g225(.a(new_n320), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g226(.a(new_n125), .b(new_n115), .c(new_n158), .out0(\s[9] ));
endmodule


