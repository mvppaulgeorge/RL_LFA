// Benchmark "adder" written by ABC on Wed Jul 17 13:01:51 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n347, new_n349, new_n352, new_n354, new_n355,
    new_n357, new_n358, new_n359, new_n361, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n12x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  nor042aa1n03x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nand42aa1n03x5               g006(.a(\b[8] ), .b(\a[9] ), .o1(new_n102));
  nor022aa1n12x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand42aa1d28x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand22aa1n12x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  norb03aa1d15x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n106));
  inv000aa1d42x5               g011(.a(new_n106), .o1(new_n107));
  xnrc02aa1n12x5               g012(.a(\b[3] ), .b(\a[4] ), .out0(new_n108));
  nor022aa1n16x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nand42aa1n03x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nanb03aa1n09x5               g015(.a(new_n109), .b(new_n110), .c(new_n104), .out0(new_n111));
  nona22aa1n09x5               g016(.a(new_n107), .b(new_n111), .c(new_n108), .out0(new_n112));
  inv020aa1n02x5               g017(.a(new_n109), .o1(new_n113));
  oao003aa1n09x5               g018(.a(\a[4] ), .b(\b[3] ), .c(new_n113), .carry(new_n114));
  nor042aa1n04x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand02aa1d24x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nor002aa1n20x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nand02aa1n12x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nano23aa1n06x5               g023(.a(new_n115), .b(new_n117), .c(new_n118), .d(new_n116), .out0(new_n119));
  nor002aa1n03x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nand02aa1d08x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  norb02aa1n03x5               g026(.a(new_n121), .b(new_n120), .out0(new_n122));
  tech160nm_fixorc02aa1n04x5   g027(.a(\a[5] ), .b(\b[4] ), .out0(new_n123));
  nanp03aa1n02x5               g028(.a(new_n119), .b(new_n122), .c(new_n123), .o1(new_n124));
  nor002aa1d32x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  tech160nm_fioaoi03aa1n03p5x5 g031(.a(\a[6] ), .b(\b[5] ), .c(new_n126), .o1(new_n127));
  aoi012aa1n02x7               g032(.a(new_n115), .b(new_n117), .c(new_n116), .o1(new_n128));
  aobi12aa1n02x5               g033(.a(new_n128), .b(new_n119), .c(new_n127), .out0(new_n129));
  aoai13aa1n04x5               g034(.a(new_n129), .b(new_n124), .c(new_n112), .d(new_n114), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n100), .b(new_n101), .c(new_n130), .d(new_n102), .o1(new_n131));
  oai013aa1d12x5               g036(.a(new_n114), .b(new_n106), .c(new_n111), .d(new_n108), .o1(new_n132));
  nona23aa1n02x4               g037(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n133));
  nano22aa1n03x7               g038(.a(new_n133), .b(new_n123), .c(new_n122), .out0(new_n134));
  nanp02aa1n06x5               g039(.a(new_n119), .b(new_n127), .o1(new_n135));
  nand02aa1d04x5               g040(.a(new_n135), .b(new_n128), .o1(new_n136));
  aoai13aa1n02x5               g041(.a(new_n102), .b(new_n136), .c(new_n132), .d(new_n134), .o1(new_n137));
  nona22aa1n02x4               g042(.a(new_n137), .b(new_n101), .c(new_n100), .out0(new_n138));
  nanp02aa1n02x5               g043(.a(new_n131), .b(new_n138), .o1(\s[10] ));
  nand02aa1d04x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nor002aa1n16x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nano22aa1n02x4               g046(.a(new_n141), .b(new_n98), .c(new_n140), .out0(new_n142));
  nanp02aa1n02x5               g047(.a(new_n138), .b(new_n142), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n141), .o1(new_n144));
  aoi022aa1n02x5               g049(.a(new_n138), .b(new_n98), .c(new_n144), .d(new_n140), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n143), .b(new_n145), .out0(\s[11] ));
  nor002aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanp02aa1n06x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  nona23aa1n02x4               g054(.a(new_n143), .b(new_n148), .c(new_n147), .d(new_n141), .out0(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n149), .c(new_n144), .d(new_n143), .o1(\s[12] ));
  nano23aa1n06x5               g056(.a(new_n147), .b(new_n141), .c(new_n148), .d(new_n140), .out0(new_n152));
  norb02aa1n03x5               g057(.a(new_n102), .b(new_n101), .out0(new_n153));
  and003aa1n02x5               g058(.a(new_n152), .b(new_n99), .c(new_n153), .o(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n136), .c(new_n132), .d(new_n134), .o1(new_n155));
  tech160nm_fiao0012aa1n02p5x5 g060(.a(new_n97), .b(new_n101), .c(new_n98), .o(new_n156));
  aoi012aa1n02x7               g061(.a(new_n147), .b(new_n141), .c(new_n148), .o1(new_n157));
  aobi12aa1n02x5               g062(.a(new_n157), .b(new_n152), .c(new_n156), .out0(new_n158));
  tech160nm_finand02aa1n05x5   g063(.a(new_n155), .b(new_n158), .o1(new_n159));
  xorc02aa1n12x5               g064(.a(\a[13] ), .b(\b[12] ), .out0(new_n160));
  nand42aa1n02x5               g065(.a(new_n152), .b(new_n156), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n160), .o1(new_n162));
  and003aa1n02x5               g067(.a(new_n161), .b(new_n162), .c(new_n157), .o(new_n163));
  aoi022aa1n02x5               g068(.a(new_n159), .b(new_n160), .c(new_n155), .d(new_n163), .o1(\s[13] ));
  nor002aa1n06x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  xorc02aa1n12x5               g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n165), .c(new_n159), .d(new_n160), .o1(new_n168));
  inv000aa1d42x5               g073(.a(\b[13] ), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\a[14] ), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n165), .b(new_n170), .c(new_n169), .o1(new_n171));
  oaib12aa1n02x5               g076(.a(new_n171), .b(new_n169), .c(\a[14] ), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n168), .b(new_n172), .c(new_n160), .d(new_n159), .o1(\s[14] ));
  and002aa1n02x5               g078(.a(new_n166), .b(new_n160), .o(new_n174));
  oaoi03aa1n12x5               g079(.a(new_n170), .b(new_n169), .c(new_n165), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  nor042aa1n12x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand42aa1n04x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  aoai13aa1n04x5               g084(.a(new_n179), .b(new_n176), .c(new_n159), .d(new_n174), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n176), .c(new_n159), .d(new_n174), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(\s[15] ));
  inv000aa1d42x5               g087(.a(new_n177), .o1(new_n183));
  nor042aa1n04x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand42aa1n06x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  norb03aa1n02x5               g091(.a(new_n185), .b(new_n177), .c(new_n184), .out0(new_n187));
  nand42aa1n03x5               g092(.a(new_n180), .b(new_n187), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n186), .c(new_n183), .d(new_n180), .o1(\s[16] ));
  nano23aa1n09x5               g094(.a(new_n177), .b(new_n184), .c(new_n185), .d(new_n178), .out0(new_n190));
  nand23aa1n06x5               g095(.a(new_n190), .b(new_n160), .c(new_n166), .o1(new_n191));
  nano32aa1n03x7               g096(.a(new_n191), .b(new_n153), .c(new_n152), .d(new_n99), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n136), .c(new_n132), .d(new_n134), .o1(new_n193));
  aoi012aa1n02x7               g098(.a(new_n191), .b(new_n161), .c(new_n157), .o1(new_n194));
  aoi012aa1n02x5               g099(.a(new_n184), .b(new_n177), .c(new_n185), .o1(new_n195));
  oaib12aa1n09x5               g100(.a(new_n195), .b(new_n175), .c(new_n190), .out0(new_n196));
  nor042aa1n06x5               g101(.a(new_n194), .b(new_n196), .o1(new_n197));
  nanp02aa1n09x5               g102(.a(new_n193), .b(new_n197), .o1(new_n198));
  tech160nm_fixorc02aa1n03p5x5 g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  nanb02aa1n02x5               g104(.a(new_n199), .b(new_n195), .out0(new_n200));
  aoi112aa1n02x5               g105(.a(new_n194), .b(new_n200), .c(new_n176), .d(new_n190), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n198), .b(new_n199), .c(new_n193), .d(new_n201), .o1(\s[17] ));
  aobi12aa1n02x5               g107(.a(new_n199), .b(new_n193), .c(new_n197), .out0(new_n203));
  nor042aa1n04x5               g108(.a(\b[16] ), .b(\a[17] ), .o1(new_n204));
  aoi012aa1n02x5               g109(.a(new_n204), .b(new_n198), .c(new_n199), .o1(new_n205));
  norp02aa1n06x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand22aa1n04x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  norb02aa1n03x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  nona22aa1n02x4               g113(.a(new_n207), .b(new_n206), .c(new_n204), .out0(new_n209));
  oai022aa1n02x5               g114(.a(new_n205), .b(new_n208), .c(new_n209), .d(new_n203), .o1(\s[18] ));
  and002aa1n02x5               g115(.a(new_n199), .b(new_n208), .o(new_n211));
  tech160nm_fiaoi012aa1n04x5   g116(.a(new_n206), .b(new_n204), .c(new_n207), .o1(new_n212));
  inv020aa1n04x5               g117(.a(new_n212), .o1(new_n213));
  nor042aa1d18x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand02aa1n03x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n213), .c(new_n198), .d(new_n211), .o1(new_n217));
  aoi112aa1n02x5               g122(.a(new_n216), .b(new_n213), .c(new_n198), .d(new_n211), .o1(new_n218));
  norb02aa1n02x7               g123(.a(new_n217), .b(new_n218), .out0(\s[19] ));
  xnrc02aa1n02x5               g124(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g125(.a(new_n214), .o1(new_n221));
  nor042aa1n04x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanp02aa1n04x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  norb03aa1n02x5               g129(.a(new_n223), .b(new_n214), .c(new_n222), .out0(new_n225));
  nanp02aa1n06x5               g130(.a(new_n217), .b(new_n225), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n224), .c(new_n221), .d(new_n217), .o1(\s[20] ));
  nona23aa1n09x5               g132(.a(new_n223), .b(new_n215), .c(new_n214), .d(new_n222), .out0(new_n228));
  nano22aa1n03x7               g133(.a(new_n228), .b(new_n199), .c(new_n208), .out0(new_n229));
  aoi012aa1n06x5               g134(.a(new_n222), .b(new_n214), .c(new_n223), .o1(new_n230));
  tech160nm_fioai012aa1n05x5   g135(.a(new_n230), .b(new_n228), .c(new_n212), .o1(new_n231));
  nor042aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n231), .c(new_n198), .d(new_n229), .o1(new_n235));
  nano23aa1n09x5               g140(.a(new_n214), .b(new_n222), .c(new_n223), .d(new_n215), .out0(new_n236));
  inv030aa1n03x5               g141(.a(new_n230), .o1(new_n237));
  aoi112aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n236), .d(new_n213), .o1(new_n238));
  aobi12aa1n02x5               g143(.a(new_n238), .b(new_n198), .c(new_n229), .out0(new_n239));
  norb02aa1n03x4               g144(.a(new_n235), .b(new_n239), .out0(\s[21] ));
  inv000aa1d42x5               g145(.a(new_n232), .o1(new_n241));
  nor042aa1n02x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  and002aa1n06x5               g147(.a(\b[21] ), .b(\a[22] ), .o(new_n243));
  norp02aa1n02x5               g148(.a(new_n243), .b(new_n242), .o1(new_n244));
  norp03aa1n02x5               g149(.a(new_n243), .b(new_n242), .c(new_n232), .o1(new_n245));
  nanp02aa1n06x5               g150(.a(new_n235), .b(new_n245), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n244), .c(new_n241), .d(new_n235), .o1(\s[22] ));
  nano23aa1n06x5               g152(.a(new_n243), .b(new_n242), .c(new_n241), .d(new_n233), .out0(new_n248));
  nano32aa1n02x4               g153(.a(new_n228), .b(new_n248), .c(new_n199), .d(new_n208), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n248), .b(new_n237), .c(new_n236), .d(new_n213), .o1(new_n250));
  oab012aa1n04x5               g155(.a(new_n242), .b(new_n241), .c(new_n243), .out0(new_n251));
  nanp02aa1n02x5               g156(.a(new_n250), .b(new_n251), .o1(new_n252));
  nor022aa1n16x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  nand42aa1n03x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n252), .c(new_n198), .d(new_n249), .o1(new_n256));
  inv040aa1n03x5               g161(.a(new_n251), .o1(new_n257));
  nona22aa1n02x4               g162(.a(new_n250), .b(new_n257), .c(new_n255), .out0(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(new_n198), .c(new_n249), .o1(new_n259));
  norb02aa1n03x4               g164(.a(new_n256), .b(new_n259), .out0(\s[23] ));
  inv000aa1d42x5               g165(.a(new_n253), .o1(new_n261));
  nor022aa1n04x5               g166(.a(\b[23] ), .b(\a[24] ), .o1(new_n262));
  and002aa1n06x5               g167(.a(\b[23] ), .b(\a[24] ), .o(new_n263));
  norp02aa1n02x5               g168(.a(new_n263), .b(new_n262), .o1(new_n264));
  norp03aa1n02x5               g169(.a(new_n263), .b(new_n262), .c(new_n253), .o1(new_n265));
  nanp02aa1n06x5               g170(.a(new_n256), .b(new_n265), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n266), .b(new_n264), .c(new_n261), .d(new_n256), .o1(\s[24] ));
  inv000aa1n02x5               g172(.a(new_n229), .o1(new_n268));
  nano23aa1d18x5               g173(.a(new_n263), .b(new_n262), .c(new_n261), .d(new_n254), .out0(new_n269));
  nano22aa1n02x5               g174(.a(new_n268), .b(new_n248), .c(new_n269), .out0(new_n270));
  inv000aa1d42x5               g175(.a(new_n269), .o1(new_n271));
  oab012aa1n02x4               g176(.a(new_n262), .b(new_n261), .c(new_n263), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n271), .c(new_n250), .d(new_n251), .o1(new_n273));
  tech160nm_fixorc02aa1n04x5   g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n198), .d(new_n270), .o1(new_n275));
  nanb02aa1n02x5               g180(.a(new_n274), .b(new_n272), .out0(new_n276));
  aoi122aa1n06x5               g181(.a(new_n276), .b(new_n252), .c(new_n269), .d(new_n198), .e(new_n270), .o1(new_n277));
  norb02aa1n02x7               g182(.a(new_n275), .b(new_n277), .out0(\s[25] ));
  nor042aa1n03x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  norp02aa1n02x5               g185(.a(\b[25] ), .b(\a[26] ), .o1(new_n281));
  and002aa1n03x5               g186(.a(\b[25] ), .b(\a[26] ), .o(new_n282));
  nor022aa1n04x5               g187(.a(new_n282), .b(new_n281), .o1(new_n283));
  norp03aa1n02x5               g188(.a(new_n282), .b(new_n281), .c(new_n279), .o1(new_n284));
  nand02aa1n04x5               g189(.a(new_n275), .b(new_n284), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n283), .c(new_n280), .d(new_n275), .o1(\s[26] ));
  and002aa1n09x5               g191(.a(new_n274), .b(new_n283), .o(new_n287));
  nano32aa1n03x7               g192(.a(new_n268), .b(new_n287), .c(new_n248), .d(new_n269), .out0(new_n288));
  aobi12aa1n06x5               g193(.a(new_n288), .b(new_n193), .c(new_n197), .out0(new_n289));
  aoai13aa1n04x5               g194(.a(new_n269), .b(new_n257), .c(new_n231), .d(new_n248), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n287), .o1(new_n291));
  oab012aa1n02x4               g196(.a(new_n281), .b(new_n280), .c(new_n282), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n291), .c(new_n290), .d(new_n272), .o1(new_n293));
  xorc02aa1n02x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  inv000aa1n02x5               g199(.a(new_n294), .o1(new_n295));
  nanp02aa1n02x5               g200(.a(new_n292), .b(new_n295), .o1(new_n296));
  aoi112aa1n03x4               g201(.a(new_n289), .b(new_n296), .c(new_n273), .d(new_n287), .o1(new_n297));
  oaoi13aa1n02x7               g202(.a(new_n297), .b(new_n294), .c(new_n289), .d(new_n293), .o1(\s[27] ));
  norp02aa1n02x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  oaih12aa1n02x5               g205(.a(new_n294), .b(new_n293), .c(new_n289), .o1(new_n301));
  norp02aa1n02x5               g206(.a(\b[27] ), .b(\a[28] ), .o1(new_n302));
  and002aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .o(new_n303));
  norp02aa1n02x5               g208(.a(new_n303), .b(new_n302), .o1(new_n304));
  oabi12aa1n03x5               g209(.a(new_n196), .b(new_n158), .c(new_n191), .out0(new_n305));
  aoai13aa1n06x5               g210(.a(new_n288), .b(new_n305), .c(new_n130), .d(new_n192), .o1(new_n306));
  aobi12aa1n06x5               g211(.a(new_n292), .b(new_n273), .c(new_n287), .out0(new_n307));
  norp03aa1n02x5               g212(.a(new_n303), .b(new_n302), .c(new_n299), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n295), .c(new_n307), .d(new_n306), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n301), .d(new_n300), .o1(\s[28] ));
  inv000aa1d42x5               g215(.a(\a[27] ), .o1(new_n311));
  inv000aa1d42x5               g216(.a(\a[28] ), .o1(new_n312));
  xroi22aa1d04x5               g217(.a(new_n311), .b(\b[26] ), .c(new_n312), .d(\b[27] ), .out0(new_n313));
  oaih12aa1n02x5               g218(.a(new_n313), .b(new_n293), .c(new_n289), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  aoi112aa1n09x5               g220(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n316));
  oai022aa1n02x5               g221(.a(\a[28] ), .b(\b[27] ), .c(\b[28] ), .d(\a[29] ), .o1(new_n317));
  aoi112aa1n02x5               g222(.a(new_n316), .b(new_n317), .c(\a[29] ), .d(\b[28] ), .o1(new_n318));
  aoai13aa1n06x5               g223(.a(new_n318), .b(new_n315), .c(new_n307), .d(new_n306), .o1(new_n319));
  nor042aa1n03x5               g224(.a(new_n316), .b(new_n302), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n319), .b(new_n321), .c(new_n314), .d(new_n320), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g228(.a(new_n295), .b(new_n321), .c(new_n304), .out0(new_n324));
  oaih12aa1n02x5               g229(.a(new_n324), .b(new_n293), .c(new_n289), .o1(new_n325));
  tech160nm_fioaoi03aa1n03p5x5 g230(.a(\a[29] ), .b(\b[28] ), .c(new_n320), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n326), .o1(new_n327));
  norp02aa1n02x5               g232(.a(\b[29] ), .b(\a[30] ), .o1(new_n328));
  nanp02aa1n02x5               g233(.a(\b[29] ), .b(\a[30] ), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n329), .b(new_n328), .out0(new_n330));
  inv000aa1n02x5               g235(.a(new_n324), .o1(new_n331));
  inv000aa1d42x5               g236(.a(\a[29] ), .o1(new_n332));
  obai22aa1n02x7               g237(.a(\b[28] ), .b(new_n332), .c(new_n316), .d(new_n302), .out0(new_n333));
  oai022aa1n02x5               g238(.a(\a[29] ), .b(\b[28] ), .c(\b[29] ), .d(\a[30] ), .o1(new_n334));
  nano22aa1n02x4               g239(.a(new_n334), .b(new_n333), .c(new_n329), .out0(new_n335));
  aoai13aa1n02x7               g240(.a(new_n335), .b(new_n331), .c(new_n307), .d(new_n306), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n330), .c(new_n325), .d(new_n327), .o1(\s[30] ));
  nano32aa1n02x4               g242(.a(new_n295), .b(new_n330), .c(new_n304), .d(new_n321), .out0(new_n338));
  oaih12aa1n02x5               g243(.a(new_n338), .b(new_n293), .c(new_n289), .o1(new_n339));
  xnrc02aa1n02x5               g244(.a(\b[30] ), .b(\a[31] ), .out0(new_n340));
  inv000aa1d42x5               g245(.a(new_n340), .o1(new_n341));
  inv000aa1n02x5               g246(.a(new_n338), .o1(new_n342));
  aoi112aa1n02x5               g247(.a(new_n328), .b(new_n340), .c(new_n326), .d(new_n330), .o1(new_n343));
  aoai13aa1n04x5               g248(.a(new_n343), .b(new_n342), .c(new_n307), .d(new_n306), .o1(new_n344));
  aoi012aa1n02x5               g249(.a(new_n328), .b(new_n326), .c(new_n330), .o1(new_n345));
  aoai13aa1n03x5               g250(.a(new_n344), .b(new_n341), .c(new_n339), .d(new_n345), .o1(\s[31] ));
  norb02aa1n02x5               g251(.a(new_n110), .b(new_n109), .out0(new_n347));
  xobna2aa1n03x5               g252(.a(new_n347), .b(new_n107), .c(new_n104), .out0(\s[3] ));
  oai112aa1n02x5               g253(.a(new_n347), .b(new_n104), .c(new_n105), .d(new_n103), .o1(new_n349));
  xobna2aa1n03x5               g254(.a(new_n108), .b(new_n349), .c(new_n113), .out0(\s[4] ));
  xnbna2aa1n03x5               g255(.a(new_n123), .b(new_n112), .c(new_n114), .out0(\s[5] ));
  nanp02aa1n02x5               g256(.a(new_n132), .b(new_n123), .o1(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n122), .b(new_n352), .c(new_n126), .out0(\s[6] ));
  nanb02aa1n02x5               g258(.a(new_n117), .b(new_n118), .out0(new_n354));
  nanp03aa1n02x5               g259(.a(new_n352), .b(new_n122), .c(new_n126), .o1(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n354), .b(new_n355), .c(new_n121), .out0(\s[7] ));
  norb02aa1n02x5               g261(.a(new_n116), .b(new_n115), .out0(new_n357));
  inv000aa1d42x5               g262(.a(new_n117), .o1(new_n358));
  nanb03aa1n02x5               g263(.a(new_n354), .b(new_n355), .c(new_n121), .out0(new_n359));
  xnbna2aa1n03x5               g264(.a(new_n357), .b(new_n359), .c(new_n358), .out0(\s[8] ));
  aoi012aa1n02x5               g265(.a(new_n124), .b(new_n112), .c(new_n114), .o1(new_n361));
  nanp03aa1n02x5               g266(.a(new_n135), .b(new_n128), .c(new_n153), .o1(new_n362));
  obai22aa1n02x7               g267(.a(new_n130), .b(new_n153), .c(new_n361), .d(new_n362), .out0(\s[9] ));
endmodule


