// Benchmark "adder" written by ABC on Thu Jul 18 08:05:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n340, new_n343, new_n345, new_n346, new_n347, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nand02aa1n06x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nor002aa1d32x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nand42aa1n04x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nona23aa1n09x5               g005(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n101));
  nor022aa1n16x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nanb02aa1n02x5               g008(.a(new_n102), .b(new_n103), .out0(new_n104));
  xnrc02aa1n02x5               g009(.a(\b[4] ), .b(\a[5] ), .out0(new_n105));
  nor043aa1n04x5               g010(.a(new_n101), .b(new_n104), .c(new_n105), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\a[2] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[1] ), .o1(new_n108));
  nand22aa1n04x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  tech160nm_fioaoi03aa1n05x5   g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  nor002aa1n06x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nand22aa1n03x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nor022aa1n06x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  nona23aa1n03x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  tech160nm_fiao0012aa1n02p5x5 g020(.a(new_n111), .b(new_n113), .c(new_n112), .o(new_n116));
  oabi12aa1n06x5               g021(.a(new_n116), .b(new_n115), .c(new_n110), .out0(new_n117));
  inv000aa1d42x5               g022(.a(new_n97), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(new_n99), .b(new_n98), .o1(new_n119));
  nor042aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  tech160nm_fioai012aa1n03p5x5 g025(.a(new_n103), .b(new_n120), .c(new_n102), .o1(new_n121));
  oai112aa1n04x5               g026(.a(new_n118), .b(new_n119), .c(new_n101), .d(new_n121), .o1(new_n122));
  aoi012aa1n06x5               g027(.a(new_n122), .b(new_n117), .c(new_n106), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .c(new_n123), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n04x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  tech160nm_finand02aa1n03p5x5 g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  norb02aa1n03x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  nor042aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  nand42aa1n03x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nor002aa1n03x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nand42aa1n06x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nano23aa1n03x7               g037(.a(new_n129), .b(new_n131), .c(new_n132), .d(new_n130), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n122), .c(new_n117), .d(new_n106), .o1(new_n134));
  oai012aa1n06x5               g039(.a(new_n132), .b(new_n131), .c(new_n129), .o1(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n128), .b(new_n134), .c(new_n135), .out0(\s[11] ));
  nanp02aa1n02x5               g041(.a(new_n134), .b(new_n135), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n126), .b(new_n137), .c(new_n127), .o1(new_n138));
  nor002aa1d24x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n138), .b(new_n141), .c(new_n140), .out0(\s[12] ));
  nand42aa1n03x5               g047(.a(new_n126), .b(new_n141), .o1(new_n143));
  nona23aa1n09x5               g048(.a(new_n141), .b(new_n127), .c(new_n126), .d(new_n139), .out0(new_n144));
  oai112aa1n06x5               g049(.a(new_n143), .b(new_n140), .c(new_n144), .d(new_n135), .o1(new_n145));
  norb02aa1n02x7               g050(.a(new_n141), .b(new_n139), .out0(new_n146));
  nano32aa1n03x7               g051(.a(new_n123), .b(new_n146), .c(new_n128), .d(new_n133), .out0(new_n147));
  nor042aa1d18x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  tech160nm_finand02aa1n03p5x5 g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nanb02aa1n02x5               g054(.a(new_n148), .b(new_n149), .out0(new_n150));
  oabi12aa1n02x5               g055(.a(new_n150), .b(new_n147), .c(new_n145), .out0(new_n151));
  inv020aa1n02x5               g056(.a(new_n148), .o1(new_n152));
  aoi112aa1n02x5               g057(.a(new_n147), .b(new_n145), .c(new_n152), .d(new_n149), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n151), .b(new_n153), .out0(\s[13] ));
  nor002aa1n02x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nand42aa1n03x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nanb02aa1n02x5               g061(.a(new_n155), .b(new_n156), .out0(new_n157));
  xobna2aa1n03x5               g062(.a(new_n157), .b(new_n151), .c(new_n152), .out0(\s[14] ));
  nano23aa1n06x5               g063(.a(new_n148), .b(new_n155), .c(new_n156), .d(new_n149), .out0(new_n159));
  oaoi03aa1n09x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n152), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n160), .b(new_n145), .c(new_n159), .o1(new_n161));
  nano23aa1n02x4               g066(.a(new_n97), .b(new_n99), .c(new_n100), .d(new_n98), .out0(new_n162));
  nona22aa1n02x4               g067(.a(new_n162), .b(new_n105), .c(new_n104), .out0(new_n163));
  oao003aa1n02x5               g068(.a(new_n107), .b(new_n108), .c(new_n109), .carry(new_n164));
  nano23aa1n02x4               g069(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n165));
  aoi012aa1n03x5               g070(.a(new_n116), .b(new_n165), .c(new_n164), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n97), .b(new_n98), .out0(new_n167));
  nanb02aa1n12x5               g072(.a(new_n99), .b(new_n100), .out0(new_n168));
  norp03aa1n02x5               g073(.a(new_n121), .b(new_n168), .c(new_n167), .o1(new_n169));
  nano22aa1n02x4               g074(.a(new_n169), .b(new_n118), .c(new_n119), .out0(new_n170));
  oai012aa1n02x5               g075(.a(new_n170), .b(new_n166), .c(new_n163), .o1(new_n171));
  nona23aa1n02x4               g076(.a(new_n132), .b(new_n130), .c(new_n129), .d(new_n131), .out0(new_n172));
  nona23aa1n02x4               g077(.a(new_n156), .b(new_n149), .c(new_n148), .d(new_n155), .out0(new_n173));
  nona32aa1n02x4               g078(.a(new_n171), .b(new_n173), .c(new_n144), .d(new_n172), .out0(new_n174));
  nor002aa1d32x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nand42aa1n04x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  xobna2aa1n03x5               g082(.a(new_n177), .b(new_n174), .c(new_n161), .out0(\s[15] ));
  inv000aa1d42x5               g083(.a(new_n175), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n179), .b(new_n177), .c(new_n174), .d(new_n161), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor002aa1n04x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nanp02aa1n12x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nano23aa1n06x5               g088(.a(new_n175), .b(new_n182), .c(new_n183), .d(new_n176), .out0(new_n184));
  aoi122aa1n12x5               g089(.a(new_n182), .b(new_n183), .c(new_n175), .d(new_n184), .e(new_n160), .o1(new_n185));
  nona23aa1n02x4               g090(.a(new_n183), .b(new_n176), .c(new_n175), .d(new_n182), .out0(new_n186));
  nona32aa1n09x5               g091(.a(new_n145), .b(new_n186), .c(new_n157), .d(new_n150), .out0(new_n187));
  nanp02aa1n03x5               g092(.a(new_n184), .b(new_n133), .o1(new_n188));
  nano32aa1n03x7               g093(.a(new_n188), .b(new_n159), .c(new_n146), .d(new_n128), .out0(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n122), .c(new_n117), .d(new_n106), .o1(new_n190));
  nand23aa1n09x5               g095(.a(new_n190), .b(new_n185), .c(new_n187), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d28x5               g097(.a(\a[17] ), .o1(new_n193));
  inv040aa1d32x5               g098(.a(\b[16] ), .o1(new_n194));
  oaoi03aa1n03x5               g099(.a(new_n193), .b(new_n194), .c(new_n191), .o1(new_n195));
  xnrb03aa1n03x5               g100(.a(new_n195), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv020aa1n03x5               g101(.a(new_n185), .o1(new_n197));
  aoi013aa1n06x4               g102(.a(new_n197), .b(new_n145), .c(new_n159), .d(new_n184), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(new_n194), .b(new_n193), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  nor002aa1d32x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand42aa1d28x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nano32aa1d12x5               g107(.a(new_n201), .b(new_n199), .c(new_n202), .d(new_n200), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n12x5               g109(.a(new_n202), .b(new_n201), .c(new_n193), .d(new_n194), .o1(new_n205));
  aoai13aa1n03x5               g110(.a(new_n205), .b(new_n204), .c(new_n198), .d(new_n190), .o1(new_n206));
  xorb03aa1n02x5               g111(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1d18x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nanp02aa1n03x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nanb02aa1n12x5               g115(.a(new_n209), .b(new_n210), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor042aa1n09x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanp02aa1n04x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1d24x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoi112aa1n03x4               g121(.a(new_n209), .b(new_n216), .c(new_n206), .d(new_n212), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n209), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n205), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n212), .b(new_n219), .c(new_n191), .d(new_n203), .o1(new_n220));
  aoi012aa1n03x5               g125(.a(new_n215), .b(new_n220), .c(new_n218), .o1(new_n221));
  norp02aa1n03x5               g126(.a(new_n221), .b(new_n217), .o1(\s[20] ));
  nona22aa1d24x5               g127(.a(new_n203), .b(new_n211), .c(new_n215), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n213), .o1(new_n224));
  nand42aa1n03x5               g129(.a(new_n209), .b(new_n214), .o1(new_n225));
  nor043aa1n03x5               g130(.a(new_n205), .b(new_n211), .c(new_n215), .o1(new_n226));
  nano22aa1n02x4               g131(.a(new_n226), .b(new_n224), .c(new_n225), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n223), .c(new_n198), .d(new_n190), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  tech160nm_fixorc02aa1n03p5x5 g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xorc02aa1n12x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  aoi112aa1n03x4               g137(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n233));
  inv020aa1n02x5               g138(.a(new_n230), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n223), .o1(new_n235));
  nona23aa1n03x5               g140(.a(new_n214), .b(new_n210), .c(new_n209), .d(new_n213), .out0(new_n236));
  oai112aa1n06x5               g141(.a(new_n225), .b(new_n224), .c(new_n236), .d(new_n205), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n231), .b(new_n237), .c(new_n191), .d(new_n235), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n232), .o1(new_n239));
  aoi012aa1n03x5               g144(.a(new_n239), .b(new_n238), .c(new_n234), .o1(new_n240));
  norp02aa1n03x5               g145(.a(new_n240), .b(new_n233), .o1(\s[22] ));
  and002aa1n06x5               g146(.a(new_n232), .b(new_n231), .o(new_n242));
  oaoi03aa1n09x5               g147(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .o1(new_n243));
  aoi012aa1n12x5               g148(.a(new_n243), .b(new_n237), .c(new_n242), .o1(new_n244));
  nano22aa1n03x7               g149(.a(new_n223), .b(new_n231), .c(new_n232), .out0(new_n245));
  inv020aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  aoai13aa1n06x5               g151(.a(new_n244), .b(new_n246), .c(new_n198), .d(new_n190), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  nand42aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n250), .b(new_n249), .out0(new_n251));
  nor042aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  nanp02aa1n02x5               g157(.a(\b[23] ), .b(\a[24] ), .o1(new_n253));
  norb02aa1n02x5               g158(.a(new_n253), .b(new_n252), .out0(new_n254));
  aoi112aa1n02x7               g159(.a(new_n249), .b(new_n254), .c(new_n247), .d(new_n251), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n249), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n244), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n251), .b(new_n257), .c(new_n191), .d(new_n245), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n254), .o1(new_n259));
  tech160nm_fiaoi012aa1n02p5x5 g164(.a(new_n259), .b(new_n258), .c(new_n256), .o1(new_n260));
  nor042aa1n03x5               g165(.a(new_n260), .b(new_n255), .o1(\s[24] ));
  nano23aa1n06x5               g166(.a(new_n249), .b(new_n252), .c(new_n253), .d(new_n250), .out0(new_n262));
  nano32aa1n03x7               g167(.a(new_n223), .b(new_n262), .c(new_n231), .d(new_n232), .out0(new_n263));
  inv000aa1n02x5               g168(.a(new_n263), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n265));
  nand42aa1n03x5               g170(.a(new_n262), .b(new_n243), .o1(new_n266));
  nona22aa1n02x4               g171(.a(new_n266), .b(new_n265), .c(new_n252), .out0(new_n267));
  nand23aa1n02x5               g172(.a(new_n262), .b(new_n231), .c(new_n232), .o1(new_n268));
  inv000aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  aoi012aa1n09x5               g174(.a(new_n267), .b(new_n237), .c(new_n269), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n264), .c(new_n198), .d(new_n190), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  tech160nm_fixorc02aa1n03p5x5 g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xorc02aa1n12x5               g179(.a(\a[26] ), .b(\b[25] ), .out0(new_n275));
  aoi112aa1n03x4               g180(.a(new_n273), .b(new_n275), .c(new_n271), .d(new_n274), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n273), .o1(new_n277));
  inv000aa1n02x5               g182(.a(new_n270), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n274), .b(new_n278), .c(new_n191), .d(new_n263), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n275), .o1(new_n280));
  aoi012aa1n03x5               g185(.a(new_n280), .b(new_n279), .c(new_n277), .o1(new_n281));
  nor002aa1n02x5               g186(.a(new_n281), .b(new_n276), .o1(\s[26] ));
  nand02aa1n02x5               g187(.a(new_n187), .b(new_n185), .o1(new_n283));
  nor002aa1n02x5               g188(.a(new_n186), .b(new_n172), .o1(new_n284));
  nona22aa1n02x4               g189(.a(new_n284), .b(new_n173), .c(new_n144), .out0(new_n285));
  oaoi13aa1n04x5               g190(.a(new_n285), .b(new_n170), .c(new_n166), .d(new_n163), .o1(new_n286));
  and002aa1n24x5               g191(.a(new_n275), .b(new_n274), .o(new_n287));
  nano32aa1d12x5               g192(.a(new_n223), .b(new_n287), .c(new_n242), .d(new_n262), .out0(new_n288));
  oai012aa1n06x5               g193(.a(new_n288), .b(new_n283), .c(new_n286), .o1(new_n289));
  norp02aa1n02x5               g194(.a(\b[25] ), .b(\a[26] ), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  aoi112aa1n02x5               g196(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n292));
  inv000aa1n02x5               g197(.a(new_n292), .o1(new_n293));
  aoi112aa1n02x5               g198(.a(new_n265), .b(new_n252), .c(new_n262), .d(new_n243), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n287), .o1(new_n295));
  oaoi13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n227), .d(new_n268), .o1(new_n296));
  nano22aa1n03x7               g201(.a(new_n296), .b(new_n291), .c(new_n293), .out0(new_n297));
  xorc02aa1n12x5               g202(.a(\a[27] ), .b(\b[26] ), .out0(new_n298));
  xnbna2aa1n03x5               g203(.a(new_n298), .b(new_n289), .c(new_n297), .out0(\s[27] ));
  nor042aa1n03x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n298), .o1(new_n302));
  tech160nm_fiaoi012aa1n02p5x5 g207(.a(new_n302), .b(new_n289), .c(new_n297), .o1(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[27] ), .b(\a[28] ), .out0(new_n304));
  nano22aa1n02x4               g209(.a(new_n303), .b(new_n301), .c(new_n304), .out0(new_n305));
  aoai13aa1n04x5               g210(.a(new_n287), .b(new_n267), .c(new_n237), .d(new_n269), .o1(new_n306));
  nona22aa1n06x5               g211(.a(new_n306), .b(new_n292), .c(new_n290), .out0(new_n307));
  aoai13aa1n06x5               g212(.a(new_n298), .b(new_n307), .c(new_n191), .d(new_n288), .o1(new_n308));
  aoi012aa1n03x5               g213(.a(new_n304), .b(new_n308), .c(new_n301), .o1(new_n309));
  nor002aa1n02x5               g214(.a(new_n309), .b(new_n305), .o1(\s[28] ));
  norb02aa1n02x5               g215(.a(new_n298), .b(new_n304), .out0(new_n311));
  aoai13aa1n06x5               g216(.a(new_n311), .b(new_n307), .c(new_n191), .d(new_n288), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[28] ), .b(\b[27] ), .c(new_n301), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .out0(new_n314));
  aoi012aa1n03x5               g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  inv000aa1n02x5               g220(.a(new_n311), .o1(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n289), .c(new_n297), .o1(new_n317));
  nano22aa1n02x4               g222(.a(new_n317), .b(new_n313), .c(new_n314), .out0(new_n318));
  nor002aa1n02x5               g223(.a(new_n315), .b(new_n318), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n03x5               g225(.a(new_n298), .b(new_n314), .c(new_n304), .out0(new_n321));
  aoai13aa1n06x5               g226(.a(new_n321), .b(new_n307), .c(new_n191), .d(new_n288), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .carry(new_n323));
  xnrc02aa1n02x5               g228(.a(\b[29] ), .b(\a[30] ), .out0(new_n324));
  tech160nm_fiaoi012aa1n05x5   g229(.a(new_n324), .b(new_n322), .c(new_n323), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n321), .o1(new_n326));
  aoi012aa1n02x7               g231(.a(new_n326), .b(new_n289), .c(new_n297), .o1(new_n327));
  nano22aa1n02x4               g232(.a(new_n327), .b(new_n323), .c(new_n324), .out0(new_n328));
  nor002aa1n02x5               g233(.a(new_n325), .b(new_n328), .o1(\s[30] ));
  norb02aa1n06x5               g234(.a(new_n321), .b(new_n324), .out0(new_n330));
  inv000aa1n02x5               g235(.a(new_n330), .o1(new_n331));
  tech160nm_fiaoi012aa1n02p5x5 g236(.a(new_n331), .b(new_n289), .c(new_n297), .o1(new_n332));
  oao003aa1n02x5               g237(.a(\a[30] ), .b(\b[29] ), .c(new_n323), .carry(new_n333));
  xnrc02aa1n02x5               g238(.a(\b[30] ), .b(\a[31] ), .out0(new_n334));
  nano22aa1n02x4               g239(.a(new_n332), .b(new_n333), .c(new_n334), .out0(new_n335));
  aoai13aa1n04x5               g240(.a(new_n330), .b(new_n307), .c(new_n191), .d(new_n288), .o1(new_n336));
  aoi012aa1n03x5               g241(.a(new_n334), .b(new_n336), .c(new_n333), .o1(new_n337));
  nor002aa1n02x5               g242(.a(new_n337), .b(new_n335), .o1(\s[31] ));
  xnrb03aa1n02x5               g243(.a(new_n110), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g244(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n340));
  xorb03aa1n02x5               g245(.a(new_n340), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g246(.a(new_n117), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g247(.a(\a[5] ), .b(\b[4] ), .c(new_n166), .o1(new_n343));
  xorb03aa1n02x5               g248(.a(new_n343), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g249(.a(new_n168), .o1(new_n345));
  aoai13aa1n03x5               g250(.a(new_n345), .b(new_n102), .c(new_n343), .d(new_n103), .o1(new_n346));
  aoi112aa1n02x5               g251(.a(new_n345), .b(new_n102), .c(new_n343), .d(new_n103), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n346), .b(new_n347), .out0(\s[7] ));
  inv000aa1d42x5               g253(.a(new_n99), .o1(new_n349));
  xobna2aa1n03x5               g254(.a(new_n167), .b(new_n346), .c(new_n349), .out0(\s[8] ));
  xnrb03aa1n02x5               g255(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


