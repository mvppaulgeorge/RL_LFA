// Benchmark "adder" written by ABC on Thu Jul 18 11:22:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n313, new_n316, new_n318, new_n320, new_n321,
    new_n322, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n03p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  nor002aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n04x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n06x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aoi012aa1d24x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor042aa1n03x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  oa0012aa1n03x5               g012(.a(new_n104), .b(new_n105), .c(new_n103), .o(new_n108));
  oabi12aa1n18x5               g013(.a(new_n108), .b(new_n102), .c(new_n107), .out0(new_n109));
  xorc02aa1n02x5               g014(.a(\a[7] ), .b(\b[6] ), .out0(new_n110));
  tech160nm_fixorc02aa1n05x5   g015(.a(\a[5] ), .b(\b[4] ), .out0(new_n111));
  nand02aa1d06x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor042aa1n04x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1n12x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand42aa1n16x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nona23aa1n02x4               g020(.a(new_n112), .b(new_n115), .c(new_n114), .d(new_n113), .out0(new_n116));
  nano22aa1n03x7               g021(.a(new_n116), .b(new_n110), .c(new_n111), .out0(new_n117));
  orn002aa1n02x5               g022(.a(\a[7] ), .b(\b[6] ), .o(new_n118));
  inv000aa1d42x5               g023(.a(new_n114), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n115), .o1(new_n120));
  nand02aa1n10x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nor042aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  aoai13aa1n06x5               g027(.a(new_n121), .b(new_n113), .c(new_n122), .d(new_n112), .o1(new_n123));
  aoai13aa1n06x5               g028(.a(new_n119), .b(new_n120), .c(new_n123), .d(new_n118), .o1(new_n124));
  tech160nm_fixorc02aa1n03p5x5 g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  nand42aa1n03x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  nor002aa1n12x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nanb02aa1n02x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  nanp02aa1n02x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  inv040aa1n02x5               g036(.a(new_n102), .o1(new_n132));
  nano23aa1n02x5               g037(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n133));
  aoi012aa1n06x5               g038(.a(new_n108), .b(new_n133), .c(new_n132), .o1(new_n134));
  nano23aa1n02x4               g039(.a(new_n114), .b(new_n113), .c(new_n115), .d(new_n112), .out0(new_n135));
  nand03aa1n02x5               g040(.a(new_n135), .b(new_n110), .c(new_n111), .o1(new_n136));
  nanp02aa1n03x5               g041(.a(new_n123), .b(new_n118), .o1(new_n137));
  tech160nm_fiaoi012aa1n03p5x5 g042(.a(new_n114), .b(new_n137), .c(new_n115), .o1(new_n138));
  oai012aa1n12x5               g043(.a(new_n138), .b(new_n134), .c(new_n136), .o1(new_n139));
  oai022aa1d18x5               g044(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n131), .b(new_n140), .c(new_n139), .d(new_n125), .o1(new_n141));
  nano22aa1n02x4               g046(.a(new_n129), .b(new_n131), .c(new_n128), .out0(new_n142));
  aoai13aa1n03x5               g047(.a(new_n142), .b(new_n140), .c(new_n139), .d(new_n125), .o1(new_n143));
  aobi12aa1n02x5               g048(.a(new_n143), .b(new_n141), .c(new_n130), .out0(\s[11] ));
  inv000aa1d42x5               g049(.a(new_n129), .o1(new_n145));
  nor042aa1n03x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n02x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanb02aa1n02x5               g052(.a(new_n146), .b(new_n147), .out0(new_n148));
  xobna2aa1n03x5               g053(.a(new_n148), .b(new_n143), .c(new_n145), .out0(\s[12] ));
  nano23aa1n06x5               g054(.a(new_n146), .b(new_n129), .c(new_n147), .d(new_n128), .out0(new_n150));
  and003aa1n02x5               g055(.a(new_n150), .b(new_n125), .c(new_n97), .o(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n152));
  aoi022aa1n02x5               g057(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n129), .c(new_n140), .d(new_n131), .o1(new_n154));
  norb02aa1n03x4               g059(.a(new_n154), .b(new_n146), .out0(new_n155));
  nor042aa1n04x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1d28x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n157), .b(new_n156), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n152), .c(new_n155), .out0(\s[13] ));
  inv000aa1d42x5               g064(.a(\a[13] ), .o1(new_n160));
  inv000aa1d42x5               g065(.a(\b[12] ), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(new_n152), .b(new_n155), .o1(new_n162));
  oaoi03aa1n02x5               g067(.a(new_n160), .b(new_n161), .c(new_n162), .o1(new_n163));
  xnrb03aa1n02x5               g068(.a(new_n163), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n12x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand42aa1n16x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nano23aa1d15x5               g071(.a(new_n156), .b(new_n165), .c(new_n166), .d(new_n157), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n06x5               g073(.a(new_n166), .b(new_n165), .c(new_n160), .d(new_n161), .o1(new_n169));
  aoai13aa1n04x5               g074(.a(new_n169), .b(new_n168), .c(new_n152), .d(new_n155), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv000aa1d42x5               g076(.a(\a[15] ), .o1(new_n172));
  nanb02aa1n09x5               g077(.a(\b[14] ), .b(new_n172), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  tech160nm_fixorc02aa1n05x5   g079(.a(\a[15] ), .b(\b[14] ), .out0(new_n175));
  xorc02aa1n12x5               g080(.a(\a[16] ), .b(\b[15] ), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n174), .c(new_n170), .d(new_n175), .o1(new_n178));
  aoi112aa1n02x5               g083(.a(new_n174), .b(new_n177), .c(new_n170), .d(new_n175), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  nand23aa1d12x5               g085(.a(new_n167), .b(new_n175), .c(new_n176), .o1(new_n181));
  nano32aa1d12x5               g086(.a(new_n181), .b(new_n150), .c(new_n125), .d(new_n97), .out0(new_n182));
  aoai13aa1n09x5               g087(.a(new_n182), .b(new_n124), .c(new_n109), .d(new_n117), .o1(new_n183));
  oai012aa1n02x5               g088(.a(new_n154), .b(\b[11] ), .c(\a[12] ), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  and002aa1n02x5               g090(.a(\b[14] ), .b(\a[15] ), .o(new_n186));
  orn002aa1n02x5               g091(.a(\a[16] ), .b(\b[15] ), .o(new_n187));
  aoai13aa1n04x5               g092(.a(new_n187), .b(new_n186), .c(new_n169), .d(new_n173), .o1(new_n188));
  aboi22aa1n09x5               g093(.a(new_n181), .b(new_n184), .c(new_n188), .d(new_n185), .out0(new_n189));
  xorc02aa1n02x5               g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n190), .b(new_n183), .c(new_n189), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(\b[16] ), .b(new_n192), .out0(new_n193));
  nanp02aa1n02x5               g098(.a(new_n188), .b(new_n185), .o1(new_n194));
  tech160nm_fioai012aa1n04x5   g099(.a(new_n194), .b(new_n155), .c(new_n181), .o1(new_n195));
  aoai13aa1n02x5               g100(.a(new_n190), .b(new_n195), .c(new_n139), .d(new_n182), .o1(new_n196));
  xnrc02aa1n02x5               g101(.a(\b[17] ), .b(\a[18] ), .out0(new_n197));
  xobna2aa1n03x5               g102(.a(new_n197), .b(new_n196), .c(new_n193), .out0(\s[18] ));
  inv040aa1d32x5               g103(.a(\a[18] ), .o1(new_n199));
  xroi22aa1d06x4               g104(.a(new_n192), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  oai022aa1n04x7               g106(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n202));
  oaib12aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(\b[17] ), .out0(new_n203));
  aoai13aa1n04x5               g108(.a(new_n203), .b(new_n201), .c(new_n183), .d(new_n189), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand02aa1n06x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nor002aa1n16x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand02aa1d04x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nanb02aa1n02x5               g115(.a(new_n209), .b(new_n210), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n207), .c(new_n204), .d(new_n208), .o1(new_n212));
  aoi112aa1n03x5               g117(.a(new_n207), .b(new_n211), .c(new_n204), .d(new_n208), .o1(new_n213));
  nanb02aa1n03x5               g118(.a(new_n213), .b(new_n212), .out0(\s[20] ));
  nano23aa1n06x5               g119(.a(new_n207), .b(new_n209), .c(new_n210), .d(new_n208), .out0(new_n215));
  nanb03aa1n02x5               g120(.a(new_n197), .b(new_n215), .c(new_n190), .out0(new_n216));
  nona23aa1n09x5               g121(.a(new_n210), .b(new_n208), .c(new_n207), .d(new_n209), .out0(new_n217));
  tech160nm_fiaoi012aa1n04x5   g122(.a(new_n209), .b(new_n207), .c(new_n210), .o1(new_n218));
  oai012aa1n12x5               g123(.a(new_n218), .b(new_n217), .c(new_n203), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n04x5               g125(.a(new_n220), .b(new_n216), .c(new_n183), .d(new_n189), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  xnrc02aa1n12x5               g128(.a(\b[20] ), .b(\a[21] ), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  tech160nm_fixnrc02aa1n05x5   g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n221), .d(new_n225), .o1(new_n227));
  aoi112aa1n03x4               g132(.a(new_n223), .b(new_n226), .c(new_n221), .d(new_n225), .o1(new_n228));
  nanb02aa1n03x5               g133(.a(new_n228), .b(new_n227), .out0(\s[22] ));
  nor042aa1n02x5               g134(.a(new_n226), .b(new_n224), .o1(new_n230));
  nand23aa1n06x5               g135(.a(new_n200), .b(new_n230), .c(new_n215), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\a[22] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\b[21] ), .o1(new_n233));
  oao003aa1n02x5               g138(.a(new_n232), .b(new_n233), .c(new_n223), .carry(new_n234));
  tech160nm_fiaoi012aa1n02p5x5 g139(.a(new_n234), .b(new_n219), .c(new_n230), .o1(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n231), .c(new_n183), .d(new_n189), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  xorc02aa1n02x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xnrc02aa1n02x5               g144(.a(\b[23] ), .b(\a[24] ), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n240), .b(new_n238), .c(new_n236), .d(new_n239), .o1(new_n241));
  aoi112aa1n03x4               g146(.a(new_n238), .b(new_n240), .c(new_n236), .d(new_n239), .o1(new_n242));
  nanb02aa1n03x5               g147(.a(new_n242), .b(new_n241), .out0(\s[24] ));
  norb02aa1n02x5               g148(.a(new_n239), .b(new_n240), .out0(new_n244));
  inv000aa1n02x5               g149(.a(new_n244), .o1(new_n245));
  nano32aa1n03x7               g150(.a(new_n245), .b(new_n200), .c(new_n230), .d(new_n215), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n195), .c(new_n139), .d(new_n182), .o1(new_n247));
  oaoi03aa1n02x5               g152(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n218), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n230), .b(new_n249), .c(new_n215), .d(new_n248), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n234), .o1(new_n251));
  oai022aa1n02x5               g156(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n252));
  aob012aa1n02x5               g157(.a(new_n252), .b(\b[23] ), .c(\a[24] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n245), .c(new_n250), .d(new_n251), .o1(new_n254));
  nanb02aa1n06x5               g159(.a(new_n254), .b(new_n247), .out0(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  tech160nm_fixorc02aa1n04x5   g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  nor002aa1n04x5               g163(.a(\b[25] ), .b(\a[26] ), .o1(new_n259));
  nand42aa1n03x5               g164(.a(\b[25] ), .b(\a[26] ), .o1(new_n260));
  norb02aa1n09x5               g165(.a(new_n260), .b(new_n259), .out0(new_n261));
  inv030aa1n04x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n263));
  nand42aa1n02x5               g168(.a(new_n255), .b(new_n258), .o1(new_n264));
  nona22aa1n02x4               g169(.a(new_n264), .b(new_n262), .c(new_n257), .out0(new_n265));
  nanp02aa1n03x5               g170(.a(new_n265), .b(new_n263), .o1(\s[26] ));
  norb02aa1n09x5               g171(.a(new_n258), .b(new_n262), .out0(new_n267));
  nano22aa1n03x7               g172(.a(new_n231), .b(new_n267), .c(new_n244), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n195), .c(new_n139), .d(new_n182), .o1(new_n269));
  oai012aa1n02x5               g174(.a(new_n260), .b(new_n259), .c(new_n257), .o1(new_n270));
  aobi12aa1n06x5               g175(.a(new_n270), .b(new_n254), .c(new_n267), .out0(new_n271));
  xorc02aa1n12x5               g176(.a(\a[27] ), .b(\b[26] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n269), .out0(\s[27] ));
  nanp02aa1n02x5               g178(.a(new_n254), .b(new_n267), .o1(new_n274));
  nand43aa1n03x5               g179(.a(new_n269), .b(new_n274), .c(new_n270), .o1(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  nor022aa1n06x5               g181(.a(\b[27] ), .b(\a[28] ), .o1(new_n277));
  nanp02aa1n04x5               g182(.a(\b[27] ), .b(\a[28] ), .o1(new_n278));
  nanb02aa1n06x5               g183(.a(new_n277), .b(new_n278), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n275), .d(new_n272), .o1(new_n280));
  aobi12aa1n06x5               g185(.a(new_n268), .b(new_n183), .c(new_n189), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n244), .b(new_n234), .c(new_n219), .d(new_n230), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n267), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n270), .b(new_n283), .c(new_n282), .d(new_n253), .o1(new_n284));
  oaih12aa1n02x5               g189(.a(new_n272), .b(new_n284), .c(new_n281), .o1(new_n285));
  nona22aa1n03x5               g190(.a(new_n285), .b(new_n279), .c(new_n276), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n280), .b(new_n286), .o1(\s[28] ));
  norb02aa1d27x5               g192(.a(new_n272), .b(new_n279), .out0(new_n288));
  oai012aa1n03x5               g193(.a(new_n288), .b(new_n284), .c(new_n281), .o1(new_n289));
  xorc02aa1n02x5               g194(.a(\a[29] ), .b(\b[28] ), .out0(new_n290));
  aoi012aa1n02x5               g195(.a(new_n277), .b(new_n276), .c(new_n278), .o1(new_n291));
  norb02aa1n02x5               g196(.a(new_n291), .b(new_n290), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n288), .o1(new_n293));
  aoai13aa1n02x7               g198(.a(new_n291), .b(new_n293), .c(new_n271), .d(new_n269), .o1(new_n294));
  aoi022aa1n03x5               g199(.a(new_n294), .b(new_n290), .c(new_n289), .d(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g201(.a(new_n279), .b(new_n272), .c(new_n290), .out0(new_n297));
  oai012aa1n03x5               g202(.a(new_n297), .b(new_n284), .c(new_n281), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .out0(new_n299));
  oao003aa1n02x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n300));
  norb02aa1n02x5               g205(.a(new_n300), .b(new_n299), .out0(new_n301));
  inv000aa1n02x5               g206(.a(new_n297), .o1(new_n302));
  aoai13aa1n02x7               g207(.a(new_n300), .b(new_n302), .c(new_n271), .d(new_n269), .o1(new_n303));
  aoi022aa1n03x5               g208(.a(new_n303), .b(new_n299), .c(new_n298), .d(new_n301), .o1(\s[30] ));
  nand03aa1n02x5               g209(.a(new_n288), .b(new_n290), .c(new_n299), .o1(new_n305));
  oabi12aa1n03x5               g210(.a(new_n305), .b(new_n284), .c(new_n281), .out0(new_n306));
  xorc02aa1n02x5               g211(.a(\a[31] ), .b(\b[30] ), .out0(new_n307));
  oao003aa1n02x5               g212(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n308));
  norb02aa1n02x5               g213(.a(new_n308), .b(new_n307), .out0(new_n309));
  aoai13aa1n02x7               g214(.a(new_n308), .b(new_n305), .c(new_n271), .d(new_n269), .o1(new_n310));
  aoi022aa1n03x5               g215(.a(new_n310), .b(new_n307), .c(new_n306), .d(new_n309), .o1(\s[31] ));
  xnrb03aa1n02x5               g216(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g217(.a(\a[3] ), .b(\b[2] ), .c(new_n102), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnrc02aa1n02x5               g219(.a(new_n134), .b(new_n111), .out0(\s[5] ));
  tech160nm_fiaoi012aa1n05x5   g220(.a(new_n122), .b(new_n109), .c(new_n111), .o1(new_n316));
  xnrb03aa1n02x5               g221(.a(new_n316), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaib12aa1n09x5               g222(.a(new_n112), .b(new_n113), .c(new_n316), .out0(new_n318));
  xnbna2aa1n03x5               g223(.a(new_n318), .b(new_n118), .c(new_n121), .out0(\s[7] ));
  inv000aa1d42x5               g224(.a(new_n121), .o1(new_n320));
  norb02aa1n02x5               g225(.a(new_n115), .b(new_n114), .out0(new_n321));
  aoi112aa1n03x5               g226(.a(new_n321), .b(new_n320), .c(new_n318), .d(new_n118), .o1(new_n322));
  aoai13aa1n02x5               g227(.a(new_n321), .b(new_n320), .c(new_n318), .d(new_n118), .o1(new_n323));
  nanb02aa1n02x5               g228(.a(new_n322), .b(new_n323), .out0(\s[8] ));
  xorb03aa1n02x5               g229(.a(new_n139), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


