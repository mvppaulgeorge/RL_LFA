// Benchmark "adder" written by ABC on Wed Jul 17 17:35:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n330, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nand02aa1d06x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nor042aa1n06x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nona23aa1n09x5               g006(.a(new_n101), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n102));
  nor042aa1n04x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nand22aa1n06x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nor042aa1n04x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  nand02aa1n03x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  nor042aa1n03x5               g012(.a(new_n107), .b(new_n102), .o1(new_n108));
  nor042aa1n06x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  inv040aa1n03x5               g014(.a(new_n109), .o1(new_n110));
  oaoi03aa1n06x5               g015(.a(\a[4] ), .b(\b[3] ), .c(new_n110), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nand42aa1n16x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  norp02aa1n06x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[0] ), .b(\a[1] ), .o1(new_n115));
  nand02aa1n03x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  aoi012aa1n06x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  nano32aa1n03x5               g022(.a(new_n117), .b(new_n110), .c(new_n112), .d(new_n113), .out0(new_n118));
  tech160nm_fioai012aa1n02p5x5 g023(.a(new_n108), .b(new_n118), .c(new_n111), .o1(new_n119));
  inv040aa1d32x5               g024(.a(\a[8] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[7] ), .o1(new_n121));
  nand42aa1n02x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(new_n100), .b(new_n99), .o1(new_n123));
  nand02aa1n02x5               g028(.a(new_n122), .b(new_n99), .o1(new_n124));
  nanb02aa1n02x5               g029(.a(new_n100), .b(new_n101), .out0(new_n125));
  tech160nm_fiaoi012aa1n05x5   g030(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n126));
  norp03aa1n02x5               g031(.a(new_n126), .b(new_n125), .c(new_n124), .o1(new_n127));
  nano22aa1n03x7               g032(.a(new_n127), .b(new_n122), .c(new_n123), .out0(new_n128));
  nanp02aa1n02x5               g033(.a(new_n119), .b(new_n128), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  aoi012aa1n02x5               g035(.a(new_n97), .b(new_n129), .c(new_n130), .o1(new_n131));
  xnrb03aa1n02x5               g036(.a(new_n131), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n06x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  nand22aa1n03x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nona23aa1n03x5               g039(.a(new_n130), .b(new_n134), .c(new_n133), .d(new_n97), .out0(new_n135));
  aoi012aa1n02x5               g040(.a(new_n133), .b(new_n97), .c(new_n134), .o1(new_n136));
  aoai13aa1n02x5               g041(.a(new_n136), .b(new_n135), .c(new_n119), .d(new_n128), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand22aa1n09x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  aoi012aa1n02x5               g045(.a(new_n139), .b(new_n137), .c(new_n140), .o1(new_n141));
  nor042aa1d18x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d24x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n15x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  xnrc02aa1n02x5               g049(.a(new_n141), .b(new_n144), .out0(\s[12] ));
  aoi112aa1n09x5               g050(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n146));
  aoi112aa1n09x5               g051(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n147));
  norb02aa1n06x5               g052(.a(new_n140), .b(new_n139), .out0(new_n148));
  oai112aa1n06x5               g053(.a(new_n148), .b(new_n144), .c(new_n147), .d(new_n133), .o1(new_n149));
  nona22aa1d18x5               g054(.a(new_n149), .b(new_n146), .c(new_n142), .out0(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  norb02aa1n02x7               g056(.a(new_n113), .b(new_n109), .out0(new_n152));
  aoi022aa1d24x5               g057(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n153));
  oai112aa1n02x7               g058(.a(new_n152), .b(new_n112), .c(new_n153), .d(new_n114), .o1(new_n154));
  nanb02aa1n06x5               g059(.a(new_n111), .b(new_n154), .out0(new_n155));
  oai112aa1n03x5               g060(.a(new_n122), .b(new_n123), .c(new_n102), .d(new_n126), .o1(new_n156));
  nano22aa1n02x4               g061(.a(new_n135), .b(new_n148), .c(new_n144), .out0(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n156), .c(new_n155), .d(new_n108), .o1(new_n158));
  nanp02aa1n02x5               g063(.a(new_n158), .b(new_n151), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n12x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nand42aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  aoi012aa1n02x5               g067(.a(new_n161), .b(new_n159), .c(new_n162), .o1(new_n163));
  xnrb03aa1n02x5               g068(.a(new_n163), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n04x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nanp02aa1n04x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  tech160nm_fiaoi012aa1n03p5x5 g071(.a(new_n165), .b(new_n161), .c(new_n166), .o1(new_n167));
  nona23aa1n09x5               g072(.a(new_n166), .b(new_n162), .c(new_n161), .d(new_n165), .out0(new_n168));
  aoai13aa1n03x5               g073(.a(new_n167), .b(new_n168), .c(new_n158), .d(new_n151), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand42aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nor042aa1d18x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  aoi122aa1n02x5               g080(.a(new_n171), .b(new_n175), .c(new_n174), .d(new_n169), .e(new_n172), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n177));
  nanb02aa1n06x5               g082(.a(new_n173), .b(new_n175), .out0(new_n178));
  norp02aa1n02x5               g083(.a(new_n177), .b(new_n178), .o1(new_n179));
  norp02aa1n02x5               g084(.a(new_n179), .b(new_n176), .o1(\s[16] ));
  nano23aa1n03x5               g085(.a(new_n133), .b(new_n97), .c(new_n130), .d(new_n134), .out0(new_n181));
  nano23aa1n06x5               g086(.a(new_n139), .b(new_n142), .c(new_n143), .d(new_n140), .out0(new_n182));
  nano23aa1n02x5               g087(.a(new_n161), .b(new_n165), .c(new_n166), .d(new_n162), .out0(new_n183));
  nano23aa1n09x5               g088(.a(new_n171), .b(new_n173), .c(new_n175), .d(new_n172), .out0(new_n184));
  nand02aa1n02x5               g089(.a(new_n184), .b(new_n183), .o1(new_n185));
  nano22aa1n03x7               g090(.a(new_n185), .b(new_n181), .c(new_n182), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n156), .c(new_n155), .d(new_n108), .o1(new_n187));
  nanb02aa1n03x5               g092(.a(new_n171), .b(new_n172), .out0(new_n188));
  nor043aa1n03x5               g093(.a(new_n168), .b(new_n178), .c(new_n188), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n190));
  oai013aa1n03x5               g095(.a(new_n174), .b(new_n167), .c(new_n188), .d(new_n178), .o1(new_n191));
  aoi112aa1n06x5               g096(.a(new_n191), .b(new_n190), .c(new_n150), .d(new_n189), .o1(new_n192));
  nanp02aa1n06x5               g097(.a(new_n192), .b(new_n187), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nona23aa1n09x5               g099(.a(new_n184), .b(new_n182), .c(new_n135), .d(new_n168), .out0(new_n195));
  aoi012aa1n06x5               g100(.a(new_n195), .b(new_n119), .c(new_n128), .o1(new_n196));
  nand42aa1n02x5               g101(.a(new_n150), .b(new_n189), .o1(new_n197));
  nona22aa1n03x5               g102(.a(new_n197), .b(new_n191), .c(new_n190), .out0(new_n198));
  nor002aa1n03x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  nand42aa1n06x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  oaoi13aa1n06x5               g105(.a(new_n199), .b(new_n200), .c(new_n198), .d(new_n196), .o1(new_n201));
  xnrb03aa1n02x5               g106(.a(new_n201), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor042aa1n04x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand42aa1n03x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nano23aa1d12x5               g109(.a(new_n199), .b(new_n203), .c(new_n204), .d(new_n200), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  tech160nm_fiao0012aa1n02p5x5 g111(.a(new_n203), .b(new_n199), .c(new_n204), .o(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  aoai13aa1n03x5               g113(.a(new_n208), .b(new_n206), .c(new_n192), .d(new_n187), .o1(new_n209));
  xorb03aa1n02x5               g114(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n03x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nand22aa1n03x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nor042aa1n04x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand22aa1n03x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  norb02aa1n09x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  aoi112aa1n02x7               g121(.a(new_n212), .b(new_n216), .c(new_n209), .d(new_n213), .o1(new_n217));
  aoai13aa1n03x5               g122(.a(new_n216), .b(new_n212), .c(new_n209), .d(new_n213), .o1(new_n218));
  norb02aa1n03x4               g123(.a(new_n218), .b(new_n217), .out0(\s[20] ));
  nano23aa1n02x5               g124(.a(new_n212), .b(new_n214), .c(new_n215), .d(new_n213), .out0(new_n220));
  nand02aa1n02x5               g125(.a(new_n220), .b(new_n205), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n222));
  aoi112aa1n03x5               g127(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n223));
  norb02aa1n03x5               g128(.a(new_n213), .b(new_n212), .out0(new_n224));
  oai112aa1n06x5               g129(.a(new_n224), .b(new_n216), .c(new_n223), .d(new_n203), .o1(new_n225));
  nona22aa1d18x5               g130(.a(new_n225), .b(new_n222), .c(new_n214), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n221), .c(new_n192), .d(new_n187), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n08x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand42aa1n08x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  nor002aa1n02x5               g137(.a(\b[21] ), .b(\a[22] ), .o1(new_n233));
  nand02aa1n06x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  norb02aa1n06x4               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  aoi112aa1n03x5               g140(.a(new_n230), .b(new_n235), .c(new_n228), .d(new_n232), .o1(new_n236));
  aoai13aa1n06x5               g141(.a(new_n235), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n237));
  norb02aa1n03x4               g142(.a(new_n237), .b(new_n236), .out0(\s[22] ));
  nano23aa1n03x5               g143(.a(new_n230), .b(new_n233), .c(new_n234), .d(new_n231), .out0(new_n239));
  aoi012aa1n03x5               g144(.a(new_n233), .b(new_n230), .c(new_n234), .o1(new_n240));
  aobi12aa1n06x5               g145(.a(new_n240), .b(new_n226), .c(new_n239), .out0(new_n241));
  nand23aa1n03x5               g146(.a(new_n220), .b(new_n205), .c(new_n239), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n241), .b(new_n242), .c(new_n192), .d(new_n187), .o1(new_n243));
  xorb03aa1n02x5               g148(.a(new_n243), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor022aa1n08x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  nand02aa1n04x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  nor022aa1n16x5               g151(.a(\b[23] ), .b(\a[24] ), .o1(new_n247));
  nanp02aa1n04x5               g152(.a(\b[23] ), .b(\a[24] ), .o1(new_n248));
  nanb02aa1n02x5               g153(.a(new_n247), .b(new_n248), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoi112aa1n02x7               g155(.a(new_n245), .b(new_n250), .c(new_n243), .d(new_n246), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n250), .b(new_n245), .c(new_n243), .d(new_n246), .o1(new_n252));
  norb02aa1n03x4               g157(.a(new_n252), .b(new_n251), .out0(\s[24] ));
  nona23aa1d18x5               g158(.a(new_n248), .b(new_n246), .c(new_n245), .d(new_n247), .out0(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  nanb03aa1n03x5               g160(.a(new_n221), .b(new_n255), .c(new_n239), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n247), .o1(new_n257));
  nanp02aa1n02x5               g162(.a(new_n245), .b(new_n248), .o1(new_n258));
  oai112aa1n02x5               g163(.a(new_n258), .b(new_n257), .c(new_n254), .d(new_n240), .o1(new_n259));
  nano22aa1n09x5               g164(.a(new_n254), .b(new_n232), .c(new_n235), .out0(new_n260));
  tech160nm_fiaoi012aa1n02p5x5 g165(.a(new_n259), .b(new_n226), .c(new_n260), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n256), .c(new_n192), .d(new_n187), .o1(new_n262));
  xorb03aa1n02x5               g167(.a(new_n262), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  xorc02aa1n02x5               g169(.a(\a[25] ), .b(\b[24] ), .out0(new_n265));
  xorc02aa1n02x5               g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  aoi112aa1n02x5               g171(.a(new_n264), .b(new_n266), .c(new_n262), .d(new_n265), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n266), .b(new_n264), .c(new_n262), .d(new_n265), .o1(new_n268));
  norb02aa1n03x4               g173(.a(new_n268), .b(new_n267), .out0(\s[26] ));
  nano32aa1n03x7               g174(.a(new_n242), .b(new_n266), .c(new_n255), .d(new_n265), .out0(new_n270));
  oai012aa1n12x5               g175(.a(new_n270), .b(new_n198), .c(new_n196), .o1(new_n271));
  nor002aa1n04x5               g176(.a(\b[25] ), .b(\a[26] ), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n272), .o1(new_n273));
  aoi112aa1n02x7               g178(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nor002aa1n02x5               g180(.a(new_n254), .b(new_n240), .o1(new_n276));
  nano22aa1n03x5               g181(.a(new_n276), .b(new_n257), .c(new_n258), .out0(new_n277));
  nanp02aa1n09x5               g182(.a(new_n226), .b(new_n260), .o1(new_n278));
  and002aa1n02x5               g183(.a(new_n266), .b(new_n265), .o(new_n279));
  aobi12aa1n09x5               g184(.a(new_n279), .b(new_n278), .c(new_n277), .out0(new_n280));
  nano22aa1n12x5               g185(.a(new_n280), .b(new_n273), .c(new_n275), .out0(new_n281));
  xnrc02aa1n12x5               g186(.a(\b[26] ), .b(\a[27] ), .out0(new_n282));
  xobna2aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n271), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  xnrc02aa1n12x5               g190(.a(\b[27] ), .b(\a[28] ), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n279), .b(new_n259), .c(new_n226), .d(new_n260), .o1(new_n287));
  nona22aa1n06x5               g192(.a(new_n287), .b(new_n274), .c(new_n272), .out0(new_n288));
  and002aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n288), .c(new_n193), .d(new_n270), .o1(new_n291));
  aoi012aa1n03x5               g196(.a(new_n286), .b(new_n291), .c(new_n285), .o1(new_n292));
  aoi012aa1n06x5               g197(.a(new_n289), .b(new_n281), .c(new_n271), .o1(new_n293));
  nano22aa1n03x7               g198(.a(new_n293), .b(new_n285), .c(new_n286), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[28] ));
  nor042aa1n03x5               g200(.a(new_n286), .b(new_n282), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n288), .c(new_n193), .d(new_n270), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .out0(new_n299));
  aoi012aa1n03x5               g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n296), .o1(new_n301));
  aoi012aa1n06x5               g206(.a(new_n301), .b(new_n281), .c(new_n271), .o1(new_n302));
  nano22aa1n03x7               g207(.a(new_n302), .b(new_n298), .c(new_n299), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n300), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n115), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nor043aa1n03x5               g210(.a(new_n299), .b(new_n286), .c(new_n282), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n288), .c(new_n193), .d(new_n270), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[29] ), .b(\a[30] ), .out0(new_n309));
  aoi012aa1n02x5               g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n306), .o1(new_n311));
  tech160nm_fiaoi012aa1n04x5   g216(.a(new_n311), .b(new_n281), .c(new_n271), .o1(new_n312));
  nano22aa1n02x4               g217(.a(new_n312), .b(new_n308), .c(new_n309), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n310), .b(new_n313), .o1(\s[30] ));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  norb03aa1n02x5               g220(.a(new_n296), .b(new_n309), .c(new_n299), .out0(new_n316));
  inv020aa1n02x5               g221(.a(new_n316), .o1(new_n317));
  aoi012aa1n06x5               g222(.a(new_n317), .b(new_n281), .c(new_n271), .o1(new_n318));
  oao003aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n319));
  nano22aa1n03x7               g224(.a(new_n318), .b(new_n315), .c(new_n319), .out0(new_n320));
  aoai13aa1n03x5               g225(.a(new_n316), .b(new_n288), .c(new_n193), .d(new_n270), .o1(new_n321));
  aoi012aa1n03x5               g226(.a(new_n315), .b(new_n321), .c(new_n319), .o1(new_n322));
  norp02aa1n03x5               g227(.a(new_n322), .b(new_n320), .o1(\s[31] ));
  xnbna2aa1n03x5               g228(.a(new_n117), .b(new_n110), .c(new_n113), .out0(\s[3] ));
  oaoi13aa1n02x5               g229(.a(new_n109), .b(new_n113), .c(new_n153), .d(new_n114), .o1(new_n325));
  xnrb03aa1n02x5               g230(.a(new_n325), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n155), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi13aa1n02x5               g232(.a(new_n105), .b(new_n106), .c(new_n118), .d(new_n111), .o1(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaib12aa1n02x5               g234(.a(new_n126), .b(new_n107), .c(new_n155), .out0(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g236(.a(new_n100), .b(new_n330), .c(new_n101), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n122), .c(new_n99), .out0(\s[8] ));
  xorb03aa1n02x5               g238(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


