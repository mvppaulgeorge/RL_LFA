// Benchmark "adder" written by ABC on Wed Jul 17 22:59:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n357, new_n358,
    new_n360, new_n362, new_n363, new_n364, new_n366, new_n368, new_n369,
    new_n370, new_n372, new_n373, new_n375, new_n376;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n12x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  nor042aa1n04x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nand02aa1d08x5               g006(.a(\b[8] ), .b(\a[9] ), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nanp02aa1n09x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  norb03aa1d15x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .out0(new_n106));
  inv040aa1d32x5               g011(.a(\a[4] ), .o1(new_n107));
  inv040aa1d28x5               g012(.a(\b[3] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(new_n108), .b(new_n107), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nand42aa1n02x5               g015(.a(new_n109), .b(new_n110), .o1(new_n111));
  nor022aa1n06x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nanb03aa1n06x5               g018(.a(new_n112), .b(new_n113), .c(new_n104), .out0(new_n114));
  nor003aa1n03x5               g019(.a(new_n106), .b(new_n114), .c(new_n111), .o1(new_n115));
  oaoi03aa1n09x5               g020(.a(new_n107), .b(new_n108), .c(new_n112), .o1(new_n116));
  inv000aa1d42x5               g021(.a(new_n116), .o1(new_n117));
  nor002aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1d28x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nor022aa1n16x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nand42aa1n08x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nona23aa1n02x4               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  xnrc02aa1n02x5               g027(.a(\b[5] ), .b(\a[6] ), .out0(new_n123));
  xnrc02aa1n12x5               g028(.a(\b[4] ), .b(\a[5] ), .out0(new_n124));
  nor043aa1n03x5               g029(.a(new_n122), .b(new_n123), .c(new_n124), .o1(new_n125));
  tech160nm_fioai012aa1n05x5   g030(.a(new_n125), .b(new_n115), .c(new_n117), .o1(new_n126));
  nano23aa1n03x5               g031(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n127));
  nor002aa1d32x5               g032(.a(\b[4] ), .b(\a[5] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  oaoi03aa1n03x5               g034(.a(\a[6] ), .b(\b[5] ), .c(new_n129), .o1(new_n130));
  inv000aa1n02x5               g035(.a(new_n120), .o1(new_n131));
  oaoi03aa1n02x5               g036(.a(\a[8] ), .b(\b[7] ), .c(new_n131), .o1(new_n132));
  tech160nm_fiaoi012aa1n04x5   g037(.a(new_n132), .b(new_n127), .c(new_n130), .o1(new_n133));
  nand02aa1n08x5               g038(.a(new_n126), .b(new_n133), .o1(new_n134));
  aoai13aa1n02x5               g039(.a(new_n100), .b(new_n101), .c(new_n134), .d(new_n102), .o1(new_n135));
  oai013aa1n06x5               g040(.a(new_n116), .b(new_n106), .c(new_n114), .d(new_n111), .o1(new_n136));
  inv040aa1n03x5               g041(.a(new_n133), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n102), .b(new_n137), .c(new_n136), .d(new_n125), .o1(new_n138));
  nona22aa1n02x4               g043(.a(new_n138), .b(new_n101), .c(new_n100), .out0(new_n139));
  nanp02aa1n02x5               g044(.a(new_n135), .b(new_n139), .o1(\s[10] ));
  nand42aa1n20x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nor002aa1d32x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nano22aa1n02x4               g047(.a(new_n142), .b(new_n98), .c(new_n141), .out0(new_n143));
  nanp02aa1n03x5               g048(.a(new_n139), .b(new_n143), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n142), .o1(new_n145));
  aoi022aa1n02x5               g050(.a(new_n139), .b(new_n98), .c(new_n145), .d(new_n141), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n144), .b(new_n146), .out0(\s[11] ));
  nor022aa1n16x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nand42aa1d28x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  nona23aa1n02x4               g055(.a(new_n144), .b(new_n149), .c(new_n148), .d(new_n142), .out0(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n150), .c(new_n145), .d(new_n144), .o1(\s[12] ));
  nano23aa1n09x5               g057(.a(new_n148), .b(new_n142), .c(new_n149), .d(new_n141), .out0(new_n153));
  norb02aa1n12x5               g058(.a(new_n102), .b(new_n101), .out0(new_n154));
  nand23aa1d12x5               g059(.a(new_n153), .b(new_n99), .c(new_n154), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nona23aa1n09x5               g061(.a(new_n141), .b(new_n149), .c(new_n148), .d(new_n142), .out0(new_n157));
  tech160nm_fiaoi012aa1n05x5   g062(.a(new_n97), .b(new_n101), .c(new_n98), .o1(new_n158));
  aoi012aa1d18x5               g063(.a(new_n148), .b(new_n142), .c(new_n149), .o1(new_n159));
  tech160nm_fioai012aa1n04x5   g064(.a(new_n159), .b(new_n157), .c(new_n158), .o1(new_n160));
  xnrc02aa1n12x5               g065(.a(\b[12] ), .b(\a[13] ), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n160), .c(new_n134), .d(new_n156), .o1(new_n163));
  oai112aa1n02x5               g068(.a(new_n159), .b(new_n161), .c(new_n157), .d(new_n158), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n164), .b(new_n134), .c(new_n156), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n163), .b(new_n165), .out0(\s[13] ));
  oai012aa1n02x5               g071(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .o1(new_n167));
  xnrc02aa1n02x5               g072(.a(\b[13] ), .b(\a[14] ), .out0(new_n168));
  inv000aa1d42x5               g073(.a(\a[14] ), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\b[13] ), .o1(new_n170));
  nor002aa1n02x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  aoi012aa1n02x5               g076(.a(new_n171), .b(new_n169), .c(new_n170), .o1(new_n172));
  oai112aa1n02x5               g077(.a(new_n163), .b(new_n172), .c(new_n170), .d(new_n169), .o1(new_n173));
  aob012aa1n02x5               g078(.a(new_n173), .b(new_n167), .c(new_n168), .out0(\s[14] ));
  nona32aa1n02x4               g079(.a(new_n134), .b(new_n168), .c(new_n161), .d(new_n155), .out0(new_n175));
  inv000aa1n03x5               g080(.a(new_n158), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n159), .o1(new_n177));
  nor042aa1n06x5               g082(.a(new_n168), .b(new_n161), .o1(new_n178));
  aoai13aa1n04x5               g083(.a(new_n178), .b(new_n177), .c(new_n153), .d(new_n176), .o1(new_n179));
  oaoi03aa1n06x5               g084(.a(new_n169), .b(new_n170), .c(new_n171), .o1(new_n180));
  nanp02aa1n02x5               g085(.a(new_n179), .b(new_n180), .o1(new_n181));
  inv020aa1n02x5               g086(.a(new_n181), .o1(new_n182));
  xnrc02aa1n12x5               g087(.a(\b[14] ), .b(\a[15] ), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  aob012aa1n03x5               g089(.a(new_n184), .b(new_n175), .c(new_n182), .out0(new_n185));
  inv000aa1n02x5               g090(.a(new_n180), .o1(new_n186));
  aoi112aa1n02x5               g091(.a(new_n184), .b(new_n186), .c(new_n160), .d(new_n178), .o1(new_n187));
  aobi12aa1n02x7               g092(.a(new_n185), .b(new_n187), .c(new_n175), .out0(\s[15] ));
  nor042aa1n04x5               g093(.a(\b[14] ), .b(\a[15] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  xnrc02aa1n12x5               g095(.a(\b[15] ), .b(\a[16] ), .out0(new_n191));
  inv000aa1d42x5               g096(.a(new_n191), .o1(new_n192));
  norp02aa1n02x5               g097(.a(\b[15] ), .b(\a[16] ), .o1(new_n193));
  and002aa1n02x5               g098(.a(\b[15] ), .b(\a[16] ), .o(new_n194));
  norp03aa1n02x5               g099(.a(new_n194), .b(new_n193), .c(new_n189), .o1(new_n195));
  aoai13aa1n02x5               g100(.a(new_n195), .b(new_n183), .c(new_n175), .d(new_n182), .o1(new_n196));
  aoai13aa1n02x5               g101(.a(new_n196), .b(new_n192), .c(new_n185), .d(new_n190), .o1(\s[16] ));
  nor042aa1d18x5               g102(.a(new_n191), .b(new_n183), .o1(new_n198));
  nano22aa1d15x5               g103(.a(new_n155), .b(new_n178), .c(new_n198), .out0(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n137), .c(new_n136), .d(new_n125), .o1(new_n200));
  aoai13aa1n06x5               g105(.a(new_n198), .b(new_n186), .c(new_n160), .d(new_n178), .o1(new_n201));
  oab012aa1n09x5               g106(.a(new_n193), .b(new_n190), .c(new_n194), .out0(new_n202));
  nand23aa1d12x5               g107(.a(new_n200), .b(new_n201), .c(new_n202), .o1(new_n203));
  tech160nm_fixorc02aa1n05x5   g108(.a(\a[17] ), .b(\b[16] ), .out0(new_n204));
  nano22aa1n02x4               g109(.a(new_n204), .b(new_n201), .c(new_n202), .out0(new_n205));
  aoi022aa1n02x5               g110(.a(new_n205), .b(new_n200), .c(new_n203), .d(new_n204), .o1(\s[17] ));
  nor042aa1n06x5               g111(.a(\b[16] ), .b(\a[17] ), .o1(new_n207));
  aoi012aa1n02x5               g112(.a(new_n207), .b(new_n203), .c(new_n204), .o1(new_n208));
  nor042aa1n04x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nand02aa1d08x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  norb02aa1n06x4               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  norb03aa1n02x5               g116(.a(new_n210), .b(new_n207), .c(new_n209), .out0(new_n212));
  aob012aa1n02x5               g117(.a(new_n212), .b(new_n203), .c(new_n204), .out0(new_n213));
  oai012aa1n02x5               g118(.a(new_n213), .b(new_n208), .c(new_n211), .o1(\s[18] ));
  inv000aa1d42x5               g119(.a(new_n198), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n202), .b(new_n215), .c(new_n179), .d(new_n180), .o1(new_n216));
  and002aa1n02x5               g121(.a(new_n204), .b(new_n211), .o(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n216), .c(new_n134), .d(new_n199), .o1(new_n218));
  aoi012aa1d24x5               g123(.a(new_n209), .b(new_n207), .c(new_n210), .o1(new_n219));
  nor042aa1d18x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nand02aa1d04x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n218), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g129(.a(new_n220), .o1(new_n225));
  inv020aa1n06x5               g130(.a(new_n219), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n222), .b(new_n226), .c(new_n203), .d(new_n217), .o1(new_n227));
  nor042aa1n04x5               g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  nand02aa1d06x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  inv000aa1n02x5               g135(.a(new_n222), .o1(new_n231));
  norb03aa1n02x5               g136(.a(new_n229), .b(new_n220), .c(new_n228), .out0(new_n232));
  aoai13aa1n02x5               g137(.a(new_n232), .b(new_n231), .c(new_n218), .d(new_n219), .o1(new_n233));
  aoai13aa1n03x5               g138(.a(new_n233), .b(new_n230), .c(new_n227), .d(new_n225), .o1(\s[20] ));
  nona23aa1d18x5               g139(.a(new_n229), .b(new_n221), .c(new_n220), .d(new_n228), .out0(new_n235));
  nano22aa1n03x7               g140(.a(new_n235), .b(new_n204), .c(new_n211), .out0(new_n236));
  aoai13aa1n04x5               g141(.a(new_n236), .b(new_n216), .c(new_n134), .d(new_n199), .o1(new_n237));
  aoi012aa1n12x5               g142(.a(new_n228), .b(new_n220), .c(new_n229), .o1(new_n238));
  oai012aa1d24x5               g143(.a(new_n238), .b(new_n235), .c(new_n219), .o1(new_n239));
  nor042aa1n12x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  nanp02aa1n02x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n239), .c(new_n203), .d(new_n236), .o1(new_n243));
  nano23aa1n06x5               g148(.a(new_n220), .b(new_n228), .c(new_n229), .d(new_n221), .out0(new_n244));
  inv000aa1n06x5               g149(.a(new_n238), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n245), .b(new_n242), .c(new_n244), .d(new_n226), .o1(new_n246));
  aobi12aa1n02x7               g151(.a(new_n243), .b(new_n246), .c(new_n237), .out0(\s[21] ));
  inv000aa1d42x5               g152(.a(new_n240), .o1(new_n248));
  nor042aa1n03x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  and002aa1n06x5               g154(.a(\b[21] ), .b(\a[22] ), .o(new_n250));
  norp02aa1n02x5               g155(.a(new_n250), .b(new_n249), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n239), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n242), .o1(new_n253));
  norp03aa1n02x5               g158(.a(new_n250), .b(new_n249), .c(new_n240), .o1(new_n254));
  aoai13aa1n02x7               g159(.a(new_n254), .b(new_n253), .c(new_n237), .d(new_n252), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n251), .c(new_n243), .d(new_n248), .o1(\s[22] ));
  nano23aa1n09x5               g161(.a(new_n250), .b(new_n249), .c(new_n248), .d(new_n241), .out0(new_n257));
  nano32aa1n02x4               g162(.a(new_n235), .b(new_n257), .c(new_n204), .d(new_n211), .out0(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n216), .c(new_n134), .d(new_n199), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n257), .b(new_n245), .c(new_n244), .d(new_n226), .o1(new_n260));
  oab012aa1d15x5               g165(.a(new_n249), .b(new_n248), .c(new_n250), .out0(new_n261));
  nand42aa1n02x5               g166(.a(new_n260), .b(new_n261), .o1(new_n262));
  xorc02aa1n12x5               g167(.a(\a[23] ), .b(\b[22] ), .out0(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n203), .d(new_n258), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n261), .o1(new_n265));
  aoi112aa1n02x5               g170(.a(new_n263), .b(new_n265), .c(new_n239), .d(new_n257), .o1(new_n266));
  aobi12aa1n02x5               g171(.a(new_n264), .b(new_n266), .c(new_n259), .out0(\s[23] ));
  nor042aa1n03x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  nor002aa1n02x5               g174(.a(\b[23] ), .b(\a[24] ), .o1(new_n270));
  and002aa1n02x5               g175(.a(\b[23] ), .b(\a[24] ), .o(new_n271));
  norp02aa1n03x5               g176(.a(new_n271), .b(new_n270), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n262), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n263), .o1(new_n274));
  norp03aa1n02x5               g179(.a(new_n271), .b(new_n270), .c(new_n268), .o1(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n274), .c(new_n259), .d(new_n273), .o1(new_n276));
  aoai13aa1n02x5               g181(.a(new_n276), .b(new_n272), .c(new_n264), .d(new_n269), .o1(\s[24] ));
  inv000aa1n02x5               g182(.a(new_n236), .o1(new_n278));
  and002aa1n06x5               g183(.a(new_n263), .b(new_n272), .o(new_n279));
  nano22aa1n02x5               g184(.a(new_n278), .b(new_n257), .c(new_n279), .out0(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n216), .c(new_n134), .d(new_n199), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n279), .o1(new_n282));
  oab012aa1n06x5               g187(.a(new_n270), .b(new_n269), .c(new_n271), .out0(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n282), .c(new_n260), .d(new_n261), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n284), .c(new_n203), .d(new_n280), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n279), .b(new_n265), .c(new_n239), .d(new_n257), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  and003aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n283), .o(new_n289));
  aobi12aa1n02x5               g194(.a(new_n286), .b(new_n289), .c(new_n281), .out0(\s[25] ));
  nor042aa1n03x5               g195(.a(\b[24] ), .b(\a[25] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  norp02aa1n02x5               g197(.a(\b[25] ), .b(\a[26] ), .o1(new_n293));
  and002aa1n02x7               g198(.a(\b[25] ), .b(\a[26] ), .o(new_n294));
  nor002aa1n02x5               g199(.a(new_n294), .b(new_n293), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n284), .o1(new_n296));
  norp03aa1n02x5               g201(.a(new_n294), .b(new_n293), .c(new_n291), .o1(new_n297));
  aoai13aa1n04x5               g202(.a(new_n297), .b(new_n288), .c(new_n281), .d(new_n296), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n295), .c(new_n286), .d(new_n292), .o1(\s[26] ));
  and002aa1n06x5               g204(.a(new_n285), .b(new_n295), .o(new_n300));
  nano32aa1n06x5               g205(.a(new_n278), .b(new_n300), .c(new_n257), .d(new_n279), .out0(new_n301));
  aoai13aa1n06x5               g206(.a(new_n301), .b(new_n216), .c(new_n134), .d(new_n199), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n300), .o1(new_n303));
  oab012aa1n04x5               g208(.a(new_n293), .b(new_n292), .c(new_n294), .out0(new_n304));
  aoai13aa1n04x5               g209(.a(new_n304), .b(new_n303), .c(new_n287), .d(new_n283), .o1(new_n305));
  xorc02aa1n12x5               g210(.a(\a[27] ), .b(\b[26] ), .out0(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n305), .c(new_n203), .d(new_n301), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n304), .o1(new_n308));
  aoi112aa1n02x5               g213(.a(new_n306), .b(new_n308), .c(new_n284), .d(new_n300), .o1(new_n309));
  aobi12aa1n03x7               g214(.a(new_n307), .b(new_n309), .c(new_n302), .out0(\s[27] ));
  norp02aa1n02x5               g215(.a(\b[26] ), .b(\a[27] ), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n311), .o1(new_n312));
  norp02aa1n02x5               g217(.a(\b[27] ), .b(\a[28] ), .o1(new_n313));
  and002aa1n03x5               g218(.a(\b[27] ), .b(\a[28] ), .o(new_n314));
  nor002aa1n02x5               g219(.a(new_n314), .b(new_n313), .o1(new_n315));
  aoi012aa1n09x5               g220(.a(new_n308), .b(new_n284), .c(new_n300), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n306), .o1(new_n317));
  norp03aa1n02x5               g222(.a(new_n314), .b(new_n313), .c(new_n311), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n302), .d(new_n316), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n315), .c(new_n307), .d(new_n312), .o1(\s[28] ));
  inv000aa1d42x5               g225(.a(\a[27] ), .o1(new_n321));
  inv000aa1d42x5               g226(.a(\a[28] ), .o1(new_n322));
  xroi22aa1d04x5               g227(.a(new_n321), .b(\b[26] ), .c(new_n322), .d(\b[27] ), .out0(new_n323));
  aoai13aa1n02x5               g228(.a(new_n323), .b(new_n305), .c(new_n203), .d(new_n301), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  aoi112aa1n09x5               g230(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n326));
  oai022aa1n02x5               g231(.a(\a[28] ), .b(\b[27] ), .c(\b[28] ), .d(\a[29] ), .o1(new_n327));
  aoi112aa1n02x5               g232(.a(new_n326), .b(new_n327), .c(\a[29] ), .d(\b[28] ), .o1(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n325), .c(new_n302), .d(new_n316), .o1(new_n329));
  nor042aa1n03x5               g234(.a(new_n326), .b(new_n313), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[29] ), .b(\b[28] ), .out0(new_n331));
  aoai13aa1n03x5               g236(.a(new_n329), .b(new_n331), .c(new_n324), .d(new_n330), .o1(\s[29] ));
  xorb03aa1n02x5               g237(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g238(.a(new_n317), .b(new_n331), .c(new_n315), .out0(new_n334));
  aoai13aa1n02x5               g239(.a(new_n334), .b(new_n305), .c(new_n203), .d(new_n301), .o1(new_n335));
  tech160nm_fioaoi03aa1n03p5x5 g240(.a(\a[29] ), .b(\b[28] ), .c(new_n330), .o1(new_n336));
  inv000aa1d42x5               g241(.a(new_n336), .o1(new_n337));
  norp02aa1n02x5               g242(.a(\b[29] ), .b(\a[30] ), .o1(new_n338));
  nand42aa1n02x5               g243(.a(\b[29] ), .b(\a[30] ), .o1(new_n339));
  norb02aa1n02x5               g244(.a(new_n339), .b(new_n338), .out0(new_n340));
  inv000aa1d42x5               g245(.a(new_n334), .o1(new_n341));
  inv000aa1d42x5               g246(.a(\a[29] ), .o1(new_n342));
  obai22aa1n02x7               g247(.a(\b[28] ), .b(new_n342), .c(new_n326), .d(new_n313), .out0(new_n343));
  oai022aa1n02x5               g248(.a(\a[29] ), .b(\b[28] ), .c(\b[29] ), .d(\a[30] ), .o1(new_n344));
  nano22aa1n02x4               g249(.a(new_n344), .b(new_n343), .c(new_n339), .out0(new_n345));
  aoai13aa1n03x5               g250(.a(new_n345), .b(new_n341), .c(new_n302), .d(new_n316), .o1(new_n346));
  aoai13aa1n03x5               g251(.a(new_n346), .b(new_n340), .c(new_n335), .d(new_n337), .o1(\s[30] ));
  nano32aa1n03x7               g252(.a(new_n317), .b(new_n340), .c(new_n315), .d(new_n331), .out0(new_n348));
  aoai13aa1n02x7               g253(.a(new_n348), .b(new_n305), .c(new_n203), .d(new_n301), .o1(new_n349));
  xnrc02aa1n02x5               g254(.a(\b[30] ), .b(\a[31] ), .out0(new_n350));
  inv000aa1d42x5               g255(.a(new_n350), .o1(new_n351));
  inv000aa1d42x5               g256(.a(new_n348), .o1(new_n352));
  aoi112aa1n03x5               g257(.a(new_n338), .b(new_n350), .c(new_n336), .d(new_n340), .o1(new_n353));
  aoai13aa1n03x5               g258(.a(new_n353), .b(new_n352), .c(new_n302), .d(new_n316), .o1(new_n354));
  aoi012aa1n02x5               g259(.a(new_n338), .b(new_n336), .c(new_n340), .o1(new_n355));
  aoai13aa1n03x5               g260(.a(new_n354), .b(new_n351), .c(new_n349), .d(new_n355), .o1(\s[31] ));
  inv000aa1d42x5               g261(.a(new_n106), .o1(new_n357));
  nanb02aa1n02x5               g262(.a(new_n112), .b(new_n113), .out0(new_n358));
  xnbna2aa1n03x5               g263(.a(new_n358), .b(new_n357), .c(new_n104), .out0(\s[3] ));
  tech160nm_fiao0012aa1n02p5x5 g264(.a(new_n358), .b(new_n357), .c(new_n104), .o(new_n360));
  xnbna2aa1n03x5               g265(.a(new_n111), .b(new_n360), .c(new_n113), .out0(\s[4] ));
  inv000aa1d42x5               g266(.a(new_n124), .o1(new_n362));
  and003aa1n02x5               g267(.a(new_n109), .b(new_n112), .c(new_n110), .o(new_n363));
  nano22aa1n02x4               g268(.a(new_n363), .b(new_n124), .c(new_n109), .out0(new_n364));
  aboi22aa1n03x5               g269(.a(new_n115), .b(new_n364), .c(new_n136), .d(new_n362), .out0(\s[5] ));
  oai012aa1n02x5               g270(.a(new_n362), .b(new_n115), .c(new_n117), .o1(new_n366));
  xobna2aa1n03x5               g271(.a(new_n123), .b(new_n366), .c(new_n129), .out0(\s[6] ));
  nanb02aa1n02x5               g272(.a(new_n120), .b(new_n121), .out0(new_n368));
  nanp02aa1n02x5               g273(.a(\b[5] ), .b(\a[6] ), .o1(new_n369));
  nona22aa1n02x4               g274(.a(new_n366), .b(new_n128), .c(new_n123), .out0(new_n370));
  xnbna2aa1n03x5               g275(.a(new_n368), .b(new_n370), .c(new_n369), .out0(\s[7] ));
  norb02aa1n02x5               g276(.a(new_n119), .b(new_n118), .out0(new_n372));
  nanb03aa1n02x5               g277(.a(new_n368), .b(new_n370), .c(new_n369), .out0(new_n373));
  xnbna2aa1n03x5               g278(.a(new_n372), .b(new_n373), .c(new_n131), .out0(\s[8] ));
  inv000aa1d42x5               g279(.a(new_n154), .o1(new_n375));
  aoi112aa1n02x5               g280(.a(new_n375), .b(new_n132), .c(new_n127), .d(new_n130), .o1(new_n376));
  ao0022aa1n03x5               g281(.a(new_n134), .b(new_n375), .c(new_n376), .d(new_n126), .o(\s[9] ));
endmodule


