// Benchmark "adder" written by ABC on Wed Jul 17 17:55:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n315, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n340, new_n341, new_n343, new_n345, new_n347, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor022aa1n16x5               g002(.a(\b[2] ), .b(\a[3] ), .o1(new_n98));
  norp02aa1n02x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  techfinor002aa1n02p5x5       g004(.a(new_n99), .b(new_n98), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nanb02aa1n06x5               g006(.a(new_n98), .b(new_n101), .out0(new_n102));
  nanp02aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oai112aa1n06x5               g008(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n104));
  nand22aa1n03x5               g009(.a(new_n104), .b(new_n103), .o1(new_n105));
  oai012aa1n12x5               g010(.a(new_n100), .b(new_n105), .c(new_n102), .o1(new_n106));
  nand42aa1n06x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nand02aa1n06x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nanb03aa1n06x5               g014(.a(new_n109), .b(new_n107), .c(new_n108), .out0(new_n110));
  aoi022aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n111));
  inv000aa1d42x5               g016(.a(\a[8] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[7] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  aoi012aa1n02x5               g019(.a(new_n114), .b(new_n112), .c(new_n113), .o1(new_n115));
  inv040aa1d32x5               g020(.a(\a[7] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[6] ), .o1(new_n117));
  nanp02aa1n04x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  nand42aa1n06x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n118), .b(new_n119), .o1(new_n120));
  nano23aa1n06x5               g025(.a(new_n110), .b(new_n120), .c(new_n115), .d(new_n111), .out0(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n106), .o1(new_n122));
  nand42aa1n06x5               g027(.a(new_n113), .b(new_n112), .o1(new_n123));
  nand42aa1n20x5               g028(.a(\b[5] ), .b(\a[6] ), .o1(new_n124));
  oai012aa1n18x5               g029(.a(new_n124), .b(new_n114), .c(new_n109), .o1(new_n125));
  aob012aa1n12x5               g030(.a(new_n119), .b(\b[7] ), .c(\a[8] ), .out0(new_n126));
  aoai13aa1n12x5               g031(.a(new_n123), .b(new_n126), .c(new_n125), .d(new_n118), .o1(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  nanp02aa1n03x5               g033(.a(new_n122), .b(new_n128), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  xnrc02aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n97), .c(new_n129), .d(new_n130), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n130), .o1(new_n133));
  nor042aa1n06x5               g038(.a(new_n131), .b(new_n97), .o1(new_n134));
  aoai13aa1n02x5               g039(.a(new_n134), .b(new_n133), .c(new_n122), .d(new_n128), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(new_n132), .b(new_n135), .o1(\s[10] ));
  nona22aa1n02x4               g041(.a(new_n129), .b(new_n133), .c(new_n131), .out0(new_n137));
  nand02aa1n06x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  oai012aa1n02x5               g043(.a(new_n138), .b(new_n131), .c(new_n97), .o1(new_n139));
  xorc02aa1n02x5               g044(.a(\a[11] ), .b(\b[10] ), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n137), .c(new_n139), .out0(\s[11] ));
  nor042aa1n09x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  inv000aa1n02x5               g047(.a(new_n142), .o1(new_n143));
  aob012aa1n03x5               g048(.a(new_n140), .b(new_n137), .c(new_n139), .out0(new_n144));
  xorc02aa1n02x5               g049(.a(\a[12] ), .b(\b[11] ), .out0(new_n145));
  nand02aa1d24x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  inv020aa1n04x5               g051(.a(new_n146), .o1(new_n147));
  oaih22aa1n04x5               g052(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n148));
  nona22aa1n02x4               g053(.a(new_n144), .b(new_n147), .c(new_n148), .out0(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n145), .c(new_n143), .d(new_n144), .o1(\s[12] ));
  inv040aa1d32x5               g055(.a(\a[12] ), .o1(new_n151));
  inv000aa1d42x5               g056(.a(\b[11] ), .o1(new_n152));
  aoi022aa1d24x5               g057(.a(new_n152), .b(new_n151), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  nona23aa1d18x5               g058(.a(new_n153), .b(new_n138), .c(new_n147), .d(new_n142), .out0(new_n154));
  nor043aa1d12x5               g059(.a(new_n154), .b(new_n133), .c(new_n131), .o1(new_n155));
  aoai13aa1n12x5               g060(.a(new_n155), .b(new_n127), .c(new_n121), .d(new_n106), .o1(new_n156));
  tech160nm_finand02aa1n03p5x5 g061(.a(new_n148), .b(new_n146), .o1(new_n157));
  oaih12aa1n12x5               g062(.a(new_n157), .b(new_n134), .c(new_n154), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  xorc02aa1n12x5               g064(.a(\a[13] ), .b(\b[12] ), .out0(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n156), .c(new_n159), .out0(\s[13] ));
  inv000aa1d42x5               g066(.a(\a[13] ), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(\b[12] ), .b(new_n162), .out0(new_n163));
  nanp02aa1n03x5               g068(.a(new_n156), .b(new_n159), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(new_n164), .b(new_n160), .o1(new_n165));
  tech160nm_fixorc02aa1n05x5   g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n165), .c(new_n163), .out0(\s[14] ));
  nanp02aa1n02x5               g072(.a(new_n166), .b(new_n160), .o1(new_n168));
  inv000aa1d42x5               g073(.a(\a[14] ), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\b[13] ), .o1(new_n170));
  nor002aa1n03x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  tech160nm_fioaoi03aa1n03p5x5 g076(.a(new_n169), .b(new_n170), .c(new_n171), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n168), .c(new_n156), .d(new_n159), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  xorc02aa1n12x5               g079(.a(\a[16] ), .b(\b[15] ), .out0(new_n175));
  norp02aa1n02x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  tech160nm_fixorc02aa1n04x5   g081(.a(\a[15] ), .b(\b[14] ), .out0(new_n177));
  tech160nm_fiaoi012aa1n02p5x5 g082(.a(new_n176), .b(new_n173), .c(new_n177), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n175), .b(new_n176), .out0(new_n179));
  aob012aa1n03x5               g084(.a(new_n179), .b(new_n173), .c(new_n177), .out0(new_n180));
  oai012aa1n03x5               g085(.a(new_n180), .b(new_n178), .c(new_n175), .o1(\s[16] ));
  xroi22aa1d06x4               g086(.a(new_n162), .b(\b[12] ), .c(new_n169), .d(\b[13] ), .out0(new_n182));
  nand23aa1n04x5               g087(.a(new_n182), .b(new_n177), .c(new_n175), .o1(new_n183));
  nano22aa1n03x7               g088(.a(new_n168), .b(new_n177), .c(new_n175), .out0(new_n184));
  inv000aa1d42x5               g089(.a(\a[16] ), .o1(new_n185));
  inv020aa1n02x5               g090(.a(new_n176), .o1(new_n186));
  nanp02aa1n03x5               g091(.a(new_n172), .b(new_n186), .o1(new_n187));
  aoi022aa1n02x5               g092(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(new_n187), .b(new_n188), .o1(new_n189));
  oaib12aa1n02x5               g094(.a(new_n189), .b(\b[15] ), .c(new_n185), .out0(new_n190));
  aoi012aa1n06x5               g095(.a(new_n190), .b(new_n158), .c(new_n184), .o1(new_n191));
  oai012aa1n18x5               g096(.a(new_n191), .b(new_n156), .c(new_n183), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g098(.a(\a[17] ), .o1(new_n194));
  inv040aa1d28x5               g099(.a(\b[16] ), .o1(new_n195));
  nand22aa1n04x5               g100(.a(new_n195), .b(new_n194), .o1(new_n196));
  inv000aa1n02x5               g101(.a(new_n153), .o1(new_n197));
  nano32aa1n03x7               g102(.a(new_n197), .b(new_n143), .c(new_n146), .d(new_n138), .out0(new_n198));
  oai012aa1n02x5               g103(.a(new_n198), .b(new_n131), .c(new_n97), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\b[15] ), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n187), .b(new_n188), .c(new_n200), .d(new_n185), .o1(new_n201));
  aoai13aa1n04x5               g106(.a(new_n201), .b(new_n183), .c(new_n199), .d(new_n157), .o1(new_n202));
  aoi012aa1n06x5               g107(.a(new_n127), .b(new_n121), .c(new_n106), .o1(new_n203));
  nano22aa1n03x7               g108(.a(new_n203), .b(new_n155), .c(new_n184), .out0(new_n204));
  oai022aa1n02x5               g109(.a(new_n204), .b(new_n202), .c(new_n195), .d(new_n194), .o1(new_n205));
  tech160nm_finor002aa1n05x5   g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand22aa1n06x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  norb02aa1n02x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n205), .c(new_n196), .out0(\s[18] ));
  nanp02aa1n02x5               g114(.a(\b[16] ), .b(\a[17] ), .o1(new_n210));
  nano32aa1n03x7               g115(.a(new_n206), .b(new_n196), .c(new_n207), .d(new_n210), .out0(new_n211));
  oaoi03aa1n09x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n196), .o1(new_n212));
  nor002aa1d32x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand02aa1n10x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n212), .c(new_n192), .d(new_n211), .o1(new_n216));
  aoi112aa1n02x7               g121(.a(new_n215), .b(new_n212), .c(new_n192), .d(new_n211), .o1(new_n217));
  norb02aa1n03x4               g122(.a(new_n216), .b(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n06x5               g124(.a(new_n213), .o1(new_n220));
  nor002aa1d32x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand02aa1n08x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  norb03aa1n02x5               g128(.a(new_n222), .b(new_n213), .c(new_n221), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n216), .b(new_n224), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n225), .b(new_n223), .c(new_n216), .d(new_n220), .o1(\s[20] ));
  nano23aa1n09x5               g131(.a(new_n213), .b(new_n221), .c(new_n222), .d(new_n214), .out0(new_n227));
  nanp02aa1n02x5               g132(.a(new_n211), .b(new_n227), .o1(new_n228));
  oabi12aa1n02x5               g133(.a(new_n228), .b(new_n204), .c(new_n202), .out0(new_n229));
  nona22aa1n02x4               g134(.a(new_n198), .b(new_n133), .c(new_n131), .out0(new_n230));
  nona22aa1n02x4               g135(.a(new_n129), .b(new_n230), .c(new_n183), .out0(new_n231));
  aoi013aa1n06x4               g136(.a(new_n206), .b(new_n207), .c(new_n194), .d(new_n195), .o1(new_n232));
  nona23aa1n09x5               g137(.a(new_n222), .b(new_n214), .c(new_n213), .d(new_n221), .out0(new_n233));
  oaoi03aa1n09x5               g138(.a(\a[20] ), .b(\b[19] ), .c(new_n220), .o1(new_n234));
  oabi12aa1n18x5               g139(.a(new_n234), .b(new_n233), .c(new_n232), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n228), .c(new_n231), .d(new_n191), .o1(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[20] ), .b(\a[21] ), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoi112aa1n02x5               g144(.a(new_n234), .b(new_n239), .c(new_n227), .d(new_n212), .o1(new_n240));
  aoi022aa1n02x5               g145(.a(new_n237), .b(new_n239), .c(new_n229), .d(new_n240), .o1(\s[21] ));
  nor042aa1d18x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  aoai13aa1n02x5               g148(.a(new_n243), .b(new_n242), .c(new_n237), .d(new_n239), .o1(new_n244));
  norp02aa1n02x5               g149(.a(new_n243), .b(new_n242), .o1(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n238), .c(new_n229), .d(new_n236), .o1(new_n246));
  nanp02aa1n03x5               g151(.a(new_n244), .b(new_n246), .o1(\s[22] ));
  nor042aa1n06x5               g152(.a(new_n243), .b(new_n238), .o1(new_n248));
  and003aa1n02x5               g153(.a(new_n248), .b(new_n211), .c(new_n227), .o(new_n249));
  tech160nm_fioai012aa1n05x5   g154(.a(new_n249), .b(new_n204), .c(new_n202), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n248), .b(new_n234), .c(new_n227), .d(new_n212), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\a[22] ), .o1(new_n252));
  inv040aa1d32x5               g157(.a(\b[21] ), .o1(new_n253));
  oao003aa1n03x5               g158(.a(new_n252), .b(new_n253), .c(new_n242), .carry(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  nand22aa1n02x5               g160(.a(new_n251), .b(new_n255), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  xnrc02aa1n12x5               g162(.a(\b[22] ), .b(\a[23] ), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n250), .c(new_n257), .out0(\s[23] ));
  norp02aa1n02x5               g165(.a(\b[22] ), .b(\a[23] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n259), .b(new_n256), .c(new_n192), .d(new_n249), .o1(new_n263));
  xorc02aa1n03x5               g168(.a(\a[24] ), .b(\b[23] ), .out0(new_n264));
  nanp02aa1n02x5               g169(.a(\b[23] ), .b(\a[24] ), .o1(new_n265));
  oai022aa1n02x5               g170(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n265), .b(new_n266), .out0(new_n267));
  aoai13aa1n02x5               g172(.a(new_n267), .b(new_n258), .c(new_n250), .d(new_n257), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n264), .c(new_n263), .d(new_n262), .o1(\s[24] ));
  nano32aa1n02x5               g174(.a(new_n228), .b(new_n264), .c(new_n248), .d(new_n259), .out0(new_n270));
  oai012aa1n02x5               g175(.a(new_n270), .b(new_n204), .c(new_n202), .o1(new_n271));
  norb02aa1n09x5               g176(.a(new_n264), .b(new_n258), .out0(new_n272));
  inv020aa1n04x5               g177(.a(new_n272), .o1(new_n273));
  nanp02aa1n02x5               g178(.a(new_n266), .b(new_n265), .o1(new_n274));
  aoai13aa1n12x5               g179(.a(new_n274), .b(new_n273), .c(new_n251), .d(new_n255), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n271), .c(new_n276), .out0(\s[25] ));
  norp02aa1n02x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n277), .b(new_n275), .c(new_n192), .d(new_n270), .o1(new_n281));
  xorc02aa1n03x5               g186(.a(\a[26] ), .b(\b[25] ), .out0(new_n282));
  nanp02aa1n02x5               g187(.a(\b[25] ), .b(\a[26] ), .o1(new_n283));
  oai022aa1n02x5               g188(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n284));
  norb02aa1n02x5               g189(.a(new_n283), .b(new_n284), .out0(new_n285));
  nand42aa1n02x5               g190(.a(new_n281), .b(new_n285), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n282), .c(new_n281), .d(new_n280), .o1(\s[26] ));
  nor002aa1d32x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  and002aa1n24x5               g193(.a(\b[26] ), .b(\a[27] ), .o(new_n289));
  nor042aa1n03x5               g194(.a(new_n289), .b(new_n288), .o1(new_n290));
  and002aa1n06x5               g195(.a(new_n282), .b(new_n277), .o(new_n291));
  nano32aa1n06x5               g196(.a(new_n228), .b(new_n291), .c(new_n248), .d(new_n272), .out0(new_n292));
  oai012aa1n06x5               g197(.a(new_n292), .b(new_n204), .c(new_n202), .o1(new_n293));
  aoi022aa1n12x5               g198(.a(new_n275), .b(new_n291), .c(new_n283), .d(new_n284), .o1(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n290), .b(new_n294), .c(new_n293), .out0(\s[27] ));
  inv000aa1d42x5               g200(.a(new_n289), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n272), .b(new_n254), .c(new_n235), .d(new_n248), .o1(new_n297));
  inv000aa1n02x5               g202(.a(new_n291), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n284), .b(new_n283), .o1(new_n299));
  aoai13aa1n02x7               g204(.a(new_n299), .b(new_n298), .c(new_n297), .d(new_n274), .o1(new_n300));
  aoai13aa1n02x5               g205(.a(new_n296), .b(new_n300), .c(new_n192), .d(new_n292), .o1(new_n301));
  inv040aa1n08x5               g206(.a(new_n288), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n289), .c(new_n294), .d(new_n293), .o1(new_n303));
  xorc02aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .out0(new_n304));
  norp02aa1n02x5               g209(.a(new_n304), .b(new_n288), .o1(new_n305));
  aoi022aa1n03x5               g210(.a(new_n303), .b(new_n304), .c(new_n301), .d(new_n305), .o1(\s[28] ));
  and002aa1n06x5               g211(.a(new_n304), .b(new_n290), .o(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n300), .c(new_n192), .d(new_n292), .o1(new_n308));
  inv000aa1n02x5               g213(.a(new_n307), .o1(new_n309));
  oao003aa1n03x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n302), .carry(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n309), .c(new_n294), .d(new_n293), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n308), .d(new_n313), .o1(\s[29] ));
  nanp02aa1n02x5               g219(.a(\b[0] ), .b(\a[1] ), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g221(.a(new_n304), .b(new_n312), .c(new_n290), .o(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n300), .c(new_n192), .d(new_n292), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  tech160nm_fioaoi03aa1n03p5x5 g224(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n319), .c(new_n294), .d(new_n293), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(\b[28] ), .b(\a[29] ), .o(new_n324));
  oabi12aa1n02x5               g229(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n325));
  oab012aa1n02x4               g230(.a(new_n325), .b(new_n310), .c(new_n324), .out0(new_n326));
  aoi022aa1n03x5               g231(.a(new_n322), .b(new_n323), .c(new_n318), .d(new_n326), .o1(\s[30] ));
  nano22aa1n09x5               g232(.a(new_n309), .b(new_n312), .c(new_n323), .out0(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n300), .c(new_n192), .d(new_n292), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  inv000aa1d42x5               g235(.a(\a[30] ), .o1(new_n331));
  inv000aa1d42x5               g236(.a(\b[29] ), .o1(new_n332));
  oabi12aa1n02x5               g237(.a(new_n330), .b(\a[30] ), .c(\b[29] ), .out0(new_n333));
  oaoi13aa1n02x5               g238(.a(new_n333), .b(new_n320), .c(new_n331), .d(new_n332), .o1(new_n334));
  inv000aa1d42x5               g239(.a(new_n328), .o1(new_n335));
  oaoi03aa1n03x5               g240(.a(new_n331), .b(new_n332), .c(new_n320), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n335), .c(new_n294), .d(new_n293), .o1(new_n337));
  aoi022aa1n03x5               g242(.a(new_n337), .b(new_n330), .c(new_n329), .d(new_n334), .o1(\s[31] ));
  xnbna2aa1n03x5               g243(.a(new_n102), .b(new_n104), .c(new_n103), .out0(\s[3] ));
  norb02aa1n02x5               g244(.a(new_n107), .b(new_n99), .out0(new_n340));
  aoi113aa1n02x5               g245(.a(new_n98), .b(new_n340), .c(new_n104), .d(new_n103), .e(new_n101), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n341), .b(new_n106), .c(new_n340), .o1(\s[4] ));
  nanb02aa1n02x5               g247(.a(new_n109), .b(new_n108), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n106), .c(new_n107), .out0(\s[5] ));
  aoai13aa1n02x5               g249(.a(new_n108), .b(new_n109), .c(new_n106), .d(new_n107), .o1(new_n345));
  xnrb03aa1n02x5               g250(.a(new_n345), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n03x5               g251(.a(\a[6] ), .b(\b[5] ), .c(new_n345), .o1(new_n347));
  xorb03aa1n02x5               g252(.a(new_n347), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g253(.a(new_n116), .b(new_n117), .c(new_n347), .o1(new_n349));
  xorb03aa1n02x5               g254(.a(new_n349), .b(\b[7] ), .c(new_n112), .out0(\s[8] ));
  xnbna2aa1n03x5               g255(.a(new_n130), .b(new_n122), .c(new_n128), .out0(\s[9] ));
endmodule


