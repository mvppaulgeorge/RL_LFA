// Benchmark "adder" written by ABC on Wed Jul 17 13:24:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n361, new_n362, new_n363, new_n365, new_n366,
    new_n368, new_n369, new_n370, new_n371, new_n373, new_n374, new_n376,
    new_n377, new_n380;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n06x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1n04x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand42aa1d28x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand22aa1n09x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  norb03aa1d15x5               g005(.a(new_n99), .b(new_n98), .c(new_n100), .out0(new_n101));
  nand02aa1d16x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nor002aa1d32x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanb03aa1d24x5               g008(.a(new_n103), .b(new_n99), .c(new_n102), .out0(new_n104));
  oai022aa1d18x5               g009(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n105));
  oabi12aa1n18x5               g010(.a(new_n105), .b(new_n101), .c(new_n104), .out0(new_n106));
  nanp02aa1n04x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nand42aa1n20x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  inv040aa1d32x5               g013(.a(\a[5] ), .o1(new_n109));
  inv040aa1d32x5               g014(.a(\b[4] ), .o1(new_n110));
  nand02aa1n10x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nand03aa1n02x5               g016(.a(new_n111), .b(new_n107), .c(new_n108), .o1(new_n112));
  nor042aa1d18x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  inv040aa1n03x5               g018(.a(new_n113), .o1(new_n114));
  nand42aa1n16x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  oai112aa1n03x5               g020(.a(new_n114), .b(new_n115), .c(\b[5] ), .d(\a[6] ), .o1(new_n116));
  aoi022aa1d24x5               g021(.a(\b[7] ), .b(\a[8] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n117));
  tech160nm_fioai012aa1n04x5   g022(.a(new_n117), .b(\b[7] ), .c(\a[8] ), .o1(new_n118));
  nona32aa1n09x5               g023(.a(new_n106), .b(new_n118), .c(new_n116), .d(new_n112), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\b[5] ), .o1(new_n120));
  nanb02aa1d24x5               g025(.a(\a[6] ), .b(new_n120), .out0(new_n121));
  oai112aa1n06x5               g026(.a(new_n121), .b(new_n108), .c(\b[4] ), .d(\a[5] ), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .out0(new_n123));
  nano22aa1n03x7               g028(.a(new_n113), .b(new_n108), .c(new_n115), .out0(new_n124));
  oaoi03aa1n03x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n114), .o1(new_n125));
  aoi013aa1n09x5               g030(.a(new_n125), .b(new_n124), .c(new_n123), .d(new_n122), .o1(new_n126));
  aoi022aa1n09x5               g031(.a(new_n119), .b(new_n126), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  inv000aa1d42x5               g032(.a(\b[8] ), .o1(new_n128));
  nanb02aa1n03x5               g033(.a(\a[9] ), .b(new_n128), .out0(new_n129));
  norb02aa1n02x5               g034(.a(new_n129), .b(new_n127), .out0(new_n130));
  orn002aa1n24x5               g035(.a(\a[10] ), .b(\b[9] ), .o(new_n131));
  nand02aa1n06x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  oai112aa1n06x5               g037(.a(new_n131), .b(new_n132), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  oai022aa1n02x5               g038(.a(new_n130), .b(new_n97), .c(new_n127), .d(new_n133), .o1(\s[10] ));
  nand42aa1n03x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor002aa1d32x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n06x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  oai012aa1n02x5               g042(.a(new_n132), .b(new_n127), .c(new_n133), .o1(new_n138));
  aoi022aa1d24x5               g043(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n139));
  oai122aa1n02x7               g044(.a(new_n139), .b(new_n127), .c(new_n133), .d(\a[11] ), .e(\b[10] ), .o1(new_n140));
  aobi12aa1n02x7               g045(.a(new_n140), .b(new_n138), .c(new_n137), .out0(\s[11] ));
  oaoi13aa1n02x5               g046(.a(new_n136), .b(new_n139), .c(new_n127), .d(new_n133), .o1(new_n142));
  nor022aa1n16x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1d06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n06x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  norb03aa1n02x5               g050(.a(new_n144), .b(new_n136), .c(new_n143), .out0(new_n146));
  nand22aa1n03x5               g051(.a(new_n140), .b(new_n146), .o1(new_n147));
  oai012aa1n02x5               g052(.a(new_n147), .b(new_n142), .c(new_n145), .o1(\s[12] ));
  nona22aa1n02x4               g053(.a(new_n99), .b(new_n98), .c(new_n100), .out0(new_n149));
  nano22aa1n02x4               g054(.a(new_n103), .b(new_n99), .c(new_n102), .out0(new_n150));
  aoi012aa1n02x5               g055(.a(new_n105), .b(new_n150), .c(new_n149), .o1(new_n151));
  inv000aa1n02x5               g056(.a(new_n107), .o1(new_n152));
  oai012aa1n02x5               g057(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .o1(new_n153));
  nor042aa1n02x5               g058(.a(new_n153), .b(new_n152), .o1(new_n154));
  norp02aa1n02x5               g059(.a(\b[5] ), .b(\a[6] ), .o1(new_n155));
  norb03aa1n02x7               g060(.a(new_n115), .b(new_n155), .c(new_n113), .out0(new_n156));
  nanb03aa1n02x5               g061(.a(new_n118), .b(new_n154), .c(new_n156), .out0(new_n157));
  oai012aa1n06x5               g062(.a(new_n126), .b(new_n151), .c(new_n157), .o1(new_n158));
  nand42aa1n04x5               g063(.a(new_n131), .b(new_n132), .o1(new_n159));
  xnrc02aa1n03x5               g064(.a(\b[8] ), .b(\a[9] ), .out0(new_n160));
  inv030aa1n03x5               g065(.a(new_n160), .o1(new_n161));
  nona23aa1d18x5               g066(.a(new_n161), .b(new_n145), .c(new_n159), .d(new_n137), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(new_n158), .b(new_n163), .o1(new_n164));
  oai022aa1n02x5               g069(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n165));
  aoai13aa1n03x5               g070(.a(new_n144), .b(new_n165), .c(new_n133), .d(new_n139), .o1(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n162), .c(new_n119), .d(new_n126), .o1(new_n167));
  nor002aa1d32x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  nand42aa1n20x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  oai012aa1n02x5               g075(.a(new_n144), .b(new_n143), .c(new_n136), .o1(new_n171));
  oaib12aa1n02x5               g076(.a(new_n171), .b(new_n168), .c(new_n169), .out0(new_n172));
  aoi013aa1n02x4               g077(.a(new_n172), .b(new_n133), .c(new_n146), .d(new_n139), .o1(new_n173));
  aoi022aa1n02x5               g078(.a(new_n167), .b(new_n170), .c(new_n164), .d(new_n173), .o1(\s[13] ));
  inv000aa1d42x5               g079(.a(new_n168), .o1(new_n175));
  nona23aa1n09x5               g080(.a(new_n139), .b(new_n144), .c(new_n143), .d(new_n136), .out0(new_n176));
  aoai13aa1n06x5               g081(.a(new_n171), .b(new_n176), .c(new_n97), .d(new_n129), .o1(new_n177));
  aoai13aa1n02x7               g082(.a(new_n170), .b(new_n177), .c(new_n158), .d(new_n163), .o1(new_n178));
  nor002aa1d32x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nand42aa1d28x5               g084(.a(\b[13] ), .b(\a[14] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  norb03aa1d15x5               g086(.a(new_n180), .b(new_n168), .c(new_n179), .out0(new_n182));
  nanp02aa1n02x5               g087(.a(new_n178), .b(new_n182), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n183), .b(new_n181), .c(new_n175), .d(new_n178), .o1(\s[14] ));
  nano23aa1n03x7               g089(.a(new_n168), .b(new_n179), .c(new_n180), .d(new_n169), .out0(new_n185));
  oaoi03aa1n02x5               g090(.a(\a[14] ), .b(\b[13] ), .c(new_n175), .o1(new_n186));
  nor002aa1d32x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  nanp02aa1n24x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  norb02aa1n12x5               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n186), .c(new_n167), .d(new_n185), .o1(new_n190));
  aoi112aa1n02x5               g095(.a(new_n189), .b(new_n186), .c(new_n167), .d(new_n185), .o1(new_n191));
  norb02aa1n02x5               g096(.a(new_n190), .b(new_n191), .out0(\s[15] ));
  inv000aa1d42x5               g097(.a(new_n187), .o1(new_n193));
  nor042aa1n12x5               g098(.a(\b[15] ), .b(\a[16] ), .o1(new_n194));
  nand22aa1n12x5               g099(.a(\b[15] ), .b(\a[16] ), .o1(new_n195));
  norb02aa1n12x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  nona23aa1n03x5               g101(.a(new_n190), .b(new_n195), .c(new_n194), .d(new_n187), .out0(new_n197));
  aoai13aa1n02x5               g102(.a(new_n197), .b(new_n196), .c(new_n193), .d(new_n190), .o1(\s[16] ));
  nand23aa1n03x5               g103(.a(new_n185), .b(new_n189), .c(new_n196), .o1(new_n199));
  nor042aa1n03x5               g104(.a(new_n162), .b(new_n199), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(new_n158), .b(new_n200), .o1(new_n201));
  nona23aa1n02x4               g106(.a(new_n135), .b(new_n144), .c(new_n143), .d(new_n136), .out0(new_n202));
  nona23aa1n03x5               g107(.a(new_n180), .b(new_n169), .c(new_n168), .d(new_n179), .out0(new_n203));
  nano22aa1n03x7               g108(.a(new_n203), .b(new_n189), .c(new_n196), .out0(new_n204));
  nona32aa1n03x5               g109(.a(new_n204), .b(new_n202), .c(new_n160), .d(new_n159), .out0(new_n205));
  oai012aa1n02x5               g110(.a(new_n180), .b(\b[14] ), .c(\a[15] ), .o1(new_n206));
  nanb03aa1n02x5               g111(.a(new_n194), .b(new_n195), .c(new_n188), .out0(new_n207));
  tech160nm_fioai012aa1n03p5x5 g112(.a(new_n195), .b(new_n194), .c(new_n187), .o1(new_n208));
  oai013aa1n03x4               g113(.a(new_n208), .b(new_n182), .c(new_n207), .d(new_n206), .o1(new_n209));
  tech160nm_fiaoi012aa1n05x5   g114(.a(new_n209), .b(new_n177), .c(new_n204), .o1(new_n210));
  aoai13aa1n12x5               g115(.a(new_n210), .b(new_n205), .c(new_n119), .d(new_n126), .o1(new_n211));
  xorc02aa1n12x5               g116(.a(\a[17] ), .b(\b[16] ), .out0(new_n212));
  inv000aa1d42x5               g117(.a(new_n182), .o1(new_n213));
  nano23aa1n02x4               g118(.a(new_n206), .b(new_n194), .c(new_n188), .d(new_n195), .out0(new_n214));
  nanb02aa1n02x5               g119(.a(new_n212), .b(new_n208), .out0(new_n215));
  aoi122aa1n02x5               g120(.a(new_n215), .b(new_n213), .c(new_n214), .d(new_n177), .e(new_n204), .o1(new_n216));
  aoi022aa1n02x5               g121(.a(new_n211), .b(new_n212), .c(new_n201), .d(new_n216), .o1(\s[17] ));
  nor002aa1d32x5               g122(.a(\b[16] ), .b(\a[17] ), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aobi12aa1n02x5               g124(.a(new_n208), .b(new_n214), .c(new_n213), .out0(new_n220));
  oai012aa1n06x5               g125(.a(new_n220), .b(new_n166), .c(new_n199), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n212), .b(new_n221), .c(new_n158), .d(new_n200), .o1(new_n222));
  nor002aa1n08x5               g127(.a(\b[17] ), .b(\a[18] ), .o1(new_n223));
  nand02aa1n03x5               g128(.a(\b[17] ), .b(\a[18] ), .o1(new_n224));
  norb02aa1n03x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  norp02aa1n02x5               g130(.a(new_n223), .b(new_n218), .o1(new_n226));
  nand03aa1n02x5               g131(.a(new_n222), .b(new_n224), .c(new_n226), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n227), .b(new_n225), .c(new_n219), .d(new_n222), .o1(\s[18] ));
  and002aa1n02x5               g133(.a(new_n212), .b(new_n225), .o(new_n229));
  oaoi03aa1n02x5               g134(.a(\a[18] ), .b(\b[17] ), .c(new_n219), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[19] ), .b(\b[18] ), .out0(new_n231));
  aoai13aa1n04x5               g136(.a(new_n231), .b(new_n230), .c(new_n211), .d(new_n229), .o1(new_n232));
  aoi112aa1n02x7               g137(.a(new_n231), .b(new_n230), .c(new_n211), .d(new_n229), .o1(new_n233));
  norb02aa1n03x4               g138(.a(new_n232), .b(new_n233), .out0(\s[19] ));
  xnrc02aa1n02x5               g139(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g140(.a(\a[19] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(\b[18] ), .o1(new_n237));
  nanp02aa1n04x5               g142(.a(new_n237), .b(new_n236), .o1(new_n238));
  nor042aa1n06x5               g143(.a(\b[19] ), .b(\a[20] ), .o1(new_n239));
  nand42aa1n04x5               g144(.a(\b[19] ), .b(\a[20] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  nano22aa1n02x4               g146(.a(new_n239), .b(new_n238), .c(new_n240), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n232), .b(new_n242), .o1(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n241), .c(new_n238), .d(new_n232), .o1(\s[20] ));
  tech160nm_finand02aa1n03p5x5 g149(.a(\b[18] ), .b(\a[19] ), .o1(new_n245));
  nano32aa1n03x7               g150(.a(new_n239), .b(new_n238), .c(new_n240), .d(new_n245), .out0(new_n246));
  nand23aa1n09x5               g151(.a(new_n246), .b(new_n212), .c(new_n225), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  nanb03aa1n06x5               g153(.a(new_n239), .b(new_n240), .c(new_n245), .out0(new_n249));
  oai112aa1n03x5               g154(.a(new_n224), .b(new_n238), .c(new_n223), .d(new_n218), .o1(new_n250));
  aoai13aa1n04x5               g155(.a(new_n240), .b(new_n239), .c(new_n236), .d(new_n237), .o1(new_n251));
  oai012aa1n06x5               g156(.a(new_n251), .b(new_n250), .c(new_n249), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[21] ), .b(\b[20] ), .out0(new_n253));
  aoai13aa1n04x5               g158(.a(new_n253), .b(new_n252), .c(new_n211), .d(new_n248), .o1(new_n254));
  nano22aa1n02x4               g159(.a(new_n239), .b(new_n245), .c(new_n240), .out0(new_n255));
  oai012aa1n02x5               g160(.a(new_n224), .b(\b[18] ), .c(\a[19] ), .o1(new_n256));
  nona22aa1n03x5               g161(.a(new_n255), .b(new_n226), .c(new_n256), .out0(new_n257));
  nano22aa1n02x4               g162(.a(new_n253), .b(new_n257), .c(new_n251), .out0(new_n258));
  aobi12aa1n02x5               g163(.a(new_n258), .b(new_n211), .c(new_n248), .out0(new_n259));
  norb02aa1n03x4               g164(.a(new_n254), .b(new_n259), .out0(\s[21] ));
  nor042aa1n09x5               g165(.a(\b[20] ), .b(\a[21] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  nor042aa1n03x5               g167(.a(\b[21] ), .b(\a[22] ), .o1(new_n263));
  and002aa1n12x5               g168(.a(\b[21] ), .b(\a[22] ), .o(new_n264));
  nor042aa1n04x5               g169(.a(new_n264), .b(new_n263), .o1(new_n265));
  norp03aa1n02x5               g170(.a(new_n264), .b(new_n263), .c(new_n261), .o1(new_n266));
  nanp02aa1n03x5               g171(.a(new_n254), .b(new_n266), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n265), .c(new_n262), .d(new_n254), .o1(\s[22] ));
  nanp02aa1n06x5               g173(.a(new_n253), .b(new_n265), .o1(new_n269));
  nano32aa1n02x4               g174(.a(new_n269), .b(new_n246), .c(new_n225), .d(new_n212), .out0(new_n270));
  oab012aa1n02x4               g175(.a(new_n264), .b(new_n261), .c(new_n263), .out0(new_n271));
  inv000aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  aoai13aa1n04x5               g177(.a(new_n272), .b(new_n269), .c(new_n257), .d(new_n251), .o1(new_n273));
  nor022aa1n08x5               g178(.a(\b[22] ), .b(\a[23] ), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(\b[22] ), .b(\a[23] ), .o1(new_n275));
  norb02aa1n02x5               g180(.a(new_n275), .b(new_n274), .out0(new_n276));
  aoai13aa1n04x5               g181(.a(new_n276), .b(new_n273), .c(new_n211), .d(new_n270), .o1(new_n277));
  inv030aa1n04x5               g182(.a(new_n269), .o1(new_n278));
  aoi112aa1n02x5               g183(.a(new_n276), .b(new_n271), .c(new_n252), .d(new_n278), .o1(new_n279));
  aobi12aa1n02x5               g184(.a(new_n279), .b(new_n211), .c(new_n270), .out0(new_n280));
  norb02aa1n03x4               g185(.a(new_n277), .b(new_n280), .out0(\s[23] ));
  inv000aa1n02x5               g186(.a(new_n274), .o1(new_n282));
  nor042aa1n02x5               g187(.a(\b[23] ), .b(\a[24] ), .o1(new_n283));
  and002aa1n02x5               g188(.a(\b[23] ), .b(\a[24] ), .o(new_n284));
  norp02aa1n02x5               g189(.a(new_n284), .b(new_n283), .o1(new_n285));
  norp03aa1n02x5               g190(.a(new_n284), .b(new_n283), .c(new_n274), .o1(new_n286));
  nanp02aa1n03x5               g191(.a(new_n277), .b(new_n286), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n285), .c(new_n282), .d(new_n277), .o1(\s[24] ));
  nano23aa1n03x7               g193(.a(new_n284), .b(new_n283), .c(new_n282), .d(new_n275), .out0(new_n289));
  nano32aa1n02x5               g194(.a(new_n247), .b(new_n289), .c(new_n253), .d(new_n265), .out0(new_n290));
  aobi12aa1n02x5               g195(.a(new_n290), .b(new_n201), .c(new_n210), .out0(new_n291));
  aoai13aa1n02x5               g196(.a(new_n289), .b(new_n271), .c(new_n252), .d(new_n278), .o1(new_n292));
  oab012aa1n04x5               g197(.a(new_n284), .b(new_n274), .c(new_n283), .out0(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  nanp02aa1n02x5               g199(.a(new_n292), .b(new_n294), .o1(new_n295));
  tech160nm_fixorc02aa1n03p5x5 g200(.a(\a[25] ), .b(\b[24] ), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n296), .b(new_n295), .c(new_n211), .d(new_n290), .o1(new_n297));
  nona22aa1n02x4               g202(.a(new_n292), .b(new_n293), .c(new_n296), .out0(new_n298));
  oa0012aa1n03x5               g203(.a(new_n297), .b(new_n298), .c(new_n291), .o(\s[25] ));
  nor042aa1n03x5               g204(.a(\b[24] ), .b(\a[25] ), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  nor002aa1n02x5               g206(.a(\b[25] ), .b(\a[26] ), .o1(new_n302));
  and002aa1n12x5               g207(.a(\b[25] ), .b(\a[26] ), .o(new_n303));
  nor022aa1n04x5               g208(.a(new_n303), .b(new_n302), .o1(new_n304));
  norp03aa1n02x5               g209(.a(new_n303), .b(new_n302), .c(new_n300), .o1(new_n305));
  nand02aa1n02x5               g210(.a(new_n297), .b(new_n305), .o1(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n304), .c(new_n301), .d(new_n297), .o1(\s[26] ));
  and002aa1n02x5               g212(.a(new_n296), .b(new_n304), .o(new_n308));
  aoai13aa1n06x5               g213(.a(new_n308), .b(new_n293), .c(new_n273), .d(new_n289), .o1(new_n309));
  nano32aa1n03x7               g214(.a(new_n247), .b(new_n308), .c(new_n278), .d(new_n289), .out0(new_n310));
  aoai13aa1n06x5               g215(.a(new_n310), .b(new_n221), .c(new_n158), .d(new_n200), .o1(new_n311));
  oab012aa1n09x5               g216(.a(new_n303), .b(new_n300), .c(new_n302), .out0(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  nand23aa1n06x5               g218(.a(new_n311), .b(new_n309), .c(new_n313), .o1(new_n314));
  xorc02aa1n12x5               g219(.a(\a[27] ), .b(\b[26] ), .out0(new_n315));
  aoi112aa1n02x7               g220(.a(new_n315), .b(new_n312), .c(new_n211), .d(new_n310), .o1(new_n316));
  aoi022aa1n03x5               g221(.a(new_n316), .b(new_n309), .c(new_n314), .d(new_n315), .o1(\s[27] ));
  norp02aa1n02x5               g222(.a(\b[26] ), .b(\a[27] ), .o1(new_n318));
  xnrc02aa1n12x5               g223(.a(\b[27] ), .b(\a[28] ), .out0(new_n319));
  aoai13aa1n02x7               g224(.a(new_n319), .b(new_n318), .c(new_n314), .d(new_n315), .o1(new_n320));
  aobi12aa1n06x5               g225(.a(new_n308), .b(new_n292), .c(new_n294), .out0(new_n321));
  aoi112aa1n06x5               g226(.a(new_n321), .b(new_n312), .c(new_n211), .d(new_n310), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n315), .o1(new_n323));
  oai022aa1d18x5               g228(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n324));
  aoi012aa1n02x5               g229(.a(new_n324), .b(\a[28] ), .c(\b[27] ), .o1(new_n325));
  oai012aa1n03x5               g230(.a(new_n325), .b(new_n322), .c(new_n323), .o1(new_n326));
  nanp02aa1n03x5               g231(.a(new_n320), .b(new_n326), .o1(\s[28] ));
  xnrc02aa1n12x5               g232(.a(\b[28] ), .b(\a[29] ), .out0(new_n328));
  norb02aa1d21x5               g233(.a(new_n315), .b(new_n319), .out0(new_n329));
  inv000aa1d42x5               g234(.a(\a[28] ), .o1(new_n330));
  inv000aa1d42x5               g235(.a(\b[27] ), .o1(new_n331));
  oao003aa1n02x5               g236(.a(new_n330), .b(new_n331), .c(new_n318), .carry(new_n332));
  aoai13aa1n02x7               g237(.a(new_n328), .b(new_n332), .c(new_n314), .d(new_n329), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n329), .o1(new_n334));
  norp02aa1n02x5               g239(.a(new_n332), .b(new_n328), .o1(new_n335));
  oai012aa1n03x5               g240(.a(new_n335), .b(new_n322), .c(new_n334), .o1(new_n336));
  nanp02aa1n03x5               g241(.a(new_n333), .b(new_n336), .o1(\s[29] ));
  xorb03aa1n02x5               g242(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1d15x5               g243(.a(new_n315), .b(new_n328), .c(new_n319), .out0(new_n339));
  nanp02aa1n02x5               g244(.a(\b[28] ), .b(\a[29] ), .o1(new_n340));
  oai112aa1n06x5               g245(.a(new_n324), .b(new_n340), .c(new_n331), .d(new_n330), .o1(new_n341));
  oai012aa1n02x5               g246(.a(new_n341), .b(\b[28] ), .c(\a[29] ), .o1(new_n342));
  norp02aa1n02x5               g247(.a(\b[29] ), .b(\a[30] ), .o1(new_n343));
  nanp02aa1n02x5               g248(.a(\b[29] ), .b(\a[30] ), .o1(new_n344));
  nanb02aa1n02x5               g249(.a(new_n343), .b(new_n344), .out0(new_n345));
  aoai13aa1n02x7               g250(.a(new_n345), .b(new_n342), .c(new_n314), .d(new_n339), .o1(new_n346));
  inv000aa1d42x5               g251(.a(new_n339), .o1(new_n347));
  norp02aa1n02x5               g252(.a(\b[28] ), .b(\a[29] ), .o1(new_n348));
  nona23aa1n06x5               g253(.a(new_n341), .b(new_n344), .c(new_n343), .d(new_n348), .out0(new_n349));
  inv000aa1d42x5               g254(.a(new_n349), .o1(new_n350));
  oai012aa1n03x5               g255(.a(new_n350), .b(new_n322), .c(new_n347), .o1(new_n351));
  nanp02aa1n03x5               g256(.a(new_n346), .b(new_n351), .o1(\s[30] ));
  norb03aa1n06x5               g257(.a(new_n329), .b(new_n328), .c(new_n345), .out0(new_n353));
  and002aa1n02x5               g258(.a(new_n349), .b(new_n344), .o(new_n354));
  xnrc02aa1n02x5               g259(.a(\b[30] ), .b(\a[31] ), .out0(new_n355));
  aoai13aa1n02x7               g260(.a(new_n355), .b(new_n354), .c(new_n314), .d(new_n353), .o1(new_n356));
  inv000aa1n02x5               g261(.a(new_n353), .o1(new_n357));
  tech160nm_fiaoi012aa1n05x5   g262(.a(new_n355), .b(new_n349), .c(new_n344), .o1(new_n358));
  oai012aa1n03x5               g263(.a(new_n358), .b(new_n322), .c(new_n357), .o1(new_n359));
  nanp02aa1n03x5               g264(.a(new_n356), .b(new_n359), .o1(\s[31] ));
  norp02aa1n02x5               g265(.a(new_n101), .b(new_n104), .o1(new_n361));
  inv000aa1d42x5               g266(.a(new_n103), .o1(new_n362));
  aoi022aa1n02x5               g267(.a(new_n149), .b(new_n99), .c(new_n362), .d(new_n102), .o1(new_n363));
  norp02aa1n02x5               g268(.a(new_n363), .b(new_n361), .o1(\s[3] ));
  inv000aa1n03x5               g269(.a(new_n361), .o1(new_n365));
  xorc02aa1n02x5               g270(.a(\a[4] ), .b(\b[3] ), .out0(new_n366));
  xnbna2aa1n03x5               g271(.a(new_n366), .b(new_n365), .c(new_n362), .out0(\s[4] ));
  inv000aa1d42x5               g272(.a(new_n111), .o1(new_n368));
  nanp02aa1n02x5               g273(.a(\b[3] ), .b(\a[4] ), .o1(new_n369));
  nona23aa1n02x4               g274(.a(new_n106), .b(new_n369), .c(new_n368), .d(new_n152), .out0(new_n370));
  aoi022aa1n02x5               g275(.a(new_n106), .b(new_n369), .c(new_n107), .d(new_n111), .o1(new_n371));
  norb02aa1n02x5               g276(.a(new_n370), .b(new_n371), .out0(\s[5] ));
  aoi013aa1n02x4               g277(.a(new_n368), .b(new_n106), .c(new_n107), .d(new_n369), .o1(new_n373));
  nanb02aa1n02x5               g278(.a(new_n122), .b(new_n370), .out0(new_n374));
  aoai13aa1n02x5               g279(.a(new_n374), .b(new_n373), .c(new_n108), .d(new_n121), .o1(\s[6] ));
  aoi022aa1n02x5               g280(.a(new_n374), .b(new_n108), .c(new_n114), .d(new_n115), .o1(new_n376));
  nanp02aa1n02x5               g281(.a(new_n374), .b(new_n124), .o1(new_n377));
  norb02aa1n02x5               g282(.a(new_n377), .b(new_n376), .out0(\s[7] ));
  xnbna2aa1n03x5               g283(.a(new_n123), .b(new_n377), .c(new_n114), .out0(\s[8] ));
  aoi113aa1n02x5               g284(.a(new_n161), .b(new_n125), .c(new_n124), .d(new_n123), .e(new_n122), .o1(new_n380));
  aoi022aa1n02x5               g285(.a(new_n158), .b(new_n161), .c(new_n119), .d(new_n380), .o1(\s[9] ));
endmodule


