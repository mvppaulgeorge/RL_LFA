// Benchmark "adder" written by ABC on Wed Jul 17 17:53:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n309, new_n310,
    new_n311, new_n313, new_n315, new_n317, new_n319, new_n320, new_n321,
    new_n322, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  oa0022aa1n06x5               g003(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n99));
  inv040aa1d24x5               g004(.a(\a[3] ), .o1(new_n100));
  inv040aa1d30x5               g005(.a(\b[2] ), .o1(new_n101));
  nand22aa1n06x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nand22aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand02aa1d04x5               g008(.a(new_n102), .b(new_n103), .o1(new_n104));
  nanp02aa1n09x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nor042aa1n06x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nand02aa1d28x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  oai012aa1d24x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .o1(new_n108));
  oai012aa1n12x5               g013(.a(new_n99), .b(new_n108), .c(new_n104), .o1(new_n109));
  nand02aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1n06x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  norp02aa1n12x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanb03aa1n06x5               g017(.a(new_n112), .b(new_n110), .c(new_n111), .out0(new_n113));
  oai022aa1n02x5               g018(.a(\a[6] ), .b(\b[5] ), .c(\b[6] ), .d(\a[7] ), .o1(new_n114));
  aoi022aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n115));
  inv040aa1d32x5               g020(.a(\a[5] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[4] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(new_n117), .b(new_n116), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[3] ), .b(\a[4] ), .o1(new_n119));
  nand03aa1n02x5               g024(.a(new_n115), .b(new_n118), .c(new_n119), .o1(new_n120));
  nor043aa1n03x5               g025(.a(new_n120), .b(new_n113), .c(new_n114), .o1(new_n121));
  inv000aa1n02x5               g026(.a(new_n112), .o1(new_n122));
  inv040aa1d32x5               g027(.a(\a[7] ), .o1(new_n123));
  inv030aa1d32x5               g028(.a(\b[6] ), .o1(new_n124));
  nanp02aa1n09x5               g029(.a(new_n124), .b(new_n123), .o1(new_n125));
  nor022aa1n04x5               g030(.a(\b[5] ), .b(\a[6] ), .o1(new_n126));
  aoai13aa1n04x5               g031(.a(new_n111), .b(new_n126), .c(new_n117), .d(new_n116), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(\b[6] ), .b(\a[7] ), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(new_n128), .b(new_n110), .o1(new_n129));
  aoai13aa1n06x5               g034(.a(new_n122), .b(new_n129), .c(new_n127), .d(new_n125), .o1(new_n130));
  aoi012aa1n12x5               g035(.a(new_n130), .b(new_n121), .c(new_n109), .o1(new_n131));
  tech160nm_fixnrc02aa1n04x5   g036(.a(\b[8] ), .b(\a[9] ), .out0(new_n132));
  orn002aa1n02x5               g037(.a(new_n131), .b(new_n132), .o(new_n133));
  xnrc02aa1n06x5               g038(.a(\b[9] ), .b(\a[10] ), .out0(new_n134));
  xobna2aa1n03x5               g039(.a(new_n134), .b(new_n133), .c(new_n98), .out0(\s[10] ));
  orn002aa1n02x5               g040(.a(new_n132), .b(new_n134), .o(new_n136));
  nor042aa1n06x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nand02aa1n04x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  oai012aa1d24x5               g043(.a(new_n138), .b(new_n137), .c(new_n97), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  oab012aa1n02x4               g045(.a(new_n140), .b(new_n131), .c(new_n136), .out0(new_n141));
  xnrb03aa1n02x5               g046(.a(new_n141), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1n08x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  oaoi03aa1n02x5               g050(.a(\a[11] ), .b(\b[10] ), .c(new_n141), .o1(new_n146));
  nor002aa1d24x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  nanp02aa1n04x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nanb02aa1n02x5               g053(.a(new_n147), .b(new_n148), .out0(new_n149));
  norb03aa1n02x5               g054(.a(new_n144), .b(new_n147), .c(new_n143), .out0(new_n150));
  oai012aa1n02x5               g055(.a(new_n150), .b(new_n141), .c(new_n149), .o1(new_n151));
  aob012aa1n02x5               g056(.a(new_n151), .b(new_n146), .c(new_n145), .out0(\s[12] ));
  nona23aa1d18x5               g057(.a(new_n144), .b(new_n148), .c(new_n147), .d(new_n143), .out0(new_n153));
  nor043aa1n03x5               g058(.a(new_n153), .b(new_n134), .c(new_n132), .o1(new_n154));
  aoai13aa1n03x5               g059(.a(new_n154), .b(new_n130), .c(new_n121), .d(new_n109), .o1(new_n155));
  oaih12aa1n12x5               g060(.a(new_n144), .b(new_n143), .c(new_n147), .o1(new_n156));
  oai012aa1d24x5               g061(.a(new_n156), .b(new_n153), .c(new_n139), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nor002aa1d32x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanp02aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n155), .c(new_n158), .out0(\s[13] ));
  nanp02aa1n02x5               g067(.a(new_n155), .b(new_n158), .o1(new_n163));
  nor002aa1d32x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nand42aa1n08x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nanb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n159), .c(new_n163), .d(new_n160), .o1(new_n167));
  nona22aa1n02x4               g072(.a(new_n165), .b(new_n164), .c(new_n159), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n167), .b(new_n168), .c(new_n161), .d(new_n163), .o1(\s[14] ));
  nona23aa1n09x5               g074(.a(new_n165), .b(new_n160), .c(new_n159), .d(new_n164), .out0(new_n170));
  tech160nm_fioai012aa1n03p5x5 g075(.a(new_n165), .b(new_n164), .c(new_n159), .o1(new_n171));
  aoai13aa1n02x7               g076(.a(new_n171), .b(new_n170), .c(new_n155), .d(new_n158), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv040aa1d32x5               g078(.a(\a[15] ), .o1(new_n174));
  inv000aa1d42x5               g079(.a(\b[14] ), .o1(new_n175));
  nand02aa1d04x5               g080(.a(new_n175), .b(new_n174), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand22aa1n04x5               g082(.a(new_n176), .b(new_n177), .o1(new_n178));
  norb02aa1n06x5               g083(.a(new_n172), .b(new_n178), .out0(new_n179));
  xnrc02aa1n12x5               g084(.a(\b[15] ), .b(\a[16] ), .out0(new_n180));
  oaoi03aa1n02x5               g085(.a(new_n174), .b(new_n175), .c(new_n172), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n180), .b(new_n176), .out0(new_n182));
  obai22aa1n02x7               g087(.a(new_n180), .b(new_n181), .c(new_n179), .d(new_n182), .out0(\s[16] ));
  nor043aa1d12x5               g088(.a(new_n170), .b(new_n178), .c(new_n180), .o1(new_n184));
  nand02aa1d04x5               g089(.a(new_n184), .b(new_n154), .o1(new_n185));
  orn002aa1n02x5               g090(.a(\a[16] ), .b(\b[15] ), .o(new_n186));
  aob012aa1n02x5               g091(.a(new_n177), .b(\b[15] ), .c(\a[16] ), .out0(new_n187));
  aoai13aa1n06x5               g092(.a(new_n186), .b(new_n187), .c(new_n171), .d(new_n176), .o1(new_n188));
  aoi012aa1d18x5               g093(.a(new_n188), .b(new_n157), .c(new_n184), .o1(new_n189));
  oai012aa1d24x5               g094(.a(new_n189), .b(new_n131), .c(new_n185), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g096(.a(\b[16] ), .b(\a[17] ), .o1(new_n192));
  inv000aa1n06x5               g097(.a(new_n192), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  oaib12aa1n02x5               g099(.a(new_n190), .b(new_n194), .c(\b[16] ), .out0(new_n195));
  xorc02aa1n02x5               g100(.a(\a[18] ), .b(\b[17] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n195), .c(new_n193), .out0(\s[18] ));
  inv040aa1d32x5               g102(.a(\a[18] ), .o1(new_n198));
  xroi22aa1d06x4               g103(.a(new_n194), .b(\b[16] ), .c(new_n198), .d(\b[17] ), .out0(new_n199));
  oaoi03aa1n09x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n200));
  xorc02aa1n12x5               g105(.a(\a[19] ), .b(\b[18] ), .out0(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n202));
  aoi112aa1n02x5               g107(.a(new_n201), .b(new_n200), .c(new_n190), .d(new_n199), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n202), .b(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(\b[18] ), .b(new_n206), .out0(new_n207));
  xorc02aa1n12x5               g112(.a(\a[20] ), .b(\b[19] ), .out0(new_n208));
  nanp02aa1n02x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  oai022aa1n02x5               g114(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n210));
  nanb03aa1n03x5               g115(.a(new_n210), .b(new_n202), .c(new_n209), .out0(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n208), .c(new_n202), .d(new_n207), .o1(\s[20] ));
  nand03aa1n02x5               g117(.a(new_n199), .b(new_n201), .c(new_n208), .o1(new_n213));
  nanb02aa1n06x5               g118(.a(new_n213), .b(new_n190), .out0(new_n214));
  nanp03aa1d12x5               g119(.a(new_n200), .b(new_n201), .c(new_n208), .o1(new_n215));
  nand42aa1n02x5               g120(.a(new_n210), .b(new_n209), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  xorc02aa1n12x5               g123(.a(\a[21] ), .b(\b[20] ), .out0(new_n219));
  xnbna2aa1n06x5               g124(.a(new_n219), .b(new_n214), .c(new_n218), .out0(\s[21] ));
  aobi12aa1n02x7               g125(.a(new_n219), .b(new_n214), .c(new_n218), .out0(new_n221));
  nand42aa1n03x5               g126(.a(new_n214), .b(new_n218), .o1(new_n222));
  norp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  tech160nm_fixnrc02aa1n05x5   g128(.a(\b[21] ), .b(\a[22] ), .out0(new_n224));
  aoai13aa1n03x5               g129(.a(new_n224), .b(new_n223), .c(new_n222), .d(new_n219), .o1(new_n225));
  norp02aa1n02x5               g130(.a(new_n224), .b(new_n223), .o1(new_n226));
  oaib12aa1n03x5               g131(.a(new_n225), .b(new_n221), .c(new_n226), .out0(\s[22] ));
  nanb02aa1n06x5               g132(.a(new_n224), .b(new_n219), .out0(new_n228));
  nano32aa1n02x4               g133(.a(new_n228), .b(new_n199), .c(new_n201), .d(new_n208), .out0(new_n229));
  orn002aa1n02x5               g134(.a(\a[21] ), .b(\b[20] ), .o(new_n230));
  oao003aa1n02x5               g135(.a(\a[22] ), .b(\b[21] ), .c(new_n230), .carry(new_n231));
  aoai13aa1n12x5               g136(.a(new_n231), .b(new_n228), .c(new_n215), .d(new_n216), .o1(new_n232));
  xorc02aa1n12x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n232), .c(new_n190), .d(new_n229), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n233), .b(new_n232), .c(new_n190), .d(new_n229), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n234), .b(new_n235), .out0(\s[23] ));
  orn002aa1n02x5               g141(.a(\a[23] ), .b(\b[22] ), .o(new_n237));
  tech160nm_fixorc02aa1n05x5   g142(.a(\a[24] ), .b(\b[23] ), .out0(new_n238));
  nanp02aa1n02x5               g143(.a(\b[23] ), .b(\a[24] ), .o1(new_n239));
  oai022aa1n02x5               g144(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n240));
  nanb03aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n239), .out0(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n238), .c(new_n234), .d(new_n237), .o1(\s[24] ));
  norb02aa1n02x5               g147(.a(new_n219), .b(new_n224), .out0(new_n243));
  and002aa1n06x5               g148(.a(new_n238), .b(new_n233), .o(new_n244));
  nano22aa1n02x4               g149(.a(new_n213), .b(new_n244), .c(new_n243), .out0(new_n245));
  nanp02aa1n03x5               g150(.a(new_n190), .b(new_n245), .o1(new_n246));
  aoi022aa1n02x5               g151(.a(new_n232), .b(new_n244), .c(new_n239), .d(new_n240), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[25] ), .b(\b[24] ), .out0(new_n248));
  xnbna2aa1n03x5               g153(.a(new_n248), .b(new_n246), .c(new_n247), .out0(\s[25] ));
  aobi12aa1n02x5               g154(.a(new_n248), .b(new_n246), .c(new_n247), .out0(new_n250));
  xorc02aa1n02x5               g155(.a(\a[26] ), .b(\b[25] ), .out0(new_n251));
  nanp02aa1n03x5               g156(.a(new_n246), .b(new_n247), .o1(new_n252));
  norp02aa1n02x5               g157(.a(\b[24] ), .b(\a[25] ), .o1(new_n253));
  aoi012aa1n03x5               g158(.a(new_n253), .b(new_n252), .c(new_n248), .o1(new_n254));
  nanp02aa1n02x5               g159(.a(\b[25] ), .b(\a[26] ), .o1(new_n255));
  oai022aa1n02x5               g160(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n256));
  nanb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  oai022aa1n03x5               g162(.a(new_n254), .b(new_n251), .c(new_n257), .d(new_n250), .o1(\s[26] ));
  oaoi03aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .o1(new_n259));
  and002aa1n02x5               g164(.a(new_n251), .b(new_n248), .o(new_n260));
  aoai13aa1n12x5               g165(.a(new_n260), .b(new_n259), .c(new_n232), .d(new_n244), .o1(new_n261));
  nor042aa1n03x5               g166(.a(\b[26] ), .b(\a[27] ), .o1(new_n262));
  and002aa1n02x5               g167(.a(\b[26] ), .b(\a[27] ), .o(new_n263));
  norp02aa1n02x5               g168(.a(new_n263), .b(new_n262), .o1(new_n264));
  nano32aa1n03x7               g169(.a(new_n213), .b(new_n260), .c(new_n243), .d(new_n244), .out0(new_n265));
  aoi122aa1n02x5               g170(.a(new_n264), .b(new_n255), .c(new_n256), .d(new_n190), .e(new_n265), .o1(new_n266));
  nand02aa1d06x5               g171(.a(new_n190), .b(new_n265), .o1(new_n267));
  nanp02aa1n02x5               g172(.a(new_n256), .b(new_n255), .o1(new_n268));
  nand03aa1n06x5               g173(.a(new_n261), .b(new_n267), .c(new_n268), .o1(new_n269));
  aoi022aa1n02x5               g174(.a(new_n261), .b(new_n266), .c(new_n269), .d(new_n264), .o1(\s[27] ));
  inv000aa1d42x5               g175(.a(\b[26] ), .o1(new_n271));
  oaib12aa1n03x5               g176(.a(new_n269), .b(new_n271), .c(\a[27] ), .out0(new_n272));
  inv000aa1n03x5               g177(.a(new_n262), .o1(new_n273));
  aoi022aa1n09x5               g178(.a(new_n190), .b(new_n265), .c(new_n255), .d(new_n256), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n273), .b(new_n263), .c(new_n274), .d(new_n261), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[28] ), .b(\b[27] ), .out0(new_n276));
  norp02aa1n02x5               g181(.a(new_n276), .b(new_n262), .o1(new_n277));
  aoi022aa1n03x5               g182(.a(new_n275), .b(new_n276), .c(new_n272), .d(new_n277), .o1(\s[28] ));
  inv000aa1d42x5               g183(.a(\a[28] ), .o1(new_n279));
  xroi22aa1d04x5               g184(.a(\a[27] ), .b(new_n271), .c(new_n279), .d(\b[27] ), .out0(new_n280));
  nanp02aa1n02x5               g185(.a(new_n269), .b(new_n280), .o1(new_n281));
  inv000aa1n06x5               g186(.a(new_n280), .o1(new_n282));
  oao003aa1n03x5               g187(.a(\a[28] ), .b(\b[27] ), .c(new_n273), .carry(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n282), .c(new_n274), .d(new_n261), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[29] ), .b(\b[28] ), .out0(new_n285));
  norb02aa1n02x5               g190(.a(new_n283), .b(new_n285), .out0(new_n286));
  aoi022aa1n03x5               g191(.a(new_n284), .b(new_n285), .c(new_n281), .d(new_n286), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g193(.a(new_n276), .b(new_n285), .c(new_n264), .o(new_n289));
  nanp02aa1n03x5               g194(.a(new_n269), .b(new_n289), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n289), .o1(new_n291));
  oaoi03aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .c(new_n283), .o1(new_n292));
  inv000aa1n03x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n291), .c(new_n274), .d(new_n261), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[30] ), .b(\b[29] ), .out0(new_n295));
  and002aa1n02x5               g200(.a(\b[28] ), .b(\a[29] ), .o(new_n296));
  oabi12aa1n02x5               g201(.a(new_n295), .b(\a[29] ), .c(\b[28] ), .out0(new_n297));
  oab012aa1n02x4               g202(.a(new_n297), .b(new_n283), .c(new_n296), .out0(new_n298));
  aoi022aa1n03x5               g203(.a(new_n294), .b(new_n295), .c(new_n290), .d(new_n298), .o1(\s[30] ));
  nano22aa1n02x4               g204(.a(new_n282), .b(new_n285), .c(new_n295), .out0(new_n300));
  nanp02aa1n02x5               g205(.a(new_n269), .b(new_n300), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[31] ), .b(\b[30] ), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n303));
  norb02aa1n02x5               g208(.a(new_n303), .b(new_n302), .out0(new_n304));
  inv000aa1n02x5               g209(.a(new_n300), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n303), .b(new_n305), .c(new_n274), .d(new_n261), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[31] ));
  xnbna2aa1n03x5               g212(.a(new_n108), .b(new_n102), .c(new_n103), .out0(\s[3] ));
  orn002aa1n02x5               g213(.a(new_n108), .b(new_n104), .o(new_n309));
  xorc02aa1n02x5               g214(.a(\a[4] ), .b(\b[3] ), .out0(new_n310));
  norb02aa1n02x5               g215(.a(new_n102), .b(new_n310), .out0(new_n311));
  aoi022aa1n02x5               g216(.a(new_n309), .b(new_n311), .c(new_n109), .d(new_n310), .o1(\s[4] ));
  and002aa1n03x5               g217(.a(new_n109), .b(new_n119), .o(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g219(.a(new_n116), .b(new_n117), .c(new_n313), .o1(new_n315));
  xnrb03aa1n02x5               g220(.a(new_n315), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fioaoi03aa1n03p5x5 g221(.a(\a[6] ), .b(\b[5] ), .c(new_n315), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  inv000aa1d42x5               g223(.a(new_n125), .o1(new_n319));
  norb02aa1n02x5               g224(.a(new_n110), .b(new_n112), .out0(new_n320));
  inv000aa1d42x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n02x5               g226(.a(new_n321), .b(new_n319), .c(new_n317), .d(new_n128), .o1(new_n322));
  aoi112aa1n03x5               g227(.a(new_n321), .b(new_n319), .c(new_n317), .d(new_n128), .o1(new_n323));
  nanb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(\s[8] ));
  xnrb03aa1n02x5               g229(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


