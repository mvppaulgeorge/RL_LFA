// Benchmark "adder" written by ABC on Wed Jul 17 21:27:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n324,
    new_n327, new_n329, new_n330, new_n332, new_n333;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n09x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n12x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\a[9] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[8] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  nor042aa1n02x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand42aa1n16x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  tech160nm_finor002aa1n05x5   g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n02x4               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  inv000aa1d42x5               g013(.a(\a[2] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[1] ), .o1(new_n110));
  nand22aa1n03x5               g015(.a(\b[0] ), .b(\a[1] ), .o1(new_n111));
  tech160nm_fioaoi03aa1n02p5x5 g016(.a(new_n109), .b(new_n110), .c(new_n111), .o1(new_n112));
  aoi012aa1n03x5               g017(.a(new_n104), .b(new_n106), .c(new_n105), .o1(new_n113));
  oai012aa1n02x7               g018(.a(new_n113), .b(new_n108), .c(new_n112), .o1(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  norp02aa1n04x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand22aa1n06x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor022aa1n06x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand42aa1n04x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nona23aa1n09x5               g024(.a(new_n119), .b(new_n117), .c(new_n116), .d(new_n118), .out0(new_n120));
  xnrc02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .out0(new_n121));
  nor003aa1n02x5               g026(.a(new_n120), .b(new_n121), .c(new_n115), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[5] ), .o1(new_n123));
  oai022aa1n02x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  oaib12aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(\a[6] ), .out0(new_n125));
  tech160nm_fiao0012aa1n02p5x5 g030(.a(new_n116), .b(new_n118), .c(new_n117), .o(new_n126));
  oabi12aa1n06x5               g031(.a(new_n126), .b(new_n120), .c(new_n125), .out0(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n114), .d(new_n122), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n100), .b(new_n129), .c(new_n103), .out0(\s[10] ));
  nano23aa1n03x5               g035(.a(new_n104), .b(new_n106), .c(new_n107), .d(new_n105), .out0(new_n131));
  oao003aa1n02x5               g036(.a(new_n109), .b(new_n110), .c(new_n111), .carry(new_n132));
  aobi12aa1n06x5               g037(.a(new_n113), .b(new_n131), .c(new_n132), .out0(new_n133));
  nano23aa1n03x7               g038(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n134));
  nona22aa1n03x5               g039(.a(new_n134), .b(new_n121), .c(new_n115), .out0(new_n135));
  inv040aa1n04x5               g040(.a(new_n127), .o1(new_n136));
  oai012aa1n12x5               g041(.a(new_n136), .b(new_n133), .c(new_n135), .o1(new_n137));
  aoai13aa1n12x5               g042(.a(new_n98), .b(new_n97), .c(new_n101), .d(new_n102), .o1(new_n138));
  inv040aa1n03x5               g043(.a(new_n138), .o1(new_n139));
  aoi013aa1n06x4               g044(.a(new_n139), .b(new_n137), .c(new_n128), .d(new_n100), .o1(new_n140));
  nor002aa1d32x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  nand22aa1n04x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  xnbna2aa1n03x5               g048(.a(new_n140), .b(new_n143), .c(new_n142), .out0(\s[11] ));
  oaoi03aa1n02x5               g049(.a(\a[11] ), .b(\b[10] ), .c(new_n140), .o1(new_n145));
  xorb03aa1n02x5               g050(.a(new_n145), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  xnrc02aa1n02x5               g051(.a(\b[8] ), .b(\a[9] ), .out0(new_n147));
  nor022aa1n16x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  nand22aa1n09x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nano23aa1n06x5               g054(.a(new_n141), .b(new_n148), .c(new_n149), .d(new_n143), .out0(new_n150));
  nona23aa1n03x5               g055(.a(new_n137), .b(new_n150), .c(new_n147), .d(new_n99), .out0(new_n151));
  nona23aa1d18x5               g056(.a(new_n149), .b(new_n143), .c(new_n141), .d(new_n148), .out0(new_n152));
  aoi012aa1n09x5               g057(.a(new_n148), .b(new_n141), .c(new_n149), .o1(new_n153));
  oai012aa1n18x5               g058(.a(new_n153), .b(new_n152), .c(new_n138), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  nor042aa1n06x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1n02x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n157), .b(new_n156), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n151), .c(new_n155), .out0(\s[13] ));
  inv000aa1n06x5               g064(.a(new_n156), .o1(new_n160));
  inv020aa1n02x5               g065(.a(new_n158), .o1(new_n161));
  aoai13aa1n03x5               g066(.a(new_n160), .b(new_n161), .c(new_n151), .d(new_n155), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n156), .b(new_n164), .c(new_n165), .d(new_n157), .out0(new_n166));
  oaoi03aa1n12x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n154), .c(new_n166), .o1(new_n168));
  nona23aa1n03x5               g073(.a(new_n165), .b(new_n157), .c(new_n156), .d(new_n164), .out0(new_n169));
  nor042aa1n06x5               g074(.a(new_n169), .b(new_n152), .o1(new_n170));
  nona23aa1n06x5               g075(.a(new_n137), .b(new_n170), .c(new_n147), .d(new_n99), .out0(new_n171));
  nor022aa1n12x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n03x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n171), .c(new_n168), .out0(\s[15] ));
  inv000aa1d42x5               g080(.a(new_n172), .o1(new_n176));
  inv000aa1n02x5               g081(.a(new_n174), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n176), .b(new_n177), .c(new_n171), .d(new_n168), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor022aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  tech160nm_finand02aa1n05x5   g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  aoi012aa1d18x5               g086(.a(new_n180), .b(new_n172), .c(new_n181), .o1(new_n182));
  nano23aa1n03x5               g087(.a(new_n172), .b(new_n180), .c(new_n181), .d(new_n173), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n167), .c(new_n154), .d(new_n166), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n166), .b(new_n150), .o1(new_n185));
  nano32aa1n03x7               g090(.a(new_n185), .b(new_n183), .c(new_n100), .d(new_n128), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n127), .c(new_n114), .d(new_n122), .o1(new_n187));
  nanp03aa1d12x5               g092(.a(new_n187), .b(new_n184), .c(new_n182), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g094(.a(\a[18] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\a[17] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[16] ), .o1(new_n192));
  oaoi03aa1n03x5               g097(.a(new_n191), .b(new_n192), .c(new_n188), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[17] ), .c(new_n190), .out0(\s[18] ));
  inv020aa1n04x5               g099(.a(new_n153), .o1(new_n195));
  aoai13aa1n04x5               g100(.a(new_n166), .b(new_n195), .c(new_n150), .d(new_n139), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n167), .o1(new_n197));
  nona23aa1n09x5               g102(.a(new_n181), .b(new_n173), .c(new_n172), .d(new_n180), .out0(new_n198));
  aoai13aa1n06x5               g103(.a(new_n182), .b(new_n198), .c(new_n196), .d(new_n197), .o1(new_n199));
  nona32aa1n09x5               g104(.a(new_n170), .b(new_n198), .c(new_n147), .d(new_n99), .out0(new_n200));
  oaoi13aa1n12x5               g105(.a(new_n200), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n201));
  xroi22aa1d04x5               g106(.a(new_n191), .b(\b[16] ), .c(new_n190), .d(\b[17] ), .out0(new_n202));
  oaih12aa1n02x5               g107(.a(new_n202), .b(new_n199), .c(new_n201), .o1(new_n203));
  oai022aa1d24x5               g108(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n204));
  oaib12aa1n18x5               g109(.a(new_n204), .b(new_n190), .c(\b[17] ), .out0(new_n205));
  xnrc02aa1n12x5               g110(.a(\b[18] ), .b(\a[19] ), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n203), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  tech160nm_fiaoi012aa1n02p5x5 g116(.a(new_n206), .b(new_n203), .c(new_n205), .o1(new_n212));
  xnrc02aa1n12x5               g117(.a(\b[19] ), .b(\a[20] ), .out0(new_n213));
  nano22aa1n02x4               g118(.a(new_n212), .b(new_n211), .c(new_n213), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n205), .o1(new_n215));
  aoai13aa1n04x5               g120(.a(new_n207), .b(new_n215), .c(new_n188), .d(new_n202), .o1(new_n216));
  tech160nm_fiaoi012aa1n04x5   g121(.a(new_n213), .b(new_n216), .c(new_n211), .o1(new_n217));
  norp02aa1n03x5               g122(.a(new_n217), .b(new_n214), .o1(\s[20] ));
  nor042aa1n03x5               g123(.a(new_n213), .b(new_n206), .o1(new_n219));
  and002aa1n02x5               g124(.a(new_n202), .b(new_n219), .o(new_n220));
  oaih12aa1n02x5               g125(.a(new_n220), .b(new_n199), .c(new_n201), .o1(new_n221));
  oao003aa1n02x5               g126(.a(\a[20] ), .b(\b[19] ), .c(new_n211), .carry(new_n222));
  oai013aa1d12x5               g127(.a(new_n222), .b(new_n206), .c(new_n213), .d(new_n205), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  xorc02aa1n12x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n221), .c(new_n224), .out0(\s[21] ));
  orn002aa1n24x5               g131(.a(\a[21] ), .b(\b[20] ), .o(new_n227));
  inv000aa1d42x5               g132(.a(new_n225), .o1(new_n228));
  aoi012aa1n03x5               g133(.a(new_n228), .b(new_n221), .c(new_n224), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[21] ), .b(\a[22] ), .out0(new_n230));
  nano22aa1n02x4               g135(.a(new_n229), .b(new_n227), .c(new_n230), .out0(new_n231));
  aoai13aa1n02x5               g136(.a(new_n225), .b(new_n223), .c(new_n188), .d(new_n220), .o1(new_n232));
  tech160nm_fiaoi012aa1n02p5x5 g137(.a(new_n230), .b(new_n232), .c(new_n227), .o1(new_n233));
  norp02aa1n02x5               g138(.a(new_n233), .b(new_n231), .o1(\s[22] ));
  norb02aa1n02x5               g139(.a(new_n225), .b(new_n230), .out0(new_n235));
  oao003aa1n12x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n227), .carry(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi012aa1n09x5               g142(.a(new_n237), .b(new_n223), .c(new_n235), .o1(new_n238));
  and003aa1n02x5               g143(.a(new_n235), .b(new_n219), .c(new_n202), .o(new_n239));
  tech160nm_fioai012aa1n03p5x5 g144(.a(new_n239), .b(new_n199), .c(new_n201), .o1(new_n240));
  xorc02aa1n12x5               g145(.a(\a[23] ), .b(\b[22] ), .out0(new_n241));
  xnbna2aa1n03x5               g146(.a(new_n241), .b(new_n240), .c(new_n238), .out0(\s[23] ));
  nor042aa1n06x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n241), .o1(new_n245));
  tech160nm_fiaoi012aa1n02p5x5 g150(.a(new_n245), .b(new_n240), .c(new_n238), .o1(new_n246));
  xorc02aa1n12x5               g151(.a(\a[24] ), .b(\b[23] ), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  nano22aa1n03x5               g153(.a(new_n246), .b(new_n244), .c(new_n248), .out0(new_n249));
  inv040aa1n02x5               g154(.a(new_n238), .o1(new_n250));
  aoai13aa1n03x5               g155(.a(new_n241), .b(new_n250), .c(new_n188), .d(new_n239), .o1(new_n251));
  tech160nm_fiaoi012aa1n02p5x5 g156(.a(new_n248), .b(new_n251), .c(new_n244), .o1(new_n252));
  norp02aa1n02x5               g157(.a(new_n252), .b(new_n249), .o1(\s[24] ));
  inv000aa1n02x5               g158(.a(new_n220), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\a[23] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(\a[24] ), .o1(new_n256));
  xroi22aa1d04x5               g161(.a(new_n255), .b(\b[22] ), .c(new_n256), .d(\b[23] ), .out0(new_n257));
  nano22aa1n02x4               g162(.a(new_n254), .b(new_n235), .c(new_n257), .out0(new_n258));
  oaih12aa1n02x5               g163(.a(new_n258), .b(new_n199), .c(new_n201), .o1(new_n259));
  oaoi03aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .c(new_n244), .o1(new_n260));
  aoib12aa1n12x5               g165(.a(new_n260), .b(new_n257), .c(new_n236), .out0(new_n261));
  nano23aa1n06x5               g166(.a(new_n248), .b(new_n230), .c(new_n225), .d(new_n241), .out0(new_n262));
  nand02aa1d08x5               g167(.a(new_n262), .b(new_n223), .o1(new_n263));
  nand02aa1d06x5               g168(.a(new_n263), .b(new_n261), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  xnrc02aa1n12x5               g170(.a(\b[24] ), .b(\a[25] ), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xnbna2aa1n03x5               g172(.a(new_n267), .b(new_n259), .c(new_n265), .out0(\s[25] ));
  nor042aa1n03x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  tech160nm_fiaoi012aa1n02p5x5 g175(.a(new_n266), .b(new_n259), .c(new_n265), .o1(new_n271));
  tech160nm_fixnrc02aa1n04x5   g176(.a(\b[25] ), .b(\a[26] ), .out0(new_n272));
  nano22aa1n03x5               g177(.a(new_n271), .b(new_n270), .c(new_n272), .out0(new_n273));
  aoai13aa1n02x5               g178(.a(new_n267), .b(new_n264), .c(new_n188), .d(new_n258), .o1(new_n274));
  tech160nm_fiaoi012aa1n02p5x5 g179(.a(new_n272), .b(new_n274), .c(new_n270), .o1(new_n275));
  norp02aa1n03x5               g180(.a(new_n275), .b(new_n273), .o1(\s[26] ));
  nor002aa1n03x5               g181(.a(new_n272), .b(new_n266), .o1(new_n277));
  inv020aa1n02x5               g182(.a(new_n277), .o1(new_n278));
  nano32aa1n03x7               g183(.a(new_n278), .b(new_n262), .c(new_n219), .d(new_n202), .out0(new_n279));
  oai012aa1n06x5               g184(.a(new_n279), .b(new_n199), .c(new_n201), .o1(new_n280));
  oao003aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .c(new_n270), .carry(new_n281));
  aobi12aa1n12x5               g186(.a(new_n281), .b(new_n264), .c(new_n277), .out0(new_n282));
  nor002aa1d32x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  nanp02aa1n04x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  nanb02aa1n12x5               g189(.a(new_n283), .b(new_n284), .out0(new_n285));
  xobna2aa1n03x5               g190(.a(new_n285), .b(new_n280), .c(new_n282), .out0(\s[27] ));
  inv000aa1d42x5               g191(.a(new_n283), .o1(new_n287));
  xnrc02aa1n12x5               g192(.a(\b[27] ), .b(\a[28] ), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n281), .b(new_n278), .c(new_n263), .d(new_n261), .o1(new_n289));
  aoai13aa1n02x5               g194(.a(new_n284), .b(new_n289), .c(new_n188), .d(new_n279), .o1(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n288), .b(new_n290), .c(new_n287), .o1(new_n291));
  aoi022aa1n02x7               g196(.a(new_n280), .b(new_n282), .c(\b[26] ), .d(\a[27] ), .o1(new_n292));
  nano22aa1n03x5               g197(.a(new_n292), .b(new_n287), .c(new_n288), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[28] ));
  nor042aa1n04x5               g199(.a(new_n288), .b(new_n285), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n289), .c(new_n188), .d(new_n279), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n297));
  xnrc02aa1n12x5               g202(.a(\b[28] ), .b(\a[29] ), .out0(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n298), .b(new_n296), .c(new_n297), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n295), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n280), .c(new_n282), .o1(new_n301));
  nano22aa1n03x5               g206(.a(new_n301), .b(new_n297), .c(new_n298), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n299), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n111), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nor043aa1n03x5               g209(.a(new_n298), .b(new_n288), .c(new_n285), .o1(new_n305));
  aoai13aa1n06x5               g210(.a(new_n305), .b(new_n289), .c(new_n188), .d(new_n279), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n305), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n310), .b(new_n280), .c(new_n282), .o1(new_n311));
  nano22aa1n03x5               g216(.a(new_n311), .b(new_n307), .c(new_n308), .out0(new_n312));
  norp02aa1n03x5               g217(.a(new_n309), .b(new_n312), .o1(\s[30] ));
  xnrc02aa1n02x5               g218(.a(\b[30] ), .b(\a[31] ), .out0(new_n314));
  norb03aa1d15x5               g219(.a(new_n295), .b(new_n308), .c(new_n298), .out0(new_n315));
  inv000aa1d42x5               g220(.a(new_n315), .o1(new_n316));
  tech160nm_fiaoi012aa1n03p5x5 g221(.a(new_n316), .b(new_n280), .c(new_n282), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n318));
  nano22aa1n03x5               g223(.a(new_n317), .b(new_n314), .c(new_n318), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n315), .b(new_n289), .c(new_n188), .d(new_n279), .o1(new_n320));
  tech160nm_fiaoi012aa1n02p5x5 g225(.a(new_n314), .b(new_n320), .c(new_n318), .o1(new_n321));
  norp02aa1n03x5               g226(.a(new_n321), .b(new_n319), .o1(\s[31] ));
  xnrb03aa1n02x5               g227(.a(new_n112), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g228(.a(\a[3] ), .b(\b[2] ), .c(new_n112), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g230(.a(new_n114), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g231(.a(\a[5] ), .b(\b[4] ), .c(new_n133), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n03x5               g233(.a(new_n115), .b(new_n327), .out0(new_n329));
  oaib12aa1n06x5               g234(.a(new_n329), .b(\a[6] ), .c(new_n123), .out0(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  inv000aa1d42x5               g236(.a(\a[8] ), .o1(new_n332));
  aoi012aa1n03x5               g237(.a(new_n118), .b(new_n330), .c(new_n119), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[7] ), .c(new_n332), .out0(\s[8] ));
  xorb03aa1n02x5               g239(.a(new_n137), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


