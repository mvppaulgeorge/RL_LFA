// Benchmark "adder" written by ABC on Thu Jul 18 03:28:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n321, new_n322, new_n325, new_n327,
    new_n328, new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor042aa1d18x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor002aa1n16x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(new_n101), .o1(new_n102));
  nand42aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  aob012aa1n06x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .out0(new_n105));
  norb02aa1n09x5               g010(.a(new_n103), .b(new_n101), .out0(new_n106));
  nand22aa1n04x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  nand42aa1n06x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nor042aa1n02x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  nona22aa1n09x5               g014(.a(new_n108), .b(new_n109), .c(new_n107), .out0(new_n110));
  nand42aa1n04x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nano22aa1n12x5               g016(.a(new_n104), .b(new_n108), .c(new_n111), .out0(new_n112));
  aoi013aa1n09x5               g017(.a(new_n105), .b(new_n112), .c(new_n110), .d(new_n106), .o1(new_n113));
  nor002aa1n03x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand42aa1n08x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor002aa1n04x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nano23aa1n03x7               g022(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n118));
  tech160nm_fixorc02aa1n03p5x5 g023(.a(\a[8] ), .b(\b[7] ), .out0(new_n119));
  tech160nm_fixorc02aa1n04x5   g024(.a(\a[7] ), .b(\b[6] ), .out0(new_n120));
  nand23aa1n03x5               g025(.a(new_n118), .b(new_n119), .c(new_n120), .o1(new_n121));
  nor042aa1n06x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(new_n122), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[8] ), .b(\b[7] ), .c(new_n123), .o1(new_n124));
  oa0012aa1n02x5               g029(.a(new_n115), .b(new_n116), .c(new_n114), .o(new_n125));
  aoi013aa1n06x4               g030(.a(new_n124), .b(new_n125), .c(new_n119), .d(new_n120), .o1(new_n126));
  tech160nm_fioai012aa1n05x5   g031(.a(new_n126), .b(new_n113), .c(new_n121), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  aoai13aa1n06x5               g033(.a(new_n99), .b(new_n100), .c(new_n127), .d(new_n128), .o1(new_n129));
  aoi112aa1n02x5               g034(.a(new_n99), .b(new_n100), .c(new_n127), .d(new_n128), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(\s[10] ));
  inv000aa1n03x5               g036(.a(new_n100), .o1(new_n132));
  oaoi03aa1n12x5               g037(.a(\a[10] ), .b(\b[9] ), .c(new_n132), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nor002aa1n06x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand22aa1n03x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  xobna2aa1n03x5               g042(.a(new_n137), .b(new_n129), .c(new_n134), .out0(\s[11] ));
  tech160nm_fiao0012aa1n02p5x5 g043(.a(new_n137), .b(new_n129), .c(new_n134), .o(new_n139));
  norp02aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1n02x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  aoib12aa1n02x5               g047(.a(new_n135), .b(new_n141), .c(new_n140), .out0(new_n143));
  inv000aa1n02x5               g048(.a(new_n135), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n137), .c(new_n129), .d(new_n134), .o1(new_n145));
  aoi022aa1n02x5               g050(.a(new_n139), .b(new_n143), .c(new_n145), .d(new_n142), .o1(\s[12] ));
  nona23aa1n03x5               g051(.a(new_n141), .b(new_n136), .c(new_n135), .d(new_n140), .out0(new_n147));
  nona23aa1n02x4               g052(.a(new_n128), .b(new_n98), .c(new_n97), .d(new_n100), .out0(new_n148));
  norp02aa1n02x5               g053(.a(new_n148), .b(new_n147), .o1(new_n149));
  oaoi03aa1n02x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n150));
  oabi12aa1n02x5               g055(.a(new_n150), .b(new_n134), .c(new_n147), .out0(new_n151));
  tech160nm_fiao0012aa1n03p5x5 g056(.a(new_n151), .b(new_n127), .c(new_n149), .o(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  xnrc02aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .out0(new_n154));
  nanb02aa1n03x5               g059(.a(new_n154), .b(new_n152), .out0(new_n155));
  xnrc02aa1n12x5               g060(.a(\b[13] ), .b(\a[14] ), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  norp02aa1n02x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  norb02aa1n02x5               g063(.a(new_n156), .b(new_n158), .out0(new_n159));
  oai012aa1n02x5               g064(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .o1(new_n160));
  aoi022aa1n02x5               g065(.a(new_n160), .b(new_n157), .c(new_n155), .d(new_n159), .o1(\s[14] ));
  nor042aa1n04x5               g066(.a(new_n156), .b(new_n154), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n151), .c(new_n127), .d(new_n149), .o1(new_n163));
  norp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  aoi012aa1n02x5               g070(.a(new_n164), .b(new_n158), .c(new_n165), .o1(new_n166));
  norp02aa1n12x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n12x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n163), .c(new_n166), .out0(\s[15] ));
  aob012aa1n03x5               g075(.a(new_n169), .b(new_n163), .c(new_n166), .out0(new_n171));
  norp02aa1n04x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand42aa1n16x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  aoib12aa1n02x5               g079(.a(new_n167), .b(new_n173), .c(new_n172), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n167), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n169), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n176), .b(new_n177), .c(new_n163), .d(new_n166), .o1(new_n178));
  aoi022aa1n03x5               g083(.a(new_n178), .b(new_n174), .c(new_n171), .d(new_n175), .o1(\s[16] ));
  nano23aa1d15x5               g084(.a(new_n167), .b(new_n172), .c(new_n173), .d(new_n168), .out0(new_n180));
  nona23aa1n09x5               g085(.a(new_n162), .b(new_n180), .c(new_n148), .d(new_n147), .out0(new_n181));
  inv030aa1n02x5               g086(.a(new_n181), .o1(new_n182));
  nanp02aa1n03x5               g087(.a(new_n127), .b(new_n182), .o1(new_n183));
  nano23aa1n02x4               g088(.a(new_n135), .b(new_n140), .c(new_n141), .d(new_n136), .out0(new_n184));
  aoai13aa1n03x5               g089(.a(new_n162), .b(new_n150), .c(new_n184), .d(new_n133), .o1(new_n185));
  aob012aa1n06x5               g090(.a(new_n180), .b(new_n185), .c(new_n166), .out0(new_n186));
  aoi012aa1n02x5               g091(.a(new_n172), .b(new_n167), .c(new_n173), .o1(new_n187));
  nand23aa1n06x5               g092(.a(new_n183), .b(new_n186), .c(new_n187), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  nanb02aa1n02x5               g095(.a(\b[16] ), .b(new_n190), .out0(new_n191));
  oaoi13aa1n12x5               g096(.a(new_n181), .b(new_n126), .c(new_n113), .d(new_n121), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n180), .o1(new_n193));
  aoai13aa1n06x5               g098(.a(new_n187), .b(new_n193), .c(new_n185), .d(new_n166), .o1(new_n194));
  xorc02aa1n02x5               g099(.a(\a[17] ), .b(\b[16] ), .out0(new_n195));
  oaih12aa1n02x5               g100(.a(new_n195), .b(new_n194), .c(new_n192), .o1(new_n196));
  tech160nm_fixorc02aa1n05x5   g101(.a(\a[18] ), .b(\b[17] ), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n196), .c(new_n191), .out0(\s[18] ));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  xroi22aa1d04x5               g104(.a(new_n190), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n200));
  oaih12aa1n02x5               g105(.a(new_n200), .b(new_n194), .c(new_n192), .o1(new_n201));
  oai022aa1n02x5               g106(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n202));
  oaib12aa1n09x5               g107(.a(new_n202), .b(new_n199), .c(\b[17] ), .out0(new_n203));
  nor042aa1n06x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanp02aa1n04x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  norb02aa1n02x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n201), .c(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n191), .o1(new_n209));
  aoai13aa1n03x5               g114(.a(new_n206), .b(new_n209), .c(new_n188), .d(new_n200), .o1(new_n210));
  nor022aa1n06x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nanp02aa1n04x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  aoib12aa1n02x5               g118(.a(new_n204), .b(new_n212), .c(new_n211), .out0(new_n214));
  inv000aa1n02x5               g119(.a(new_n204), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n206), .o1(new_n216));
  aoai13aa1n02x5               g121(.a(new_n215), .b(new_n216), .c(new_n201), .d(new_n203), .o1(new_n217));
  aoi022aa1n03x5               g122(.a(new_n217), .b(new_n213), .c(new_n210), .d(new_n214), .o1(\s[20] ));
  nano23aa1n06x5               g123(.a(new_n204), .b(new_n211), .c(new_n212), .d(new_n205), .out0(new_n219));
  nand23aa1n04x5               g124(.a(new_n219), .b(new_n195), .c(new_n197), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  oaih12aa1n02x5               g126(.a(new_n221), .b(new_n194), .c(new_n192), .o1(new_n222));
  nona23aa1n06x5               g127(.a(new_n212), .b(new_n205), .c(new_n204), .d(new_n211), .out0(new_n223));
  oaoi03aa1n03x5               g128(.a(\a[20] ), .b(\b[19] ), .c(new_n215), .o1(new_n224));
  oabi12aa1n18x5               g129(.a(new_n224), .b(new_n223), .c(new_n203), .out0(new_n225));
  inv000aa1d42x5               g130(.a(new_n225), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  xnbna2aa1n03x5               g133(.a(new_n228), .b(new_n222), .c(new_n226), .out0(\s[21] ));
  aoai13aa1n03x5               g134(.a(new_n228), .b(new_n225), .c(new_n188), .d(new_n221), .o1(new_n230));
  xnrc02aa1n12x5               g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  nor042aa1n06x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n231), .b(new_n233), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n233), .o1(new_n235));
  aoai13aa1n02x5               g140(.a(new_n235), .b(new_n227), .c(new_n222), .d(new_n226), .o1(new_n236));
  aoi022aa1n03x5               g141(.a(new_n236), .b(new_n232), .c(new_n230), .d(new_n234), .o1(\s[22] ));
  nor042aa1n06x5               g142(.a(new_n231), .b(new_n227), .o1(new_n238));
  norb02aa1n03x5               g143(.a(new_n238), .b(new_n220), .out0(new_n239));
  oaih12aa1n02x5               g144(.a(new_n239), .b(new_n194), .c(new_n192), .o1(new_n240));
  oao003aa1n12x5               g145(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .carry(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  aoi012aa1n12x5               g147(.a(new_n242), .b(new_n225), .c(new_n238), .o1(new_n243));
  nanp02aa1n02x5               g148(.a(new_n240), .b(new_n243), .o1(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  aoi112aa1n02x5               g150(.a(new_n245), .b(new_n242), .c(new_n225), .d(new_n238), .o1(new_n246));
  aoi022aa1n02x5               g151(.a(new_n244), .b(new_n245), .c(new_n240), .d(new_n246), .o1(\s[23] ));
  inv000aa1d42x5               g152(.a(new_n243), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n245), .b(new_n248), .c(new_n188), .d(new_n239), .o1(new_n249));
  tech160nm_fixorc02aa1n04x5   g154(.a(\a[24] ), .b(\b[23] ), .out0(new_n250));
  nor042aa1n03x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  norp02aa1n02x5               g156(.a(new_n250), .b(new_n251), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n251), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n245), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n253), .b(new_n254), .c(new_n240), .d(new_n243), .o1(new_n255));
  aoi022aa1n03x5               g160(.a(new_n255), .b(new_n250), .c(new_n249), .d(new_n252), .o1(\s[24] ));
  nano32aa1d12x5               g161(.a(new_n220), .b(new_n250), .c(new_n238), .d(new_n245), .out0(new_n257));
  oaih12aa1n02x5               g162(.a(new_n257), .b(new_n194), .c(new_n192), .o1(new_n258));
  aoai13aa1n06x5               g163(.a(new_n238), .b(new_n224), .c(new_n219), .d(new_n209), .o1(new_n259));
  and002aa1n06x5               g164(.a(new_n250), .b(new_n245), .o(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  oao003aa1n02x5               g166(.a(\a[24] ), .b(\b[23] ), .c(new_n253), .carry(new_n262));
  aoai13aa1n12x5               g167(.a(new_n262), .b(new_n261), .c(new_n259), .d(new_n241), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  xorc02aa1n12x5               g169(.a(\a[25] ), .b(\b[24] ), .out0(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n258), .c(new_n264), .out0(\s[25] ));
  aoai13aa1n03x5               g171(.a(new_n265), .b(new_n263), .c(new_n188), .d(new_n257), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  nor042aa1n03x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  norp02aa1n02x5               g174(.a(new_n268), .b(new_n269), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n269), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n265), .o1(new_n272));
  aoai13aa1n02x5               g177(.a(new_n271), .b(new_n272), .c(new_n258), .d(new_n264), .o1(new_n273));
  aoi022aa1n03x5               g178(.a(new_n273), .b(new_n268), .c(new_n267), .d(new_n270), .o1(\s[26] ));
  and002aa1n06x5               g179(.a(new_n268), .b(new_n265), .o(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  nano23aa1d12x5               g181(.a(new_n276), .b(new_n220), .c(new_n260), .d(new_n238), .out0(new_n277));
  oai012aa1n06x5               g182(.a(new_n277), .b(new_n194), .c(new_n192), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  aoi012aa1n12x5               g185(.a(new_n280), .b(new_n263), .c(new_n275), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n278), .c(new_n281), .out0(\s[27] ));
  aoai13aa1n06x5               g188(.a(new_n260), .b(new_n242), .c(new_n225), .d(new_n238), .o1(new_n284));
  aoai13aa1n04x5               g189(.a(new_n279), .b(new_n276), .c(new_n284), .d(new_n262), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n282), .b(new_n285), .c(new_n188), .d(new_n277), .o1(new_n286));
  tech160nm_fixorc02aa1n04x5   g191(.a(\a[28] ), .b(\b[27] ), .out0(new_n287));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  norp02aa1n02x5               g193(.a(new_n287), .b(new_n288), .o1(new_n289));
  inv000aa1n03x5               g194(.a(new_n288), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n282), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n290), .b(new_n291), .c(new_n278), .d(new_n281), .o1(new_n292));
  aoi022aa1n03x5               g197(.a(new_n292), .b(new_n287), .c(new_n286), .d(new_n289), .o1(\s[28] ));
  and002aa1n02x5               g198(.a(new_n287), .b(new_n282), .o(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n285), .c(new_n188), .d(new_n277), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n294), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n290), .carry(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n296), .c(new_n278), .d(new_n281), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  norb02aa1n02x5               g204(.a(new_n297), .b(new_n299), .out0(new_n300));
  aoi022aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n295), .d(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g206(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g207(.a(new_n291), .b(new_n287), .c(new_n299), .out0(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n285), .c(new_n188), .d(new_n277), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n303), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n305), .c(new_n278), .d(new_n281), .o1(new_n307));
  xorc02aa1n02x5               g212(.a(\a[30] ), .b(\b[29] ), .out0(new_n308));
  norb02aa1n02x5               g213(.a(new_n306), .b(new_n308), .out0(new_n309));
  aoi022aa1n03x5               g214(.a(new_n307), .b(new_n308), .c(new_n304), .d(new_n309), .o1(\s[30] ));
  nano32aa1n02x4               g215(.a(new_n291), .b(new_n308), .c(new_n287), .d(new_n299), .out0(new_n311));
  aoai13aa1n04x5               g216(.a(new_n311), .b(new_n285), .c(new_n188), .d(new_n277), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[31] ), .b(\b[30] ), .out0(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n314));
  norb02aa1n02x5               g219(.a(new_n314), .b(new_n313), .out0(new_n315));
  inv000aa1n02x5               g220(.a(new_n311), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n314), .b(new_n316), .c(new_n278), .d(new_n281), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n312), .d(new_n315), .o1(\s[31] ));
  norb02aa1n02x5               g223(.a(new_n111), .b(new_n104), .out0(new_n319));
  xobna2aa1n03x5               g224(.a(new_n319), .b(new_n110), .c(new_n108), .out0(\s[3] ));
  oai112aa1n02x5               g225(.a(new_n319), .b(new_n108), .c(new_n109), .d(new_n107), .o1(new_n321));
  aoi012aa1n02x5               g226(.a(new_n104), .b(new_n102), .c(new_n103), .o1(new_n322));
  aboi22aa1n03x5               g227(.a(new_n113), .b(new_n102), .c(new_n322), .d(new_n321), .out0(\s[4] ));
  xnrb03aa1n02x5               g228(.a(new_n113), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g229(.a(\a[5] ), .b(\b[4] ), .c(new_n113), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g231(.a(new_n113), .o1(new_n327));
  aoai13aa1n02x5               g232(.a(new_n120), .b(new_n125), .c(new_n327), .d(new_n118), .o1(new_n328));
  aoi112aa1n02x5               g233(.a(new_n125), .b(new_n120), .c(new_n327), .d(new_n118), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n328), .b(new_n329), .out0(\s[7] ));
  xnbna2aa1n03x5               g235(.a(new_n119), .b(new_n328), .c(new_n123), .out0(\s[8] ));
  xorb03aa1n02x5               g236(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


