// Benchmark "adder" written by ABC on Thu Jul 18 12:31:11 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n355, new_n356, new_n358, new_n361,
    new_n362, new_n363, new_n365, new_n366, new_n367, new_n369, new_n371,
    new_n372;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[1] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[0] ), .o1(new_n98));
  norp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oaoi13aa1n02x5               g005(.a(new_n99), .b(new_n100), .c(new_n97), .d(new_n98), .o1(new_n101));
  norp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n02x4               g010(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n106));
  tech160nm_fioai012aa1n04x5   g011(.a(new_n103), .b(new_n104), .c(new_n102), .o1(new_n107));
  tech160nm_fioai012aa1n05x5   g012(.a(new_n107), .b(new_n106), .c(new_n101), .o1(new_n108));
  norp02aa1n04x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  norp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nona23aa1n02x4               g017(.a(new_n111), .b(new_n110), .c(new_n112), .d(new_n109), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  nor043aa1n02x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[8] ), .o1(new_n117));
  oai022aa1n02x5               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  aoi022aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n119));
  aoai13aa1n02x5               g024(.a(new_n111), .b(new_n109), .c(new_n118), .d(new_n119), .o1(new_n120));
  oaib12aa1n02x5               g025(.a(new_n120), .b(\b[7] ), .c(new_n117), .out0(new_n121));
  nor002aa1n02x5               g026(.a(\b[8] ), .b(\a[9] ), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(\b[8] ), .b(\a[9] ), .o1(new_n123));
  norb02aa1n02x5               g028(.a(new_n123), .b(new_n122), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n125));
  oai012aa1n02x5               g030(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand42aa1n03x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nor042aa1n02x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  norp02aa1n02x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nona22aa1n02x4               g037(.a(new_n125), .b(new_n122), .c(new_n132), .out0(new_n133));
  xobna2aa1n03x5               g038(.a(new_n131), .b(new_n133), .c(new_n128), .out0(\s[11] ));
  norp02aa1n02x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nand42aa1n03x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  nano22aa1n02x4               g042(.a(new_n129), .b(new_n128), .c(new_n130), .out0(new_n138));
  aoi012aa1n02x5               g043(.a(new_n129), .b(new_n133), .c(new_n138), .o1(new_n139));
  norb03aa1n02x5               g044(.a(new_n136), .b(new_n129), .c(new_n135), .out0(new_n140));
  aob012aa1n02x5               g045(.a(new_n140), .b(new_n133), .c(new_n138), .out0(new_n141));
  oai012aa1n02x5               g046(.a(new_n141), .b(new_n139), .c(new_n137), .o1(\s[12] ));
  nano23aa1n03x5               g047(.a(new_n132), .b(new_n135), .c(new_n136), .d(new_n128), .out0(new_n143));
  nano23aa1n03x5               g048(.a(new_n122), .b(new_n129), .c(new_n130), .d(new_n123), .out0(new_n144));
  nand02aa1d06x5               g049(.a(new_n144), .b(new_n143), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  aoai13aa1n02x5               g051(.a(new_n146), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n147));
  aoi022aa1n02x5               g052(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n148));
  oai012aa1n02x5               g053(.a(new_n148), .b(new_n122), .c(new_n132), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n140), .b(new_n149), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n150), .b(new_n136), .o1(new_n151));
  nor022aa1n06x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1n03x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  norb02aa1n02x5               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  xnbna2aa1n03x5               g059(.a(new_n154), .b(new_n147), .c(new_n151), .out0(\s[13] ));
  nand42aa1n03x5               g060(.a(new_n147), .b(new_n151), .o1(new_n156));
  nor022aa1n04x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand42aa1n03x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n157), .b(new_n158), .out0(new_n159));
  aoai13aa1n02x5               g064(.a(new_n159), .b(new_n152), .c(new_n156), .d(new_n153), .o1(new_n160));
  nona22aa1n02x4               g065(.a(new_n158), .b(new_n157), .c(new_n152), .out0(new_n161));
  aoai13aa1n02x5               g066(.a(new_n160), .b(new_n161), .c(new_n154), .d(new_n156), .o1(\s[14] ));
  nano23aa1n02x5               g067(.a(new_n152), .b(new_n157), .c(new_n158), .d(new_n153), .out0(new_n163));
  oa0012aa1n02x5               g068(.a(new_n158), .b(new_n157), .c(new_n152), .o(new_n164));
  xorc02aa1n02x5               g069(.a(\a[15] ), .b(\b[14] ), .out0(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n164), .c(new_n156), .d(new_n163), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n165), .b(new_n164), .c(new_n156), .d(new_n163), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(\s[15] ));
  inv000aa1d42x5               g073(.a(\a[15] ), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\b[14] ), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(new_n170), .b(new_n169), .o1(new_n171));
  nor002aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  and002aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o(new_n173));
  norp02aa1n02x5               g078(.a(new_n173), .b(new_n172), .o1(new_n174));
  oai022aa1n02x5               g079(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n175));
  nona22aa1n02x4               g080(.a(new_n166), .b(new_n173), .c(new_n175), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n174), .c(new_n171), .d(new_n166), .o1(\s[16] ));
  nano32aa1n03x7               g082(.a(new_n145), .b(new_n174), .c(new_n163), .d(new_n165), .out0(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n179));
  aoi112aa1n02x5               g084(.a(new_n173), .b(new_n172), .c(\a[15] ), .d(\b[14] ), .o1(new_n180));
  oai012aa1n02x5               g085(.a(new_n136), .b(\b[12] ), .c(\a[13] ), .o1(new_n181));
  nano23aa1n02x4               g086(.a(new_n159), .b(new_n181), .c(new_n171), .d(new_n153), .out0(new_n182));
  oai122aa1n02x7               g087(.a(new_n158), .b(new_n157), .c(new_n152), .d(new_n170), .e(new_n169), .o1(new_n183));
  aoi022aa1n02x5               g088(.a(new_n183), .b(new_n171), .c(\a[16] ), .d(\b[15] ), .o1(new_n184));
  aoi113aa1n06x5               g089(.a(new_n172), .b(new_n184), .c(new_n182), .d(new_n180), .e(new_n150), .o1(new_n185));
  nand42aa1n06x5               g090(.a(new_n179), .b(new_n185), .o1(new_n186));
  nor042aa1n06x5               g091(.a(\b[16] ), .b(\a[17] ), .o1(new_n187));
  nand42aa1n03x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  norb02aa1n02x5               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  obai22aa1n02x7               g094(.a(new_n188), .b(new_n187), .c(\a[16] ), .d(\b[15] ), .out0(new_n190));
  aoi113aa1n02x5               g095(.a(new_n190), .b(new_n184), .c(new_n182), .d(new_n180), .e(new_n150), .o1(new_n191));
  aoi022aa1n02x5               g096(.a(new_n186), .b(new_n189), .c(new_n179), .d(new_n191), .o1(\s[17] ));
  inv000aa1d42x5               g097(.a(new_n187), .o1(new_n193));
  and002aa1n02x5               g098(.a(\b[0] ), .b(\a[1] ), .o(new_n194));
  oaoi03aa1n02x5               g099(.a(\a[2] ), .b(\b[1] ), .c(new_n194), .o1(new_n195));
  norb02aa1n06x4               g100(.a(new_n103), .b(new_n102), .out0(new_n196));
  norb02aa1n02x5               g101(.a(new_n105), .b(new_n104), .out0(new_n197));
  nanp03aa1n02x5               g102(.a(new_n195), .b(new_n196), .c(new_n197), .o1(new_n198));
  nano23aa1n02x4               g103(.a(new_n112), .b(new_n109), .c(new_n110), .d(new_n111), .out0(new_n199));
  xorc02aa1n02x5               g104(.a(\a[5] ), .b(\b[4] ), .out0(new_n200));
  xorc02aa1n02x5               g105(.a(\a[6] ), .b(\b[5] ), .out0(new_n201));
  nanp03aa1n02x5               g106(.a(new_n199), .b(new_n200), .c(new_n201), .o1(new_n202));
  norp02aa1n02x5               g107(.a(\b[4] ), .b(\a[5] ), .o1(new_n203));
  norp02aa1n02x5               g108(.a(\b[5] ), .b(\a[6] ), .o1(new_n204));
  oai012aa1n02x5               g109(.a(new_n119), .b(new_n204), .c(new_n203), .o1(new_n205));
  oai012aa1n02x5               g110(.a(new_n205), .b(\b[6] ), .c(\a[7] ), .o1(new_n206));
  aoi012aa1n02x5               g111(.a(new_n112), .b(new_n206), .c(new_n111), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n198), .d(new_n107), .o1(new_n208));
  nanp03aa1n02x5               g113(.a(new_n182), .b(new_n150), .c(new_n180), .o1(new_n209));
  nona22aa1n02x4               g114(.a(new_n209), .b(new_n184), .c(new_n172), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n189), .b(new_n210), .c(new_n208), .d(new_n178), .o1(new_n211));
  nor042aa1n02x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  nand02aa1n03x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  norb02aa1n02x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  oai022aa1n02x5               g119(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n215));
  nanb03aa1n02x5               g120(.a(new_n215), .b(new_n211), .c(new_n213), .out0(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n214), .c(new_n193), .d(new_n211), .o1(\s[18] ));
  nano23aa1d15x5               g122(.a(new_n187), .b(new_n212), .c(new_n213), .d(new_n188), .out0(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  oaoi03aa1n02x5               g124(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n02x7               g126(.a(new_n221), .b(new_n219), .c(new_n179), .d(new_n185), .o1(new_n222));
  norp02aa1n02x5               g127(.a(\b[18] ), .b(\a[19] ), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  aoi112aa1n02x5               g130(.a(new_n225), .b(new_n220), .c(new_n186), .d(new_n218), .o1(new_n226));
  aoi012aa1n02x5               g131(.a(new_n226), .b(new_n222), .c(new_n225), .o1(\s[19] ));
  xnrc02aa1n02x5               g132(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n06x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  nand42aa1n04x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  inv000aa1d42x5               g136(.a(\a[19] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\b[18] ), .o1(new_n233));
  oaoi03aa1n02x5               g138(.a(new_n232), .b(new_n233), .c(new_n222), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(new_n222), .b(new_n225), .o1(new_n235));
  norp02aa1n02x5               g140(.a(new_n229), .b(new_n223), .o1(new_n236));
  nanp03aa1n02x5               g141(.a(new_n235), .b(new_n230), .c(new_n236), .o1(new_n237));
  oaih12aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n231), .o1(\s[20] ));
  nano23aa1n03x7               g143(.a(new_n223), .b(new_n229), .c(new_n230), .d(new_n224), .out0(new_n239));
  nand22aa1n03x5               g144(.a(new_n239), .b(new_n218), .o1(new_n240));
  inv000aa1n06x5               g145(.a(new_n240), .o1(new_n241));
  nanb03aa1n02x5               g146(.a(new_n229), .b(new_n230), .c(new_n224), .out0(new_n242));
  oai112aa1n02x5               g147(.a(new_n215), .b(new_n213), .c(\b[18] ), .d(\a[19] ), .o1(new_n243));
  aoai13aa1n04x5               g148(.a(new_n230), .b(new_n229), .c(new_n232), .d(new_n233), .o1(new_n244));
  tech160nm_fioai012aa1n03p5x5 g149(.a(new_n244), .b(new_n243), .c(new_n242), .o1(new_n245));
  nor002aa1d32x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  nanp02aa1n02x5               g151(.a(\b[20] ), .b(\a[21] ), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n245), .c(new_n186), .d(new_n241), .o1(new_n249));
  nano22aa1n02x4               g154(.a(new_n229), .b(new_n224), .c(new_n230), .out0(new_n250));
  oai012aa1n02x5               g155(.a(new_n213), .b(\b[18] ), .c(\a[19] ), .o1(new_n251));
  oab012aa1n02x4               g156(.a(new_n251), .b(new_n187), .c(new_n212), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n244), .o1(new_n253));
  aoi112aa1n02x5               g158(.a(new_n253), .b(new_n248), .c(new_n252), .d(new_n250), .o1(new_n254));
  aobi12aa1n02x5               g159(.a(new_n254), .b(new_n186), .c(new_n241), .out0(new_n255));
  norb02aa1n02x5               g160(.a(new_n249), .b(new_n255), .out0(\s[21] ));
  inv000aa1d42x5               g161(.a(new_n246), .o1(new_n257));
  nor042aa1n02x5               g162(.a(\b[21] ), .b(\a[22] ), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(\b[21] ), .b(\a[22] ), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n259), .b(new_n258), .out0(new_n260));
  norb03aa1n02x5               g165(.a(new_n259), .b(new_n246), .c(new_n258), .out0(new_n261));
  nand42aa1n03x5               g166(.a(new_n249), .b(new_n261), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n260), .c(new_n257), .d(new_n249), .o1(\s[22] ));
  nano23aa1d15x5               g168(.a(new_n246), .b(new_n258), .c(new_n259), .d(new_n247), .out0(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  nano22aa1n02x4               g170(.a(new_n265), .b(new_n218), .c(new_n239), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n264), .b(new_n253), .c(new_n252), .d(new_n250), .o1(new_n267));
  oaoi03aa1n09x5               g172(.a(\a[22] ), .b(\b[21] ), .c(new_n257), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(new_n267), .b(new_n269), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[23] ), .b(\b[22] ), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n270), .c(new_n186), .d(new_n266), .o1(new_n272));
  nona22aa1n02x4               g177(.a(new_n267), .b(new_n268), .c(new_n271), .out0(new_n273));
  aoi012aa1n02x5               g178(.a(new_n273), .b(new_n186), .c(new_n266), .o1(new_n274));
  norb02aa1n02x5               g179(.a(new_n272), .b(new_n274), .out0(\s[23] ));
  norp02aa1n02x5               g180(.a(\b[22] ), .b(\a[23] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .out0(new_n278));
  oai022aa1n02x5               g183(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n279));
  aoi012aa1n02x5               g184(.a(new_n279), .b(\a[24] ), .c(\b[23] ), .o1(new_n280));
  tech160nm_finand02aa1n03p5x5 g185(.a(new_n272), .b(new_n280), .o1(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n278), .c(new_n277), .d(new_n272), .o1(\s[24] ));
  nano32aa1n02x4               g187(.a(new_n240), .b(new_n278), .c(new_n264), .d(new_n271), .out0(new_n283));
  nanp02aa1n03x5               g188(.a(new_n278), .b(new_n271), .o1(new_n284));
  aob012aa1n02x5               g189(.a(new_n279), .b(\b[23] ), .c(\a[24] ), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n284), .c(new_n267), .d(new_n269), .o1(new_n286));
  xorc02aa1n12x5               g191(.a(\a[25] ), .b(\b[24] ), .out0(new_n287));
  aoai13aa1n06x5               g192(.a(new_n287), .b(new_n286), .c(new_n186), .d(new_n283), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n284), .o1(new_n289));
  aoai13aa1n02x5               g194(.a(new_n289), .b(new_n268), .c(new_n245), .d(new_n264), .o1(new_n290));
  nanb03aa1n02x5               g195(.a(new_n287), .b(new_n290), .c(new_n285), .out0(new_n291));
  aoi012aa1n02x5               g196(.a(new_n291), .b(new_n186), .c(new_n283), .o1(new_n292));
  norb02aa1n02x5               g197(.a(new_n288), .b(new_n292), .out0(\s[25] ));
  norp02aa1n02x5               g198(.a(\b[24] ), .b(\a[25] ), .o1(new_n294));
  inv000aa1n03x5               g199(.a(new_n294), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[26] ), .b(\b[25] ), .out0(new_n296));
  nanp02aa1n02x5               g201(.a(\b[25] ), .b(\a[26] ), .o1(new_n297));
  oai022aa1n02x5               g202(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n298));
  norb02aa1n02x5               g203(.a(new_n297), .b(new_n298), .out0(new_n299));
  tech160nm_finand02aa1n03p5x5 g204(.a(new_n288), .b(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n288), .o1(\s[26] ));
  nanp02aa1n02x5               g206(.a(new_n296), .b(new_n287), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n302), .o1(new_n303));
  nona23aa1n03x5               g208(.a(new_n241), .b(new_n303), .c(new_n284), .d(new_n265), .out0(new_n304));
  inv040aa1n02x5               g209(.a(new_n304), .o1(new_n305));
  aoai13aa1n06x5               g210(.a(new_n305), .b(new_n210), .c(new_n208), .d(new_n178), .o1(new_n306));
  tech160nm_fiaoi012aa1n03p5x5 g211(.a(new_n304), .b(new_n179), .c(new_n185), .o1(new_n307));
  oaoi03aa1n02x5               g212(.a(\a[26] ), .b(\b[25] ), .c(new_n295), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n308), .o1(new_n309));
  aoai13aa1n06x5               g214(.a(new_n309), .b(new_n302), .c(new_n290), .d(new_n285), .o1(new_n310));
  xorc02aa1n12x5               g215(.a(\a[27] ), .b(\b[26] ), .out0(new_n311));
  oaih12aa1n02x5               g216(.a(new_n311), .b(new_n310), .c(new_n307), .o1(new_n312));
  aoi112aa1n02x5               g217(.a(new_n311), .b(new_n308), .c(new_n286), .d(new_n303), .o1(new_n313));
  aobi12aa1n02x5               g218(.a(new_n312), .b(new_n313), .c(new_n306), .out0(\s[27] ));
  norp02aa1n02x5               g219(.a(\b[26] ), .b(\a[27] ), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n315), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[28] ), .b(\b[27] ), .out0(new_n317));
  aoi022aa1n02x7               g222(.a(new_n286), .b(new_n303), .c(new_n297), .d(new_n298), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n311), .o1(new_n319));
  oai022aa1n02x5               g224(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n320));
  aoi012aa1n02x5               g225(.a(new_n320), .b(\a[28] ), .c(\b[27] ), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n319), .c(new_n318), .d(new_n306), .o1(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n317), .c(new_n312), .d(new_n316), .o1(\s[28] ));
  and002aa1n02x5               g228(.a(new_n317), .b(new_n311), .o(new_n324));
  oai012aa1n02x5               g229(.a(new_n324), .b(new_n310), .c(new_n307), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n324), .o1(new_n326));
  aob012aa1n02x5               g231(.a(new_n320), .b(\b[27] ), .c(\a[28] ), .out0(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n326), .c(new_n318), .d(new_n306), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[29] ), .b(\b[28] ), .out0(new_n329));
  norb02aa1n02x5               g234(.a(new_n327), .b(new_n329), .out0(new_n330));
  aoi022aa1n03x5               g235(.a(new_n328), .b(new_n329), .c(new_n325), .d(new_n330), .o1(\s[29] ));
  xnrb03aa1n02x5               g236(.a(new_n194), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g237(.a(new_n319), .b(new_n317), .c(new_n329), .out0(new_n333));
  oaih12aa1n02x5               g238(.a(new_n333), .b(new_n310), .c(new_n307), .o1(new_n334));
  inv000aa1d42x5               g239(.a(new_n333), .o1(new_n335));
  inv000aa1d42x5               g240(.a(\a[29] ), .o1(new_n336));
  inv000aa1d42x5               g241(.a(\b[28] ), .o1(new_n337));
  aoi022aa1n02x5               g242(.a(\b[28] ), .b(\a[29] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n338));
  aoi022aa1n02x5               g243(.a(new_n320), .b(new_n338), .c(new_n337), .d(new_n336), .o1(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n335), .c(new_n318), .d(new_n306), .o1(new_n340));
  xorc02aa1n02x5               g245(.a(\a[30] ), .b(\b[29] ), .out0(new_n341));
  aoi122aa1n02x5               g246(.a(new_n341), .b(new_n320), .c(new_n338), .d(new_n336), .e(new_n337), .o1(new_n342));
  aoi022aa1n02x5               g247(.a(new_n340), .b(new_n341), .c(new_n334), .d(new_n342), .o1(\s[30] ));
  nano32aa1n02x4               g248(.a(new_n319), .b(new_n341), .c(new_n317), .d(new_n329), .out0(new_n344));
  oai012aa1n02x5               g249(.a(new_n344), .b(new_n310), .c(new_n307), .o1(new_n345));
  inv000aa1n02x5               g250(.a(new_n344), .o1(new_n346));
  oao003aa1n02x5               g251(.a(\a[30] ), .b(\b[29] ), .c(new_n339), .carry(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n346), .c(new_n318), .d(new_n306), .o1(new_n348));
  xorc02aa1n02x5               g253(.a(\a[31] ), .b(\b[30] ), .out0(new_n349));
  nanp02aa1n02x5               g254(.a(\b[29] ), .b(\a[30] ), .o1(new_n350));
  oabi12aa1n02x5               g255(.a(new_n349), .b(\a[30] ), .c(\b[29] ), .out0(new_n351));
  aoib12aa1n02x5               g256(.a(new_n351), .b(new_n350), .c(new_n339), .out0(new_n352));
  aoi022aa1n02x5               g257(.a(new_n348), .b(new_n349), .c(new_n345), .d(new_n352), .o1(\s[31] ));
  norb03aa1n02x5               g258(.a(new_n100), .b(new_n194), .c(new_n99), .out0(new_n354));
  inv000aa1d42x5               g259(.a(new_n104), .o1(new_n355));
  aoi012aa1n02x5               g260(.a(new_n99), .b(new_n355), .c(new_n105), .o1(new_n356));
  aboi22aa1n03x5               g261(.a(new_n354), .b(new_n356), .c(new_n195), .d(new_n197), .out0(\s[3] ));
  nanp02aa1n02x5               g262(.a(new_n195), .b(new_n197), .o1(new_n358));
  xnbna2aa1n03x5               g263(.a(new_n196), .b(new_n358), .c(new_n355), .out0(\s[4] ));
  xnbna2aa1n03x5               g264(.a(new_n200), .b(new_n198), .c(new_n107), .out0(\s[5] ));
  aoai13aa1n02x5               g265(.a(new_n115), .b(new_n203), .c(new_n108), .d(new_n200), .o1(new_n361));
  aoi012aa1n02x5               g266(.a(new_n118), .b(\a[6] ), .c(\b[5] ), .o1(new_n362));
  aoai13aa1n02x5               g267(.a(new_n362), .b(new_n114), .c(new_n198), .d(new_n107), .o1(new_n363));
  nanp02aa1n02x5               g268(.a(new_n361), .b(new_n363), .o1(\s[6] ));
  nanb02aa1n02x5               g269(.a(new_n109), .b(new_n110), .out0(new_n365));
  aob012aa1n02x5               g270(.a(new_n363), .b(\b[5] ), .c(\a[6] ), .out0(new_n366));
  norb02aa1n02x5               g271(.a(new_n119), .b(new_n109), .out0(new_n367));
  aoi022aa1n02x5               g272(.a(new_n366), .b(new_n365), .c(new_n363), .d(new_n367), .o1(\s[7] ));
  aoi012aa1n02x5               g273(.a(new_n109), .b(new_n363), .c(new_n119), .o1(new_n369));
  xorb03aa1n02x5               g274(.a(new_n369), .b(\b[7] ), .c(new_n117), .out0(\s[8] ));
  nanp02aa1n02x5               g275(.a(new_n108), .b(new_n116), .o1(new_n371));
  aoi112aa1n02x5               g276(.a(new_n124), .b(new_n112), .c(new_n206), .d(new_n111), .o1(new_n372));
  aoi022aa1n02x5               g277(.a(new_n208), .b(new_n124), .c(new_n371), .d(new_n372), .o1(\s[9] ));
endmodule


