// Benchmark "adder" written by ABC on Wed Jul 17 20:35:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n317,
    new_n318, new_n321, new_n323, new_n325, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  orn002aa1n24x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  xnrc02aa1n02x5               g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nor002aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  tech160nm_fioai012aa1n04x5   g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  inv000aa1d42x5               g008(.a(\a[3] ), .o1(new_n104));
  inv000aa1d42x5               g009(.a(\a[4] ), .o1(new_n105));
  inv000aa1d42x5               g010(.a(\b[2] ), .o1(new_n106));
  aboi22aa1n03x5               g011(.a(\b[3] ), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n107));
  tech160nm_fioai012aa1n04x5   g012(.a(new_n107), .b(new_n99), .c(new_n103), .o1(new_n108));
  nand42aa1n03x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\a[6] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[5] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  oai112aa1n02x5               g017(.a(new_n112), .b(new_n109), .c(\b[6] ), .d(\a[7] ), .o1(new_n113));
  tech160nm_fixorc02aa1n03p5x5 g018(.a(\a[5] ), .b(\b[4] ), .out0(new_n114));
  aoi022aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n115));
  nand02aa1d06x5               g020(.a(\b[3] ), .b(\a[4] ), .o1(new_n116));
  oai112aa1n02x5               g021(.a(new_n115), .b(new_n116), .c(\b[7] ), .d(\a[8] ), .o1(new_n117));
  norb03aa1n03x5               g022(.a(new_n114), .b(new_n113), .c(new_n117), .out0(new_n118));
  nanp02aa1n02x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  oai022aa1n02x7               g024(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  and003aa1n02x5               g026(.a(new_n109), .b(new_n121), .c(new_n119), .o(new_n122));
  nor002aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  aoi012aa1n02x5               g028(.a(new_n123), .b(new_n110), .c(new_n111), .o1(new_n124));
  nona22aa1n02x4               g029(.a(new_n122), .b(new_n124), .c(new_n120), .out0(new_n125));
  aob012aa1n02x5               g030(.a(new_n125), .b(new_n120), .c(new_n119), .out0(new_n126));
  xorc02aa1n02x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n126), .c(new_n118), .d(new_n108), .o1(new_n128));
  xobna2aa1n03x5               g033(.a(new_n97), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  oaoi03aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n97), .c(new_n128), .d(new_n98), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  norp02aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand02aa1n03x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor042aa1n02x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanp02aa1n03x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nanb02aa1n02x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n134), .c(new_n132), .d(new_n135), .o1(new_n139));
  aoi112aa1n02x5               g044(.a(new_n134), .b(new_n138), .c(new_n132), .d(new_n135), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(\s[12] ));
  nona23aa1n09x5               g046(.a(new_n137), .b(new_n135), .c(new_n134), .d(new_n136), .out0(new_n142));
  norb03aa1n02x7               g047(.a(new_n127), .b(new_n142), .c(new_n97), .out0(new_n143));
  aoai13aa1n06x5               g048(.a(new_n143), .b(new_n126), .c(new_n118), .d(new_n108), .o1(new_n144));
  nano23aa1n06x5               g049(.a(new_n134), .b(new_n136), .c(new_n137), .d(new_n135), .out0(new_n145));
  aoi012aa1n02x5               g050(.a(new_n136), .b(new_n134), .c(new_n137), .o1(new_n146));
  aobi12aa1n09x5               g051(.a(new_n146), .b(new_n145), .c(new_n130), .out0(new_n147));
  xorc02aa1n02x5               g052(.a(\a[13] ), .b(\b[12] ), .out0(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n144), .c(new_n147), .out0(\s[13] ));
  orn002aa1n24x5               g054(.a(\a[13] ), .b(\b[12] ), .o(new_n150));
  xorc02aa1n02x5               g055(.a(\a[3] ), .b(\b[2] ), .out0(new_n151));
  nanb02aa1n02x5               g056(.a(new_n103), .b(new_n151), .out0(new_n152));
  oai012aa1n02x5               g057(.a(new_n116), .b(\b[7] ), .c(\a[8] ), .o1(new_n153));
  nano22aa1n02x4               g058(.a(new_n153), .b(new_n119), .c(new_n121), .out0(new_n154));
  nanb03aa1n02x5               g059(.a(new_n113), .b(new_n154), .c(new_n114), .out0(new_n155));
  norp02aa1n02x5               g060(.a(new_n124), .b(new_n120), .o1(new_n156));
  aoi022aa1n02x5               g061(.a(new_n156), .b(new_n122), .c(new_n119), .d(new_n120), .o1(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n155), .c(new_n152), .d(new_n107), .o1(new_n158));
  oaib12aa1n02x5               g063(.a(new_n146), .b(new_n142), .c(new_n130), .out0(new_n159));
  aoai13aa1n02x5               g064(.a(new_n148), .b(new_n159), .c(new_n158), .d(new_n143), .o1(new_n160));
  xorc02aa1n02x5               g065(.a(\a[14] ), .b(\b[13] ), .out0(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n160), .c(new_n150), .out0(\s[14] ));
  xnrc02aa1n03x5               g067(.a(\b[12] ), .b(\a[13] ), .out0(new_n163));
  xnrc02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .out0(new_n164));
  nor042aa1n04x5               g069(.a(new_n164), .b(new_n163), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  oaoi03aa1n09x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n150), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n04x5               g073(.a(new_n168), .b(new_n166), .c(new_n144), .d(new_n147), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  xorc02aa1n02x5               g076(.a(\a[15] ), .b(\b[14] ), .out0(new_n172));
  tech160nm_fixnrc02aa1n04x5   g077(.a(\b[15] ), .b(\a[16] ), .out0(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n171), .c(new_n169), .d(new_n172), .o1(new_n174));
  aoi112aa1n02x5               g079(.a(new_n171), .b(new_n173), .c(new_n169), .d(new_n172), .o1(new_n175));
  nanb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[16] ));
  inv000aa1d42x5               g081(.a(\a[17] ), .o1(new_n177));
  nanb03aa1n02x5               g082(.a(new_n97), .b(new_n145), .c(new_n127), .out0(new_n178));
  xnrc02aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .out0(new_n179));
  nona22aa1n06x5               g084(.a(new_n165), .b(new_n179), .c(new_n173), .out0(new_n180));
  nor042aa1n03x5               g085(.a(new_n180), .b(new_n178), .o1(new_n181));
  norp02aa1n02x5               g086(.a(new_n173), .b(new_n179), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\a[16] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[15] ), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(new_n183), .b(new_n184), .c(new_n171), .o1(new_n185));
  aobi12aa1n06x5               g090(.a(new_n185), .b(new_n182), .c(new_n167), .out0(new_n186));
  oai012aa1n12x5               g091(.a(new_n186), .b(new_n180), .c(new_n147), .o1(new_n187));
  aoi012aa1n12x5               g092(.a(new_n187), .b(new_n158), .c(new_n181), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(new_n177), .out0(\s[17] ));
  oaoi03aa1n02x5               g094(.a(\a[17] ), .b(\b[16] ), .c(new_n188), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  norp02aa1n02x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  nand42aa1n03x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  norb02aa1n02x5               g100(.a(new_n192), .b(new_n195), .out0(new_n196));
  norp02aa1n02x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  tech160nm_fioai012aa1n04x5   g102(.a(new_n194), .b(new_n193), .c(new_n197), .o1(new_n198));
  oaib12aa1n06x5               g103(.a(new_n198), .b(new_n188), .c(new_n196), .out0(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand42aa1n03x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  nor002aa1n02x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nanp02aa1n04x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n03x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  aoai13aa1n03x5               g112(.a(new_n207), .b(new_n202), .c(new_n199), .d(new_n204), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(new_n199), .b(new_n204), .o1(new_n209));
  nona22aa1n02x4               g114(.a(new_n209), .b(new_n207), .c(new_n202), .out0(new_n210));
  nanp02aa1n02x5               g115(.a(new_n210), .b(new_n208), .o1(\s[20] ));
  nona23aa1n06x5               g116(.a(new_n204), .b(new_n192), .c(new_n207), .d(new_n195), .out0(new_n212));
  nona23aa1n02x4               g117(.a(new_n206), .b(new_n203), .c(new_n202), .d(new_n205), .out0(new_n213));
  tech160nm_fiaoi012aa1n05x5   g118(.a(new_n205), .b(new_n202), .c(new_n206), .o1(new_n214));
  tech160nm_fioai012aa1n05x5   g119(.a(new_n214), .b(new_n213), .c(new_n198), .o1(new_n215));
  oabi12aa1n06x5               g120(.a(new_n215), .b(new_n188), .c(new_n212), .out0(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  xnrc02aa1n02x5               g125(.a(\b[21] ), .b(\a[22] ), .out0(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n218), .c(new_n216), .d(new_n220), .o1(new_n222));
  aoi112aa1n03x4               g127(.a(new_n218), .b(new_n221), .c(new_n216), .d(new_n220), .o1(new_n223));
  nanb02aa1n03x5               g128(.a(new_n223), .b(new_n222), .out0(\s[22] ));
  nor042aa1n02x5               g129(.a(new_n221), .b(new_n219), .o1(new_n225));
  nona23aa1n02x4               g130(.a(new_n225), .b(new_n192), .c(new_n213), .d(new_n195), .out0(new_n226));
  inv000aa1n02x5               g131(.a(new_n198), .o1(new_n227));
  nano23aa1n02x4               g132(.a(new_n202), .b(new_n205), .c(new_n206), .d(new_n203), .out0(new_n228));
  inv000aa1n02x5               g133(.a(new_n214), .o1(new_n229));
  aoai13aa1n06x5               g134(.a(new_n225), .b(new_n229), .c(new_n228), .d(new_n227), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\a[22] ), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\b[21] ), .o1(new_n232));
  oao003aa1n06x5               g137(.a(new_n231), .b(new_n232), .c(new_n218), .carry(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(new_n230), .b(new_n234), .o1(new_n235));
  oabi12aa1n06x5               g140(.a(new_n235), .b(new_n188), .c(new_n226), .out0(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[22] ), .b(\a[23] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  xnrc02aa1n02x5               g145(.a(\b[23] ), .b(\a[24] ), .out0(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n238), .c(new_n236), .d(new_n240), .o1(new_n242));
  aoi112aa1n03x4               g147(.a(new_n238), .b(new_n241), .c(new_n236), .d(new_n240), .o1(new_n243));
  nanb02aa1n03x5               g148(.a(new_n243), .b(new_n242), .out0(\s[24] ));
  inv000aa1n02x5               g149(.a(new_n225), .o1(new_n245));
  norp02aa1n06x5               g150(.a(new_n212), .b(new_n245), .o1(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n187), .c(new_n158), .d(new_n181), .o1(new_n247));
  nor002aa1n03x5               g152(.a(new_n241), .b(new_n239), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  oai022aa1n02x5               g154(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n250));
  aob012aa1n02x5               g155(.a(new_n250), .b(\b[23] ), .c(\a[24] ), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n249), .c(new_n230), .d(new_n234), .o1(new_n252));
  oabi12aa1n06x5               g157(.a(new_n252), .b(new_n247), .c(new_n249), .out0(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g159(.a(\b[24] ), .b(\a[25] ), .o1(new_n255));
  xorc02aa1n06x5               g160(.a(\a[25] ), .b(\b[24] ), .out0(new_n256));
  xnrc02aa1n02x5               g161(.a(\b[25] ), .b(\a[26] ), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n255), .c(new_n253), .d(new_n256), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(new_n253), .b(new_n256), .o1(new_n259));
  nona22aa1n02x4               g164(.a(new_n259), .b(new_n257), .c(new_n255), .out0(new_n260));
  nanp02aa1n02x5               g165(.a(new_n260), .b(new_n258), .o1(\s[26] ));
  norb02aa1n02x5               g166(.a(new_n256), .b(new_n257), .out0(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  nona22aa1n02x4               g168(.a(new_n246), .b(new_n263), .c(new_n249), .out0(new_n264));
  nanp02aa1n02x5               g169(.a(new_n252), .b(new_n262), .o1(new_n265));
  oai022aa1n02x5               g170(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n266));
  aob012aa1n02x5               g171(.a(new_n266), .b(\b[25] ), .c(\a[26] ), .out0(new_n267));
  oai112aa1n06x5               g172(.a(new_n265), .b(new_n267), .c(new_n188), .d(new_n264), .o1(new_n268));
  xorb03aa1n03x5               g173(.a(new_n268), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n06x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[27] ), .b(\b[26] ), .out0(new_n271));
  xnrc02aa1n02x5               g176(.a(\b[27] ), .b(\a[28] ), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n270), .c(new_n268), .d(new_n271), .o1(new_n273));
  aoi012aa1n02x5               g178(.a(new_n126), .b(new_n118), .c(new_n108), .o1(new_n274));
  nano32aa1n02x4               g179(.a(new_n173), .b(new_n172), .c(new_n161), .d(new_n148), .out0(new_n275));
  nanp02aa1n02x5               g180(.a(new_n275), .b(new_n143), .o1(new_n276));
  oai013aa1n02x4               g181(.a(new_n185), .b(new_n168), .c(new_n179), .d(new_n173), .o1(new_n277));
  aoi012aa1n02x7               g182(.a(new_n277), .b(new_n159), .c(new_n275), .o1(new_n278));
  oaoi13aa1n04x5               g183(.a(new_n264), .b(new_n278), .c(new_n274), .d(new_n276), .o1(new_n279));
  aoai13aa1n04x5               g184(.a(new_n248), .b(new_n233), .c(new_n215), .d(new_n225), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n267), .b(new_n263), .c(new_n280), .d(new_n251), .o1(new_n281));
  oaih12aa1n02x5               g186(.a(new_n271), .b(new_n281), .c(new_n279), .o1(new_n282));
  nona22aa1n02x4               g187(.a(new_n282), .b(new_n272), .c(new_n270), .out0(new_n283));
  nanp02aa1n03x5               g188(.a(new_n273), .b(new_n283), .o1(\s[28] ));
  norb02aa1n02x5               g189(.a(new_n271), .b(new_n272), .out0(new_n285));
  oaih12aa1n02x5               g190(.a(new_n285), .b(new_n281), .c(new_n279), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\a[28] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[27] ), .o1(new_n288));
  oaoi03aa1n12x5               g193(.a(new_n287), .b(new_n288), .c(new_n270), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[29] ), .b(\b[28] ), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  tech160nm_fiaoi012aa1n03p5x5 g196(.a(new_n291), .b(new_n286), .c(new_n289), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n289), .o1(new_n293));
  aoi112aa1n03x4               g198(.a(new_n290), .b(new_n293), .c(new_n268), .d(new_n285), .o1(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g201(.a(new_n272), .b(new_n271), .c(new_n290), .out0(new_n297));
  oaih12aa1n02x5               g202(.a(new_n297), .b(new_n281), .c(new_n279), .o1(new_n298));
  tech160nm_fioaoi03aa1n03p5x5 g203(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .o1(new_n299));
  inv040aa1n03x5               g204(.a(new_n299), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  tech160nm_fiaoi012aa1n03p5x5 g207(.a(new_n302), .b(new_n298), .c(new_n300), .o1(new_n303));
  aoi112aa1n03x4               g208(.a(new_n301), .b(new_n299), .c(new_n268), .d(new_n297), .o1(new_n304));
  nor042aa1n03x5               g209(.a(new_n303), .b(new_n304), .o1(\s[30] ));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  nano23aa1n02x4               g211(.a(new_n302), .b(new_n272), .c(new_n271), .d(new_n290), .out0(new_n307));
  oaih12aa1n02x5               g212(.a(new_n307), .b(new_n281), .c(new_n279), .o1(new_n308));
  tech160nm_fioaoi03aa1n03p5x5 g213(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .o1(new_n309));
  inv000aa1n02x5               g214(.a(new_n309), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n306), .b(new_n308), .c(new_n310), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n306), .o1(new_n312));
  aoi112aa1n03x4               g217(.a(new_n312), .b(new_n309), .c(new_n268), .d(new_n307), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[31] ));
  xorb03aa1n02x5               g219(.a(new_n103), .b(\b[2] ), .c(new_n104), .out0(\s[3] ));
  nanb02aa1n02x5               g220(.a(\b[3] ), .b(new_n105), .out0(new_n316));
  aoi022aa1n02x5               g221(.a(new_n316), .b(new_n116), .c(new_n106), .d(new_n104), .o1(new_n317));
  nanp02aa1n02x5               g222(.a(new_n108), .b(new_n116), .o1(new_n318));
  aboi22aa1n03x5               g223(.a(new_n318), .b(new_n316), .c(new_n152), .d(new_n317), .out0(\s[4] ));
  xobna2aa1n03x5               g224(.a(new_n114), .b(new_n108), .c(new_n116), .out0(\s[5] ));
  aoi013aa1n02x4               g225(.a(new_n123), .b(new_n108), .c(new_n114), .d(new_n116), .o1(new_n321));
  xnbna2aa1n03x5               g226(.a(new_n321), .b(new_n109), .c(new_n112), .out0(\s[6] ));
  oaoi03aa1n02x5               g227(.a(\a[6] ), .b(\b[5] ), .c(new_n321), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  norp02aa1n02x5               g229(.a(\b[6] ), .b(\a[7] ), .o1(new_n325));
  aoi012aa1n02x5               g230(.a(new_n325), .b(new_n323), .c(new_n121), .o1(new_n326));
  xnrb03aa1n02x5               g231(.a(new_n326), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n158), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


