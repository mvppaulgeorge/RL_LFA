// Benchmark "adder" written by ABC on Thu Jul 18 09:57:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n331, new_n333, new_n334, new_n335, new_n336, new_n339, new_n341,
    new_n343;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d30x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[8] ), .o1(new_n98));
  oa0022aa1n03x5               g003(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n99));
  inv020aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  xnrc02aa1n12x5               g005(.a(\b[2] ), .b(\a[3] ), .out0(new_n101));
  nand42aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand02aa1d16x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor042aa1n09x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oai012aa1n12x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  oab012aa1n09x5               g010(.a(new_n100), .b(new_n101), .c(new_n105), .out0(new_n106));
  nanp02aa1n09x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nor042aa1n06x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand42aa1n10x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  nano22aa1n12x5               g014(.a(new_n108), .b(new_n107), .c(new_n109), .out0(new_n110));
  tech160nm_fixnrc02aa1n02p5x5 g015(.a(\b[7] ), .b(\a[8] ), .out0(new_n111));
  nor002aa1d32x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nanp02aa1n24x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n12x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nanb03aa1n09x5               g021(.a(new_n111), .b(new_n116), .c(new_n110), .out0(new_n117));
  inv000aa1n02x5               g022(.a(new_n108), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[8] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[7] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  tech160nm_fioai012aa1n03p5x5 g026(.a(new_n113), .b(new_n114), .c(new_n112), .o1(new_n122));
  aob012aa1n02x5               g027(.a(new_n107), .b(\b[7] ), .c(\a[8] ), .out0(new_n123));
  aoai13aa1n06x5               g028(.a(new_n121), .b(new_n123), .c(new_n122), .d(new_n118), .o1(new_n124));
  oabi12aa1n18x5               g029(.a(new_n124), .b(new_n117), .c(new_n106), .out0(new_n125));
  oaoi03aa1n09x5               g030(.a(new_n97), .b(new_n98), .c(new_n125), .o1(new_n126));
  nor042aa1d18x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1d28x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n15x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnrc02aa1n02x5               g034(.a(new_n126), .b(new_n129), .out0(\s[10] ));
  nanp02aa1n06x5               g035(.a(new_n126), .b(new_n129), .o1(new_n131));
  inv040aa1d32x5               g036(.a(\a[11] ), .o1(new_n132));
  inv040aa1d32x5               g037(.a(\b[10] ), .o1(new_n133));
  nand02aa1d28x5               g038(.a(new_n133), .b(new_n132), .o1(new_n134));
  nand22aa1n12x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand22aa1n09x5               g040(.a(new_n134), .b(new_n135), .o1(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n131), .c(new_n128), .out0(\s[11] ));
  xorc02aa1n12x5               g042(.a(\a[11] ), .b(\b[10] ), .out0(new_n138));
  nand03aa1n02x5               g043(.a(new_n131), .b(new_n128), .c(new_n138), .o1(new_n139));
  inv000aa1d42x5               g044(.a(\b[11] ), .o1(new_n140));
  nanb02aa1d36x5               g045(.a(\a[12] ), .b(new_n140), .out0(new_n141));
  nand42aa1d28x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n04x5               g047(.a(new_n141), .b(new_n142), .o1(new_n143));
  tech160nm_fiaoi012aa1n02p5x5 g048(.a(new_n143), .b(new_n139), .c(new_n134), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n134), .o1(new_n145));
  nor002aa1n03x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  norb02aa1n06x5               g051(.a(new_n142), .b(new_n146), .out0(new_n147));
  aoi113aa1n03x5               g052(.a(new_n147), .b(new_n145), .c(new_n131), .d(new_n138), .e(new_n128), .o1(new_n148));
  nor002aa1n02x5               g053(.a(new_n144), .b(new_n148), .o1(\s[12] ));
  tech160nm_fioai012aa1n03p5x5 g054(.a(new_n99), .b(new_n101), .c(new_n105), .o1(new_n150));
  nona23aa1n03x5               g055(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n151));
  nor042aa1n02x5               g056(.a(new_n151), .b(new_n111), .o1(new_n152));
  aoi013aa1n06x4               g057(.a(new_n124), .b(new_n152), .c(new_n150), .d(new_n110), .o1(new_n153));
  tech160nm_fixnrc02aa1n04x5   g058(.a(\b[8] ), .b(\a[9] ), .out0(new_n154));
  nona23aa1n02x4               g059(.a(new_n147), .b(new_n129), .c(new_n154), .d(new_n136), .out0(new_n155));
  nona22aa1n03x5               g060(.a(new_n142), .b(\b[10] ), .c(\a[11] ), .out0(new_n156));
  aoai13aa1n06x5               g061(.a(new_n128), .b(new_n127), .c(new_n97), .d(new_n98), .o1(new_n157));
  nor003aa1n03x5               g062(.a(new_n157), .b(new_n143), .c(new_n136), .o1(new_n158));
  nano22aa1n03x7               g063(.a(new_n158), .b(new_n141), .c(new_n156), .out0(new_n159));
  tech160nm_fioai012aa1n05x5   g064(.a(new_n159), .b(new_n153), .c(new_n155), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  orn002aa1n02x5               g066(.a(\a[13] ), .b(\b[12] ), .o(new_n162));
  nano23aa1n03x7               g067(.a(new_n154), .b(new_n136), .c(new_n147), .d(new_n129), .out0(new_n163));
  nanb03aa1n06x5               g068(.a(new_n157), .b(new_n138), .c(new_n147), .out0(new_n164));
  nand23aa1n06x5               g069(.a(new_n164), .b(new_n141), .c(new_n156), .o1(new_n165));
  xorc02aa1n12x5               g070(.a(\a[13] ), .b(\b[12] ), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n165), .c(new_n125), .d(new_n163), .o1(new_n167));
  xnrc02aa1n12x5               g072(.a(\b[13] ), .b(\a[14] ), .out0(new_n168));
  xobna2aa1n03x5               g073(.a(new_n168), .b(new_n167), .c(new_n162), .out0(\s[14] ));
  nand22aa1n03x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  xnrc02aa1n12x5               g075(.a(\b[14] ), .b(\a[15] ), .out0(new_n171));
  oai022aa1d18x5               g076(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n172));
  nanb02aa1n03x5               g077(.a(new_n172), .b(new_n167), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n171), .b(new_n173), .c(new_n170), .out0(\s[15] ));
  nor002aa1n16x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  and002aa1n06x5               g080(.a(\b[14] ), .b(\a[15] ), .o(new_n176));
  aoi112aa1n02x5               g081(.a(new_n176), .b(new_n175), .c(\a[14] ), .d(\b[13] ), .o1(new_n177));
  xorc02aa1n12x5               g082(.a(\a[16] ), .b(\b[15] ), .out0(new_n178));
  aoi112aa1n03x4               g083(.a(new_n178), .b(new_n175), .c(new_n173), .d(new_n177), .o1(new_n179));
  inv000aa1d42x5               g084(.a(new_n175), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n177), .b(new_n172), .c(new_n160), .d(new_n166), .o1(new_n181));
  aobi12aa1n02x7               g086(.a(new_n178), .b(new_n181), .c(new_n180), .out0(new_n182));
  norp02aa1n03x5               g087(.a(new_n182), .b(new_n179), .o1(\s[16] ));
  nona23aa1n03x5               g088(.a(new_n166), .b(new_n178), .c(new_n171), .d(new_n168), .out0(new_n184));
  nor042aa1n03x5               g089(.a(new_n184), .b(new_n155), .o1(new_n185));
  nanp02aa1n06x5               g090(.a(new_n125), .b(new_n185), .o1(new_n186));
  nanp02aa1n02x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nano23aa1n09x5               g092(.a(new_n171), .b(new_n168), .c(new_n178), .d(new_n166), .out0(new_n188));
  aoi012aa1n06x5               g093(.a(new_n175), .b(new_n172), .c(new_n170), .o1(new_n189));
  oai022aa1n12x5               g094(.a(new_n189), .b(new_n176), .c(\b[15] ), .d(\a[16] ), .o1(new_n190));
  aoi022aa1d18x5               g095(.a(new_n165), .b(new_n188), .c(new_n187), .d(new_n190), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n192), .b(new_n186), .c(new_n191), .out0(\s[17] ));
  inv040aa1d32x5               g098(.a(\a[18] ), .o1(new_n194));
  inv040aa1d28x5               g099(.a(\a[17] ), .o1(new_n195));
  inv000aa1d42x5               g100(.a(\b[16] ), .o1(new_n196));
  nand02aa1n02x5               g101(.a(new_n188), .b(new_n163), .o1(new_n197));
  oai012aa1n12x5               g102(.a(new_n191), .b(new_n197), .c(new_n153), .o1(new_n198));
  oaoi03aa1n03x5               g103(.a(new_n195), .b(new_n196), .c(new_n198), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[17] ), .c(new_n194), .out0(\s[18] ));
  nand42aa1d28x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand42aa1d28x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nor002aa1d32x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  nand42aa1n03x5               g109(.a(new_n190), .b(new_n187), .o1(new_n205));
  tech160nm_fioai012aa1n05x5   g110(.a(new_n205), .b(new_n159), .c(new_n184), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n192), .b(new_n206), .c(new_n125), .d(new_n185), .o1(new_n207));
  oai022aa1d24x5               g112(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n208));
  nanb02aa1n03x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  aoi022aa1n03x5               g114(.a(new_n209), .b(new_n201), .c(new_n202), .d(new_n204), .o1(new_n210));
  nano22aa1d15x5               g115(.a(new_n203), .b(new_n201), .c(new_n202), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n208), .c(new_n198), .d(new_n192), .o1(new_n212));
  norb02aa1n02x7               g117(.a(new_n212), .b(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nand42aa1d28x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  norb02aa1n06x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  aobi12aa1n03x5               g122(.a(new_n217), .b(new_n212), .c(new_n204), .out0(new_n218));
  aoi112aa1n03x4               g123(.a(new_n217), .b(new_n203), .c(new_n209), .d(new_n211), .o1(new_n219));
  norp02aa1n03x5               g124(.a(new_n218), .b(new_n219), .o1(\s[20] ));
  xroi22aa1d06x4               g125(.a(new_n195), .b(\b[16] ), .c(new_n194), .d(\b[17] ), .out0(new_n221));
  nanb03aa1n02x5               g126(.a(new_n215), .b(new_n216), .c(new_n202), .out0(new_n222));
  nona22aa1n09x5               g127(.a(new_n221), .b(new_n222), .c(new_n203), .out0(new_n223));
  nanb03aa1d18x5               g128(.a(new_n203), .b(new_n201), .c(new_n202), .out0(new_n224));
  oai012aa1n12x5               g129(.a(new_n216), .b(new_n215), .c(new_n203), .o1(new_n225));
  inv020aa1n10x5               g130(.a(\b[19] ), .o1(new_n226));
  nanb02aa1n12x5               g131(.a(\a[20] ), .b(new_n226), .out0(new_n227));
  nand23aa1n06x5               g132(.a(new_n208), .b(new_n227), .c(new_n216), .o1(new_n228));
  oai012aa1d24x5               g133(.a(new_n225), .b(new_n228), .c(new_n224), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n04x5               g135(.a(new_n230), .b(new_n223), .c(new_n186), .d(new_n191), .o1(new_n231));
  xorb03aa1n02x5               g136(.a(new_n231), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  xorc02aa1n12x5               g138(.a(\a[21] ), .b(\b[20] ), .out0(new_n234));
  xorc02aa1n12x5               g139(.a(\a[22] ), .b(\b[21] ), .out0(new_n235));
  aoi112aa1n03x4               g140(.a(new_n233), .b(new_n235), .c(new_n231), .d(new_n234), .o1(new_n236));
  inv040aa1n08x5               g141(.a(new_n233), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n223), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n234), .b(new_n229), .c(new_n198), .d(new_n238), .o1(new_n239));
  aobi12aa1n02x7               g144(.a(new_n235), .b(new_n239), .c(new_n237), .out0(new_n240));
  nor002aa1n02x5               g145(.a(new_n240), .b(new_n236), .o1(\s[22] ));
  inv030aa1d32x5               g146(.a(\a[21] ), .o1(new_n242));
  inv030aa1d32x5               g147(.a(\a[22] ), .o1(new_n243));
  xroi22aa1d06x4               g148(.a(new_n242), .b(\b[20] ), .c(new_n243), .d(\b[21] ), .out0(new_n244));
  nona23aa1n06x5               g149(.a(new_n244), .b(new_n221), .c(new_n203), .d(new_n222), .out0(new_n245));
  nanp03aa1d12x5               g150(.a(new_n211), .b(new_n208), .c(new_n217), .o1(new_n246));
  nand02aa1n03x5               g151(.a(new_n235), .b(new_n234), .o1(new_n247));
  oaoi03aa1n09x5               g152(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n247), .c(new_n246), .d(new_n225), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n04x5               g156(.a(new_n251), .b(new_n245), .c(new_n186), .d(new_n191), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n09x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  nanp02aa1n04x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  aoi112aa1n03x4               g161(.a(new_n254), .b(new_n256), .c(new_n252), .d(new_n255), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n254), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n245), .o1(new_n259));
  norb02aa1n02x7               g164(.a(new_n255), .b(new_n254), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n250), .c(new_n198), .d(new_n259), .o1(new_n261));
  aobi12aa1n02x7               g166(.a(new_n256), .b(new_n261), .c(new_n258), .out0(new_n262));
  nor002aa1n02x5               g167(.a(new_n262), .b(new_n257), .o1(\s[24] ));
  nano32aa1n03x7               g168(.a(new_n223), .b(new_n256), .c(new_n244), .d(new_n260), .out0(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n206), .c(new_n125), .d(new_n185), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n255), .b(new_n248), .c(new_n229), .d(new_n244), .o1(new_n266));
  inv000aa1d42x5               g171(.a(\a[24] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(\b[23] ), .o1(new_n268));
  aoi012aa1d18x5               g173(.a(new_n254), .b(new_n267), .c(new_n268), .o1(new_n269));
  aoi022aa1n03x5               g174(.a(new_n266), .b(new_n269), .c(\b[23] ), .d(\a[24] ), .o1(new_n270));
  xnrc02aa1n12x5               g175(.a(\b[24] ), .b(\a[25] ), .out0(new_n271));
  aoib12aa1n06x5               g176(.a(new_n271), .b(new_n265), .c(new_n270), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n271), .o1(new_n273));
  aoi112aa1n02x5               g178(.a(new_n273), .b(new_n270), .c(new_n198), .d(new_n264), .o1(new_n274));
  nor002aa1n02x5               g179(.a(new_n272), .b(new_n274), .o1(\s[25] ));
  orn002aa1n02x5               g180(.a(\a[25] ), .b(\b[24] ), .o(new_n276));
  aoai13aa1n03x5               g181(.a(new_n273), .b(new_n270), .c(new_n198), .d(new_n264), .o1(new_n277));
  xnrc02aa1n12x5               g182(.a(\b[25] ), .b(\a[26] ), .out0(new_n278));
  tech160nm_fiaoi012aa1n02p5x5 g183(.a(new_n278), .b(new_n277), .c(new_n276), .o1(new_n279));
  nano22aa1n03x7               g184(.a(new_n272), .b(new_n276), .c(new_n278), .out0(new_n280));
  norp02aa1n03x5               g185(.a(new_n279), .b(new_n280), .o1(\s[26] ));
  and002aa1n02x5               g186(.a(\b[23] ), .b(\a[24] ), .o(new_n282));
  nor043aa1d12x5               g187(.a(new_n278), .b(new_n271), .c(new_n282), .o1(new_n283));
  nano32aa1n03x7               g188(.a(new_n245), .b(new_n283), .c(new_n260), .d(new_n256), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n206), .c(new_n125), .d(new_n185), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n269), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n283), .b(new_n286), .c(new_n250), .d(new_n255), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[26] ), .b(\b[25] ), .c(new_n276), .carry(new_n288));
  xorc02aa1n12x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  inv000aa1d42x5               g194(.a(new_n289), .o1(new_n290));
  aoi013aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n287), .d(new_n288), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n283), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n288), .b(new_n292), .c(new_n266), .d(new_n269), .o1(new_n293));
  aoi112aa1n02x5               g198(.a(new_n293), .b(new_n289), .c(new_n198), .d(new_n284), .o1(new_n294));
  nor002aa1n02x5               g199(.a(new_n291), .b(new_n294), .o1(\s[27] ));
  nor042aa1n03x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  inv040aa1n03x5               g201(.a(new_n296), .o1(new_n297));
  xnrc02aa1n12x5               g202(.a(\b[27] ), .b(\a[28] ), .out0(new_n298));
  nano22aa1n03x5               g203(.a(new_n291), .b(new_n297), .c(new_n298), .out0(new_n299));
  aoai13aa1n02x5               g204(.a(new_n289), .b(new_n293), .c(new_n198), .d(new_n284), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  norp02aa1n03x5               g206(.a(new_n301), .b(new_n299), .o1(\s[28] ));
  norb02aa1n02x5               g207(.a(new_n289), .b(new_n298), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n293), .c(new_n198), .d(new_n284), .o1(new_n304));
  oao003aa1n03x5               g209(.a(\a[28] ), .b(\b[27] ), .c(new_n297), .carry(new_n305));
  xnrc02aa1n12x5               g210(.a(\b[28] ), .b(\a[29] ), .out0(new_n306));
  tech160nm_fiaoi012aa1n02p5x5 g211(.a(new_n306), .b(new_n304), .c(new_n305), .o1(new_n307));
  inv000aa1n02x5               g212(.a(new_n303), .o1(new_n308));
  aoi013aa1n02x5               g213(.a(new_n308), .b(new_n285), .c(new_n287), .d(new_n288), .o1(new_n309));
  nano22aa1n03x5               g214(.a(new_n309), .b(new_n305), .c(new_n306), .out0(new_n310));
  norp02aa1n03x5               g215(.a(new_n307), .b(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g216(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g217(.a(new_n289), .b(new_n306), .c(new_n298), .out0(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n293), .c(new_n198), .d(new_n284), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[29] ), .b(\a[30] ), .out0(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n314), .c(new_n315), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n313), .o1(new_n318));
  aoi013aa1n03x5               g223(.a(new_n318), .b(new_n285), .c(new_n287), .d(new_n288), .o1(new_n319));
  nano22aa1n02x4               g224(.a(new_n319), .b(new_n315), .c(new_n316), .out0(new_n320));
  norp02aa1n03x5               g225(.a(new_n317), .b(new_n320), .o1(\s[30] ));
  norb02aa1n02x5               g226(.a(new_n313), .b(new_n316), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n293), .c(new_n198), .d(new_n284), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n324));
  xnrc02aa1n02x5               g229(.a(\b[30] ), .b(\a[31] ), .out0(new_n325));
  tech160nm_fiaoi012aa1n02p5x5 g230(.a(new_n325), .b(new_n323), .c(new_n324), .o1(new_n326));
  inv000aa1n02x5               g231(.a(new_n322), .o1(new_n327));
  aoi013aa1n02x5               g232(.a(new_n327), .b(new_n285), .c(new_n287), .d(new_n288), .o1(new_n328));
  nano22aa1n02x4               g233(.a(new_n328), .b(new_n324), .c(new_n325), .out0(new_n329));
  norp02aa1n03x5               g234(.a(new_n326), .b(new_n329), .o1(\s[31] ));
  inv000aa1d42x5               g235(.a(\a[3] ), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n105), .b(\b[2] ), .c(new_n331), .out0(\s[3] ));
  norb02aa1n02x5               g237(.a(new_n109), .b(new_n106), .out0(new_n333));
  xorc02aa1n02x5               g238(.a(\a[4] ), .b(\b[3] ), .out0(new_n334));
  oabi12aa1n02x5               g239(.a(new_n334), .b(new_n101), .c(new_n105), .out0(new_n335));
  aoib12aa1n02x5               g240(.a(new_n335), .b(new_n331), .c(\b[2] ), .out0(new_n336));
  oaoi13aa1n02x5               g241(.a(new_n336), .b(new_n333), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g242(.a(new_n333), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi013aa1n02x4               g243(.a(new_n114), .b(new_n150), .c(new_n109), .d(new_n115), .o1(new_n339));
  xnrb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n03x5               g245(.a(\a[6] ), .b(\b[5] ), .c(new_n339), .o1(new_n341));
  xorb03aa1n02x5               g246(.a(new_n341), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g247(.a(new_n108), .b(new_n341), .c(new_n107), .o1(new_n343));
  xorb03aa1n02x5               g248(.a(new_n343), .b(\b[7] ), .c(new_n119), .out0(\s[8] ));
  xorb03aa1n02x5               g249(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


