// Benchmark "adder" written by ABC on Thu Jul 18 05:14:13 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n320, new_n321, new_n322, new_n324,
    new_n325, new_n326, new_n328, new_n329, new_n330, new_n332, new_n334,
    new_n335, new_n336, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n04x5   g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\a[9] ), .b(new_n98), .out0(new_n99));
  and002aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o(new_n100));
  oaoi03aa1n09x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  xorc02aa1n12x5               g006(.a(\a[3] ), .b(\b[2] ), .out0(new_n102));
  oai022aa1n02x5               g007(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  aoi012aa1n12x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .o1(new_n104));
  nor042aa1n06x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  and002aa1n12x5               g010(.a(\b[6] ), .b(\a[7] ), .o(new_n106));
  aoi112aa1n03x5               g011(.a(new_n106), .b(new_n105), .c(\a[8] ), .d(\b[7] ), .o1(new_n107));
  inv040aa1d32x5               g012(.a(\a[5] ), .o1(new_n108));
  inv040aa1d28x5               g013(.a(\b[4] ), .o1(new_n109));
  aoi022aa1n02x5               g014(.a(new_n109), .b(new_n108), .c(\a[4] ), .d(\b[3] ), .o1(new_n110));
  and002aa1n03x5               g015(.a(\b[4] ), .b(\a[5] ), .o(new_n111));
  and002aa1n02x5               g016(.a(\b[5] ), .b(\a[6] ), .o(new_n112));
  oaih22aa1n04x5               g017(.a(\a[6] ), .b(\b[5] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n113));
  nor043aa1n02x5               g018(.a(new_n113), .b(new_n112), .c(new_n111), .o1(new_n114));
  nand23aa1n03x5               g019(.a(new_n114), .b(new_n107), .c(new_n110), .o1(new_n115));
  tech160nm_fixorc02aa1n04x5   g020(.a(\a[8] ), .b(\b[7] ), .out0(new_n116));
  nor042aa1n02x5               g021(.a(new_n106), .b(new_n105), .o1(new_n117));
  nand02aa1d04x5               g022(.a(new_n109), .b(new_n108), .o1(new_n118));
  oaoi03aa1n02x5               g023(.a(\a[6] ), .b(\b[5] ), .c(new_n118), .o1(new_n119));
  inv000aa1n02x5               g024(.a(new_n105), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  aoi013aa1n06x4               g026(.a(new_n121), .b(new_n119), .c(new_n116), .d(new_n117), .o1(new_n122));
  oai012aa1n18x5               g027(.a(new_n122), .b(new_n104), .c(new_n115), .o1(new_n123));
  oaib12aa1n06x5               g028(.a(new_n123), .b(new_n98), .c(\a[9] ), .out0(new_n124));
  xnbna2aa1n03x5               g029(.a(new_n97), .b(new_n124), .c(new_n99), .out0(\s[10] ));
  nanp02aa1n02x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nor002aa1d32x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  oaih22aa1d12x5               g033(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n129));
  nanb02aa1n02x5               g034(.a(new_n129), .b(new_n124), .out0(new_n130));
  aob012aa1n02x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n127), .o1(new_n132));
  aoi022aa1n06x5               g037(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n133));
  nanp03aa1n03x5               g038(.a(new_n130), .b(new_n132), .c(new_n133), .o1(new_n134));
  aobi12aa1n02x5               g039(.a(new_n134), .b(new_n131), .c(new_n128), .out0(\s[11] ));
  nor002aa1n02x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand42aa1n08x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x7               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  nor002aa1n02x5               g043(.a(new_n136), .b(new_n127), .o1(new_n139));
  nanp03aa1n02x5               g044(.a(new_n134), .b(new_n137), .c(new_n139), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n140), .b(new_n138), .c(new_n132), .d(new_n134), .o1(\s[12] ));
  xnrc02aa1n02x5               g046(.a(\b[8] ), .b(\a[9] ), .out0(new_n142));
  nona23aa1n09x5               g047(.a(new_n138), .b(new_n97), .c(new_n142), .d(new_n128), .out0(new_n143));
  nanb02aa1n06x5               g048(.a(new_n143), .b(new_n123), .out0(new_n144));
  aob012aa1n03x5               g049(.a(new_n139), .b(new_n129), .c(new_n133), .out0(new_n145));
  nanp02aa1n02x5               g050(.a(new_n145), .b(new_n137), .o1(new_n146));
  xnrc02aa1n12x5               g051(.a(\b[12] ), .b(\a[13] ), .out0(new_n147));
  xobna2aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n146), .out0(\s[13] ));
  nor042aa1n09x5               g053(.a(\b[13] ), .b(\a[14] ), .o1(new_n149));
  nand02aa1d28x5               g054(.a(\b[13] ), .b(\a[14] ), .o1(new_n150));
  norb02aa1n12x5               g055(.a(new_n150), .b(new_n149), .out0(new_n151));
  inv000aa1d42x5               g056(.a(\a[13] ), .o1(new_n152));
  inv000aa1d42x5               g057(.a(\b[12] ), .o1(new_n153));
  nand22aa1n03x5               g058(.a(new_n144), .b(new_n146), .o1(new_n154));
  oaoi03aa1n02x5               g059(.a(new_n152), .b(new_n153), .c(new_n154), .o1(new_n155));
  oai022aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n150), .b(new_n156), .out0(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n147), .c(new_n144), .d(new_n146), .o1(new_n158));
  oai012aa1n02x5               g063(.a(new_n158), .b(new_n155), .c(new_n151), .o1(\s[14] ));
  norb02aa1d21x5               g064(.a(new_n151), .b(new_n147), .out0(new_n160));
  nanp02aa1n03x5               g065(.a(new_n154), .b(new_n160), .o1(new_n161));
  aoai13aa1n04x5               g066(.a(new_n150), .b(new_n149), .c(new_n152), .d(new_n153), .o1(new_n162));
  inv040aa1d32x5               g067(.a(\a[15] ), .o1(new_n163));
  inv000aa1d42x5               g068(.a(\b[14] ), .o1(new_n164));
  nand02aa1d28x5               g069(.a(new_n164), .b(new_n163), .o1(new_n165));
  tech160nm_finand02aa1n05x5   g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nanp02aa1n03x5               g071(.a(new_n165), .b(new_n166), .o1(new_n167));
  xobna2aa1n03x5               g072(.a(new_n167), .b(new_n161), .c(new_n162), .out0(\s[15] ));
  inv000aa1d42x5               g073(.a(new_n160), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n162), .b(new_n169), .c(new_n144), .d(new_n146), .o1(new_n170));
  inv000aa1d42x5               g075(.a(new_n165), .o1(new_n171));
  xnrc02aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .out0(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n171), .c(new_n170), .d(new_n166), .o1(new_n173));
  norp02aa1n02x5               g078(.a(new_n172), .b(new_n171), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n167), .c(new_n161), .d(new_n162), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n173), .b(new_n175), .o1(\s[16] ));
  nor002aa1n02x5               g081(.a(new_n172), .b(new_n167), .o1(new_n177));
  nano22aa1n12x5               g082(.a(new_n143), .b(new_n160), .c(new_n177), .out0(new_n178));
  nand02aa1d04x5               g083(.a(new_n123), .b(new_n178), .o1(new_n179));
  oai012aa1n02x5               g084(.a(new_n137), .b(\b[12] ), .c(\a[13] ), .o1(new_n180));
  oai022aa1n02x5               g085(.a(new_n152), .b(new_n153), .c(\b[13] ), .d(\a[14] ), .o1(new_n181));
  nano23aa1n06x5               g086(.a(new_n181), .b(new_n180), .c(new_n165), .d(new_n150), .out0(new_n182));
  norp02aa1n02x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  aob012aa1n02x5               g088(.a(new_n166), .b(\b[15] ), .c(\a[16] ), .out0(new_n184));
  nor002aa1n02x5               g089(.a(new_n184), .b(new_n183), .o1(new_n185));
  nanp03aa1n06x5               g090(.a(new_n182), .b(new_n145), .c(new_n185), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n183), .o1(new_n187));
  aoai13aa1n03x5               g092(.a(new_n187), .b(new_n184), .c(new_n162), .d(new_n165), .o1(new_n188));
  nanb02aa1n18x5               g093(.a(new_n188), .b(new_n186), .out0(new_n189));
  inv000aa1n03x5               g094(.a(new_n189), .o1(new_n190));
  xorc02aa1n06x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n179), .c(new_n190), .out0(\s[17] ));
  inv020aa1n10x5               g097(.a(\a[17] ), .o1(new_n193));
  nanb02aa1n12x5               g098(.a(\b[16] ), .b(new_n193), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n191), .b(new_n189), .c(new_n123), .d(new_n178), .o1(new_n195));
  xorc02aa1n12x5               g100(.a(\a[18] ), .b(\b[17] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n195), .c(new_n194), .out0(\s[18] ));
  and002aa1n02x5               g102(.a(new_n196), .b(new_n191), .o(new_n198));
  aoai13aa1n02x5               g103(.a(new_n198), .b(new_n189), .c(new_n123), .d(new_n178), .o1(new_n199));
  oaoi03aa1n12x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n194), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  nor042aa1n06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1n06x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n06x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n199), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g111(.a(new_n202), .o1(new_n207));
  nand02aa1d06x5               g112(.a(new_n179), .b(new_n190), .o1(new_n208));
  aoai13aa1n06x5               g113(.a(new_n204), .b(new_n200), .c(new_n208), .d(new_n198), .o1(new_n209));
  nor002aa1n03x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  tech160nm_finand02aa1n03p5x5 g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  norb02aa1n02x7               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  norb03aa1n02x5               g117(.a(new_n211), .b(new_n202), .c(new_n210), .out0(new_n213));
  nand42aa1n02x5               g118(.a(new_n209), .b(new_n213), .o1(new_n214));
  aoai13aa1n02x5               g119(.a(new_n214), .b(new_n212), .c(new_n209), .d(new_n207), .o1(\s[20] ));
  nano23aa1n06x5               g120(.a(new_n202), .b(new_n210), .c(new_n211), .d(new_n203), .out0(new_n216));
  nand23aa1n06x5               g121(.a(new_n216), .b(new_n191), .c(new_n196), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n189), .c(new_n123), .d(new_n178), .o1(new_n219));
  oaoi03aa1n09x5               g124(.a(\a[20] ), .b(\b[19] ), .c(new_n207), .o1(new_n220));
  aoi012aa1n02x5               g125(.a(new_n220), .b(new_n216), .c(new_n200), .o1(new_n221));
  xorc02aa1n03x5               g126(.a(\a[21] ), .b(\b[20] ), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n219), .c(new_n221), .out0(\s[21] ));
  norp02aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  aob012aa1n03x5               g130(.a(new_n222), .b(new_n219), .c(new_n221), .out0(new_n226));
  xorc02aa1n02x5               g131(.a(\a[22] ), .b(\b[21] ), .out0(new_n227));
  xnrc02aa1n02x5               g132(.a(\b[20] ), .b(\a[21] ), .out0(new_n228));
  nanp02aa1n02x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  oai022aa1n02x5               g134(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n229), .b(new_n230), .out0(new_n231));
  aoai13aa1n02x5               g136(.a(new_n231), .b(new_n228), .c(new_n219), .d(new_n221), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n227), .c(new_n226), .d(new_n225), .o1(\s[22] ));
  nanp02aa1n02x5               g138(.a(new_n227), .b(new_n222), .o1(new_n234));
  nano32aa1n02x4               g139(.a(new_n234), .b(new_n216), .c(new_n196), .d(new_n191), .out0(new_n235));
  norp02aa1n02x5               g140(.a(\b[17] ), .b(\a[18] ), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n237));
  oai112aa1n03x5               g142(.a(new_n204), .b(new_n212), .c(new_n237), .d(new_n236), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n220), .o1(new_n239));
  nanp02aa1n02x5               g144(.a(new_n230), .b(new_n229), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n238), .d(new_n239), .o1(new_n241));
  xorc02aa1n02x5               g146(.a(\a[23] ), .b(\b[22] ), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n241), .c(new_n208), .d(new_n235), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(new_n242), .b(new_n241), .c(new_n208), .d(new_n235), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n243), .b(new_n244), .out0(\s[23] ));
  nor042aa1n06x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  inv020aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[24] ), .b(\b[23] ), .out0(new_n248));
  nanp02aa1n02x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  oai022aa1n02x5               g154(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n250));
  norb02aa1n02x5               g155(.a(new_n249), .b(new_n250), .out0(new_n251));
  nanp02aa1n03x5               g156(.a(new_n243), .b(new_n251), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n248), .c(new_n247), .d(new_n243), .o1(\s[24] ));
  orn002aa1n02x5               g158(.a(\a[22] ), .b(\b[21] ), .o(new_n254));
  nano22aa1n02x5               g159(.a(new_n228), .b(new_n254), .c(new_n229), .out0(new_n255));
  nano32aa1n02x5               g160(.a(new_n217), .b(new_n248), .c(new_n255), .d(new_n242), .out0(new_n256));
  aoai13aa1n06x5               g161(.a(new_n255), .b(new_n220), .c(new_n216), .d(new_n200), .o1(new_n257));
  tech160nm_fixnrc02aa1n04x5   g162(.a(\b[22] ), .b(\a[23] ), .out0(new_n258));
  norb02aa1n09x5               g163(.a(new_n248), .b(new_n258), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  oaoi03aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .c(new_n247), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n262), .b(new_n260), .c(new_n257), .d(new_n240), .o1(new_n263));
  tech160nm_fixorc02aa1n03p5x5 g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n263), .c(new_n208), .d(new_n256), .o1(new_n265));
  aoi112aa1n02x5               g170(.a(new_n264), .b(new_n263), .c(new_n208), .d(new_n256), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n265), .b(new_n266), .out0(\s[25] ));
  norp02aa1n02x5               g172(.a(\b[24] ), .b(\a[25] ), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n268), .o1(new_n269));
  tech160nm_fixorc02aa1n02p5x5 g174(.a(\a[26] ), .b(\b[25] ), .out0(new_n270));
  nanp02aa1n02x5               g175(.a(\b[25] ), .b(\a[26] ), .o1(new_n271));
  oai022aa1n02x5               g176(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n272));
  norb02aa1n02x5               g177(.a(new_n271), .b(new_n272), .out0(new_n273));
  nanp02aa1n03x5               g178(.a(new_n265), .b(new_n273), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n270), .c(new_n269), .d(new_n265), .o1(\s[26] ));
  and002aa1n02x5               g180(.a(new_n270), .b(new_n264), .o(new_n276));
  nano32aa1n03x7               g181(.a(new_n217), .b(new_n276), .c(new_n255), .d(new_n259), .out0(new_n277));
  aoai13aa1n12x5               g182(.a(new_n277), .b(new_n189), .c(new_n123), .d(new_n178), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n276), .b(new_n261), .c(new_n241), .d(new_n259), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(new_n272), .b(new_n271), .o1(new_n280));
  nand03aa1n06x5               g185(.a(new_n278), .b(new_n279), .c(new_n280), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  aoi122aa1n02x5               g187(.a(new_n282), .b(new_n271), .c(new_n272), .d(new_n263), .e(new_n276), .o1(new_n283));
  aoi022aa1n02x5               g188(.a(new_n283), .b(new_n278), .c(new_n281), .d(new_n282), .o1(\s[27] ));
  nor042aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  xnrc02aa1n12x5               g190(.a(\b[27] ), .b(\a[28] ), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n281), .d(new_n282), .o1(new_n287));
  aoi022aa1n06x5               g192(.a(new_n263), .b(new_n276), .c(new_n271), .d(new_n272), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n282), .o1(new_n289));
  nor042aa1n03x5               g194(.a(new_n286), .b(new_n285), .o1(new_n290));
  aoai13aa1n02x5               g195(.a(new_n290), .b(new_n289), .c(new_n288), .d(new_n278), .o1(new_n291));
  nanp02aa1n03x5               g196(.a(new_n287), .b(new_n291), .o1(\s[28] ));
  norb02aa1n03x5               g197(.a(new_n282), .b(new_n286), .out0(new_n293));
  nanp02aa1n03x5               g198(.a(new_n281), .b(new_n293), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n293), .o1(new_n295));
  tech160nm_fiao0012aa1n05x5   g200(.a(new_n290), .b(\a[28] ), .c(\b[27] ), .o(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n295), .c(new_n288), .d(new_n278), .o1(new_n297));
  xorc02aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .out0(new_n298));
  norb02aa1n02x5               g203(.a(new_n296), .b(new_n298), .out0(new_n299));
  aoi022aa1n03x5               g204(.a(new_n297), .b(new_n298), .c(new_n294), .d(new_n299), .o1(\s[29] ));
  xnrb03aa1n02x5               g205(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g206(.a(new_n286), .b(new_n282), .c(new_n298), .out0(new_n302));
  nanp02aa1n03x5               g207(.a(new_n281), .b(new_n302), .o1(new_n303));
  inv000aa1n02x5               g208(.a(new_n302), .o1(new_n304));
  oaoi03aa1n12x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n305), .o1(new_n306));
  aoai13aa1n02x7               g211(.a(new_n306), .b(new_n304), .c(new_n288), .d(new_n278), .o1(new_n307));
  xorc02aa1n02x5               g212(.a(\a[30] ), .b(\b[29] ), .out0(new_n308));
  norp02aa1n02x5               g213(.a(new_n305), .b(new_n308), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n307), .b(new_n308), .c(new_n303), .d(new_n309), .o1(\s[30] ));
  nanp03aa1n02x5               g215(.a(new_n293), .b(new_n298), .c(new_n308), .o1(new_n311));
  nanb02aa1n03x5               g216(.a(new_n311), .b(new_n281), .out0(new_n312));
  inv000aa1d42x5               g217(.a(\a[30] ), .o1(new_n313));
  inv000aa1d42x5               g218(.a(\b[29] ), .o1(new_n314));
  oaoi03aa1n09x5               g219(.a(new_n313), .b(new_n314), .c(new_n305), .o1(new_n315));
  aoai13aa1n02x7               g220(.a(new_n315), .b(new_n311), .c(new_n288), .d(new_n278), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[31] ), .b(\b[30] ), .out0(new_n317));
  norb02aa1n03x4               g222(.a(new_n315), .b(new_n317), .out0(new_n318));
  aoi022aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n312), .d(new_n318), .o1(\s[31] ));
  orn002aa1n02x5               g224(.a(\a[2] ), .b(\b[1] ), .o(new_n320));
  nanp02aa1n02x5               g225(.a(\b[1] ), .b(\a[2] ), .o1(new_n321));
  nanb03aa1n02x5               g226(.a(new_n100), .b(new_n320), .c(new_n321), .out0(new_n322));
  xnbna2aa1n03x5               g227(.a(new_n102), .b(new_n322), .c(new_n320), .out0(\s[3] ));
  nanp02aa1n02x5               g228(.a(new_n101), .b(new_n102), .o1(new_n324));
  xorc02aa1n02x5               g229(.a(\a[4] ), .b(\b[3] ), .out0(new_n325));
  oab012aa1n02x4               g230(.a(new_n325), .b(\a[3] ), .c(\b[2] ), .out0(new_n326));
  aboi22aa1n03x5               g231(.a(new_n104), .b(new_n325), .c(new_n326), .d(new_n324), .out0(\s[4] ));
  nona22aa1n02x4               g232(.a(new_n110), .b(new_n104), .c(new_n111), .out0(new_n328));
  xorc02aa1n02x5               g233(.a(\a[5] ), .b(\b[4] ), .out0(new_n329));
  aoi012aa1n02x5               g234(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .o1(new_n330));
  oa0012aa1n02x5               g235(.a(new_n328), .b(new_n330), .c(new_n329), .o(\s[5] ));
  xorc02aa1n02x5               g236(.a(\a[6] ), .b(\b[5] ), .out0(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n332), .b(new_n328), .c(new_n118), .out0(\s[6] ));
  and002aa1n02x5               g238(.a(new_n332), .b(new_n118), .o(new_n334));
  aoi022aa1n02x5               g239(.a(new_n328), .b(new_n334), .c(\a[6] ), .d(\b[5] ), .o1(new_n335));
  aoi112aa1n02x5               g240(.a(new_n106), .b(new_n105), .c(\a[6] ), .d(\b[5] ), .o1(new_n336));
  aob012aa1n02x5               g241(.a(new_n336), .b(new_n328), .c(new_n334), .out0(new_n337));
  oa0012aa1n02x5               g242(.a(new_n337), .b(new_n335), .c(new_n117), .o(\s[7] ));
  xnbna2aa1n03x5               g243(.a(new_n116), .b(new_n337), .c(new_n120), .out0(\s[8] ));
  xorb03aa1n02x5               g244(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


