// Benchmark "adder" written by ABC on Wed Jul 17 21:07:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n320, new_n321, new_n322, new_n324, new_n325, new_n326,
    new_n328, new_n329, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  and002aa1n06x5               g003(.a(\b[2] ), .b(\a[3] ), .o(new_n99));
  nor002aa1n06x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nand42aa1n06x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand22aa1n12x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nor002aa1n20x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  oaih12aa1n12x5               g009(.a(new_n102), .b(new_n104), .c(new_n103), .o1(new_n105));
  xorc02aa1n12x5               g010(.a(\a[4] ), .b(\b[3] ), .out0(new_n106));
  oai112aa1n06x5               g011(.a(new_n106), .b(new_n101), .c(new_n105), .d(new_n99), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  aoi012aa1n02x7               g013(.a(new_n108), .b(\a[4] ), .c(\b[3] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1d28x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanb02aa1n02x5               g016(.a(new_n110), .b(new_n111), .out0(new_n112));
  aoi022aa1d24x5               g017(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\a[5] ), .o1(new_n114));
  inv040aa1d32x5               g019(.a(\b[4] ), .o1(new_n115));
  nor002aa1n16x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  inv000aa1n12x5               g021(.a(new_n116), .o1(new_n117));
  oai122aa1n06x5               g022(.a(new_n117), .b(\a[6] ), .c(\b[5] ), .d(new_n114), .e(new_n115), .o1(new_n118));
  nano23aa1n06x5               g023(.a(new_n118), .b(new_n112), .c(new_n109), .d(new_n113), .out0(new_n119));
  norb03aa1d15x5               g024(.a(new_n111), .b(new_n110), .c(new_n116), .out0(new_n120));
  nanp02aa1n04x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nor002aa1d32x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  nona22aa1n09x5               g027(.a(new_n121), .b(new_n122), .c(new_n108), .out0(new_n123));
  nanp03aa1d12x5               g028(.a(new_n123), .b(new_n120), .c(new_n113), .o1(new_n124));
  oaib12aa1n18x5               g029(.a(new_n124), .b(new_n120), .c(new_n111), .out0(new_n125));
  nand42aa1n16x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n97), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n107), .d(new_n119), .o1(new_n128));
  nor002aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  oai022aa1d18x5               g036(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n132));
  nanb03aa1n02x5               g037(.a(new_n132), .b(new_n128), .c(new_n130), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n131), .c(new_n98), .d(new_n128), .o1(\s[10] ));
  nanp02aa1n03x5               g039(.a(new_n119), .b(new_n107), .o1(new_n135));
  nanb02aa1n03x5               g040(.a(new_n125), .b(new_n135), .out0(new_n136));
  nano23aa1n06x5               g041(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n126), .out0(new_n137));
  aoi022aa1n06x5               g042(.a(new_n136), .b(new_n137), .c(new_n130), .d(new_n132), .o1(new_n138));
  nor002aa1n12x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n138), .b(new_n141), .c(new_n140), .out0(\s[11] ));
  norb02aa1n02x5               g047(.a(new_n141), .b(new_n139), .out0(new_n143));
  nanb02aa1n02x5               g048(.a(new_n138), .b(new_n143), .out0(new_n144));
  nor042aa1n02x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand02aa1n08x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  norb03aa1n02x5               g052(.a(new_n146), .b(new_n139), .c(new_n145), .out0(new_n148));
  oaib12aa1n02x5               g053(.a(new_n148), .b(new_n138), .c(new_n143), .out0(new_n149));
  aoai13aa1n03x5               g054(.a(new_n149), .b(new_n147), .c(new_n144), .d(new_n140), .o1(\s[12] ));
  inv000aa1d42x5               g055(.a(new_n125), .o1(new_n151));
  nano23aa1n06x5               g056(.a(new_n139), .b(new_n145), .c(new_n146), .d(new_n141), .out0(new_n152));
  nand22aa1n04x5               g057(.a(new_n152), .b(new_n137), .o1(new_n153));
  oai022aa1d18x5               g058(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n154));
  aoi022aa1d24x5               g059(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n155));
  aoai13aa1n12x5               g060(.a(new_n146), .b(new_n154), .c(new_n132), .d(new_n155), .o1(new_n156));
  aoai13aa1n02x5               g061(.a(new_n156), .b(new_n153), .c(new_n151), .d(new_n135), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nanp02aa1n04x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nanp03aa1n03x5               g066(.a(new_n157), .b(new_n160), .c(new_n161), .o1(new_n162));
  nor002aa1n16x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand02aa1n06x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  nona23aa1n02x4               g070(.a(new_n162), .b(new_n164), .c(new_n163), .d(new_n159), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n165), .c(new_n160), .d(new_n162), .o1(\s[14] ));
  nona23aa1n12x5               g072(.a(new_n164), .b(new_n161), .c(new_n159), .d(new_n163), .out0(new_n168));
  oai012aa1n12x5               g073(.a(new_n164), .b(new_n163), .c(new_n159), .o1(new_n169));
  oai012aa1d24x5               g074(.a(new_n169), .b(new_n156), .c(new_n168), .o1(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  nona22aa1n02x4               g076(.a(new_n136), .b(new_n153), .c(new_n168), .out0(new_n172));
  nor022aa1n06x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1d28x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n172), .c(new_n171), .out0(\s[15] ));
  nand02aa1n02x5               g081(.a(new_n172), .b(new_n171), .o1(new_n177));
  tech160nm_fiaoi012aa1n02p5x5 g082(.a(new_n173), .b(new_n177), .c(new_n174), .o1(new_n178));
  nor002aa1n04x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand42aa1d28x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  norb03aa1n02x5               g086(.a(new_n180), .b(new_n173), .c(new_n179), .out0(new_n182));
  aob012aa1n02x5               g087(.a(new_n182), .b(new_n177), .c(new_n175), .out0(new_n183));
  oai012aa1n02x5               g088(.a(new_n183), .b(new_n178), .c(new_n181), .o1(\s[16] ));
  nano23aa1n02x5               g089(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n161), .out0(new_n185));
  nano23aa1n06x5               g090(.a(new_n173), .b(new_n179), .c(new_n180), .d(new_n174), .out0(new_n186));
  nano22aa1n03x7               g091(.a(new_n153), .b(new_n185), .c(new_n186), .out0(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n125), .c(new_n107), .d(new_n119), .o1(new_n188));
  oai022aa1n02x5               g093(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n189));
  aoi022aa1d18x5               g094(.a(new_n170), .b(new_n186), .c(new_n180), .d(new_n189), .o1(new_n190));
  xorc02aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n190), .c(new_n188), .out0(\s[17] ));
  norp02aa1n24x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  nanp02aa1n24x5               g099(.a(new_n190), .b(new_n188), .o1(new_n195));
  nanp02aa1n06x5               g100(.a(new_n195), .b(new_n191), .o1(new_n196));
  xorc02aa1n02x5               g101(.a(\a[18] ), .b(\b[17] ), .out0(new_n197));
  nand42aa1n16x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  oai022aa1d18x5               g103(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n199));
  nanb03aa1n03x5               g104(.a(new_n199), .b(new_n196), .c(new_n198), .out0(new_n200));
  aoai13aa1n03x5               g105(.a(new_n200), .b(new_n197), .c(new_n194), .d(new_n196), .o1(\s[18] ));
  nand42aa1n20x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  nor042aa1n03x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nano23aa1d15x5               g108(.a(new_n193), .b(new_n203), .c(new_n198), .d(new_n202), .out0(new_n204));
  oaoi03aa1n02x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n194), .o1(new_n205));
  xorc02aa1n12x5               g110(.a(\a[19] ), .b(\b[18] ), .out0(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n205), .c(new_n195), .d(new_n204), .o1(new_n207));
  aoi112aa1n02x5               g112(.a(new_n206), .b(new_n205), .c(new_n195), .d(new_n204), .o1(new_n208));
  norb02aa1n03x4               g113(.a(new_n207), .b(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g115(.a(\a[19] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(\b[18] ), .o1(new_n212));
  nanp02aa1n02x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  xorc02aa1n12x5               g118(.a(\a[20] ), .b(\b[19] ), .out0(new_n214));
  nand02aa1d06x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  oai022aa1n02x5               g121(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n217));
  nona22aa1n02x5               g122(.a(new_n207), .b(new_n216), .c(new_n217), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n214), .c(new_n213), .d(new_n207), .o1(\s[20] ));
  nand23aa1n06x5               g124(.a(new_n204), .b(new_n206), .c(new_n214), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  oai112aa1n02x5               g126(.a(new_n199), .b(new_n198), .c(new_n212), .d(new_n211), .o1(new_n222));
  aoib12aa1n02x5               g127(.a(new_n216), .b(new_n222), .c(new_n217), .out0(new_n223));
  orn002aa1n24x5               g128(.a(\a[21] ), .b(\b[20] ), .o(new_n224));
  nanp02aa1n06x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  nand42aa1n06x5               g130(.a(new_n224), .b(new_n225), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n223), .c(new_n195), .d(new_n221), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n227), .b(new_n223), .c(new_n195), .d(new_n221), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n228), .b(new_n229), .out0(\s[21] ));
  xnrc02aa1n12x5               g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  and002aa1n02x5               g137(.a(\b[21] ), .b(\a[22] ), .o(new_n233));
  oai022aa1n02x5               g138(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n234));
  nona22aa1n02x5               g139(.a(new_n228), .b(new_n233), .c(new_n234), .out0(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n232), .c(new_n224), .d(new_n228), .o1(\s[22] ));
  nor022aa1n04x5               g141(.a(new_n231), .b(new_n226), .o1(new_n237));
  norb02aa1n09x5               g142(.a(new_n237), .b(new_n220), .out0(new_n238));
  nanb02aa1n02x5               g143(.a(new_n217), .b(new_n222), .out0(new_n239));
  nano32aa1n03x7               g144(.a(new_n231), .b(new_n224), .c(new_n225), .d(new_n215), .out0(new_n240));
  nanp02aa1n02x5               g145(.a(new_n239), .b(new_n240), .o1(new_n241));
  oaib12aa1n02x5               g146(.a(new_n241), .b(new_n233), .c(new_n234), .out0(new_n242));
  xorc02aa1n12x5               g147(.a(\a[23] ), .b(\b[22] ), .out0(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n242), .c(new_n195), .d(new_n238), .o1(new_n244));
  oaoi03aa1n02x5               g149(.a(\a[22] ), .b(\b[21] ), .c(new_n224), .o1(new_n245));
  nona22aa1n02x4               g150(.a(new_n241), .b(new_n245), .c(new_n243), .out0(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(new_n195), .c(new_n238), .o1(new_n247));
  norb02aa1n03x4               g152(.a(new_n244), .b(new_n247), .out0(\s[23] ));
  norp02aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  tech160nm_fixorc02aa1n02p5x5 g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  and002aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o(new_n252));
  oai022aa1n02x5               g157(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n253));
  nona22aa1n02x5               g158(.a(new_n244), .b(new_n252), .c(new_n253), .out0(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n251), .c(new_n250), .d(new_n244), .o1(\s[24] ));
  nano32aa1n02x5               g160(.a(new_n220), .b(new_n251), .c(new_n237), .d(new_n243), .out0(new_n256));
  and002aa1n02x5               g161(.a(new_n251), .b(new_n243), .o(new_n257));
  aoai13aa1n04x5               g162(.a(new_n257), .b(new_n245), .c(new_n239), .d(new_n240), .o1(new_n258));
  aob012aa1n02x5               g163(.a(new_n253), .b(\b[23] ), .c(\a[24] ), .out0(new_n259));
  nanp02aa1n02x5               g164(.a(new_n258), .b(new_n259), .o1(new_n260));
  xnrc02aa1n12x5               g165(.a(\b[24] ), .b(\a[25] ), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n262), .b(new_n260), .c(new_n195), .d(new_n256), .o1(new_n263));
  aoi112aa1n02x5               g168(.a(new_n262), .b(new_n260), .c(new_n195), .d(new_n256), .o1(new_n264));
  norb02aa1n03x4               g169(.a(new_n263), .b(new_n264), .out0(\s[25] ));
  norp02aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  and002aa1n02x5               g173(.a(\b[25] ), .b(\a[26] ), .o(new_n269));
  oai022aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n270));
  nona22aa1n02x5               g175(.a(new_n263), .b(new_n269), .c(new_n270), .out0(new_n271));
  aoai13aa1n03x5               g176(.a(new_n271), .b(new_n268), .c(new_n267), .d(new_n263), .o1(\s[26] ));
  norb02aa1n02x5               g177(.a(new_n268), .b(new_n261), .out0(new_n273));
  nand03aa1n03x5               g178(.a(new_n238), .b(new_n257), .c(new_n273), .o1(new_n274));
  inv040aa1n06x5               g179(.a(new_n274), .o1(new_n275));
  inv000aa1n02x5               g180(.a(new_n273), .o1(new_n276));
  aob012aa1n02x5               g181(.a(new_n270), .b(\b[25] ), .c(\a[26] ), .out0(new_n277));
  aoai13aa1n12x5               g182(.a(new_n277), .b(new_n276), .c(new_n258), .d(new_n259), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  aoai13aa1n06x5               g184(.a(new_n279), .b(new_n278), .c(new_n195), .d(new_n275), .o1(new_n280));
  aoi112aa1n02x5               g185(.a(new_n279), .b(new_n278), .c(new_n195), .d(new_n275), .o1(new_n281));
  norb02aa1n03x4               g186(.a(new_n280), .b(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g187(.a(\b[26] ), .b(\a[27] ), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[28] ), .b(\b[27] ), .out0(new_n285));
  oai022aa1d24x5               g190(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n286));
  aoi012aa1n02x5               g191(.a(new_n286), .b(\a[28] ), .c(\b[27] ), .o1(new_n287));
  tech160nm_finand02aa1n03p5x5 g192(.a(new_n280), .b(new_n287), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n285), .c(new_n284), .d(new_n280), .o1(\s[28] ));
  xorc02aa1n02x5               g194(.a(\a[29] ), .b(\b[28] ), .out0(new_n290));
  and002aa1n02x5               g195(.a(new_n285), .b(new_n279), .o(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n278), .c(new_n195), .d(new_n275), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\b[27] ), .o1(new_n293));
  oaib12aa1n09x5               g198(.a(new_n286), .b(new_n293), .c(\a[28] ), .out0(new_n294));
  nanp03aa1n03x5               g199(.a(new_n292), .b(new_n294), .c(new_n290), .o1(new_n295));
  aoi012aa1n06x5               g200(.a(new_n274), .b(new_n190), .c(new_n188), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n294), .o1(new_n297));
  oaoi13aa1n03x5               g202(.a(new_n297), .b(new_n291), .c(new_n296), .d(new_n278), .o1(new_n298));
  oaih12aa1n02x5               g203(.a(new_n295), .b(new_n298), .c(new_n290), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g205(.a(new_n279), .b(new_n290), .c(new_n285), .o(new_n301));
  tech160nm_fioaoi03aa1n03p5x5 g206(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .o1(new_n302));
  oaoi13aa1n03x5               g207(.a(new_n302), .b(new_n301), .c(new_n296), .d(new_n278), .o1(new_n303));
  xorc02aa1n02x5               g208(.a(\a[30] ), .b(\b[29] ), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n301), .b(new_n278), .c(new_n195), .d(new_n275), .o1(new_n305));
  norb02aa1n02x5               g210(.a(new_n304), .b(new_n302), .out0(new_n306));
  nand42aa1n02x5               g211(.a(new_n305), .b(new_n306), .o1(new_n307));
  oaih12aa1n02x5               g212(.a(new_n307), .b(new_n303), .c(new_n304), .o1(\s[30] ));
  and003aa1n02x5               g213(.a(new_n291), .b(new_n304), .c(new_n290), .o(new_n309));
  aoi012aa1n02x5               g214(.a(new_n306), .b(\a[30] ), .c(\b[29] ), .o1(new_n310));
  oaoi13aa1n03x5               g215(.a(new_n310), .b(new_n309), .c(new_n296), .d(new_n278), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[31] ), .b(\b[30] ), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n309), .b(new_n278), .c(new_n195), .d(new_n275), .o1(new_n313));
  norb02aa1n02x5               g218(.a(new_n312), .b(new_n310), .out0(new_n314));
  nand42aa1n02x5               g219(.a(new_n313), .b(new_n314), .o1(new_n315));
  oaih12aa1n02x5               g220(.a(new_n315), .b(new_n311), .c(new_n312), .o1(\s[31] ));
  xnrb03aa1n02x5               g221(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oab012aa1n02x4               g222(.a(new_n100), .b(new_n105), .c(new_n99), .out0(new_n318));
  oai012aa1n02x5               g223(.a(new_n107), .b(new_n318), .c(new_n106), .o1(\s[4] ));
  aob012aa1n02x5               g224(.a(new_n107), .b(\b[3] ), .c(\a[4] ), .out0(new_n320));
  xnrc02aa1n02x5               g225(.a(\b[4] ), .b(\a[5] ), .out0(new_n321));
  oai112aa1n02x5               g226(.a(new_n107), .b(new_n109), .c(new_n115), .d(new_n114), .o1(new_n322));
  aobi12aa1n02x5               g227(.a(new_n322), .b(new_n321), .c(new_n320), .out0(\s[5] ));
  nanb02aa1n02x5               g228(.a(new_n122), .b(new_n121), .out0(new_n324));
  oaib12aa1n02x5               g229(.a(new_n322), .b(\b[4] ), .c(new_n114), .out0(new_n325));
  nanb02aa1n06x5               g230(.a(new_n123), .b(new_n322), .out0(new_n326));
  aob012aa1n02x5               g231(.a(new_n326), .b(new_n325), .c(new_n324), .out0(\s[6] ));
  nanp02aa1n02x5               g232(.a(\b[6] ), .b(\a[7] ), .o1(new_n328));
  aoi022aa1n02x5               g233(.a(new_n326), .b(new_n121), .c(new_n328), .d(new_n117), .o1(new_n329));
  aoi013aa1n02x4               g234(.a(new_n329), .b(new_n326), .c(new_n117), .d(new_n113), .o1(\s[7] ));
  nanp03aa1n02x5               g235(.a(new_n326), .b(new_n113), .c(new_n117), .o1(new_n331));
  xobna2aa1n03x5               g236(.a(new_n112), .b(new_n331), .c(new_n117), .out0(\s[8] ));
  xnbna2aa1n03x5               g237(.a(new_n127), .b(new_n151), .c(new_n135), .out0(\s[9] ));
endmodule


