// Benchmark "adder" written by ABC on Thu Jul 18 08:51:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n149,
    new_n150, new_n152, new_n153, new_n154, new_n155, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n175, new_n176, new_n177, new_n178, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n306, new_n307, new_n308, new_n311, new_n313,
    new_n315;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n03p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1n04x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv030aa1n02x5               g003(.a(new_n98), .o1(new_n99));
  nor002aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  tech160nm_fiaoi012aa1n05x5   g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand02aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n09x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nona23aa1n09x5               g012(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n108));
  tech160nm_fiaoi012aa1n03p5x5 g013(.a(new_n104), .b(new_n106), .c(new_n105), .o1(new_n109));
  oai012aa1n12x5               g014(.a(new_n109), .b(new_n108), .c(new_n103), .o1(new_n110));
  nor022aa1n16x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n03x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .out0(new_n116));
  tech160nm_fixnrc02aa1n02p5x5 g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nor043aa1n06x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  inv040aa1d32x5               g023(.a(\a[5] ), .o1(new_n119));
  inv040aa1d28x5               g024(.a(\b[4] ), .o1(new_n120));
  nand22aa1n02x5               g025(.a(new_n120), .b(new_n119), .o1(new_n121));
  tech160nm_fioaoi03aa1n02p5x5 g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  aoi012aa1n06x5               g027(.a(new_n111), .b(new_n113), .c(new_n112), .o1(new_n123));
  oaib12aa1n09x5               g028(.a(new_n123), .b(new_n115), .c(new_n122), .out0(new_n124));
  tech160nm_fixorc02aa1n02p5x5 g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  and002aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  nor042aa1n04x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nand42aa1n04x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  oab012aa1n02x4               g036(.a(new_n98), .b(\a[10] ), .c(\b[9] ), .out0(new_n132));
  aoi112aa1n03x5               g037(.a(new_n131), .b(new_n128), .c(new_n126), .d(new_n132), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n131), .b(new_n128), .c(new_n126), .d(new_n132), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(\s[11] ));
  nor042aa1n03x5               g040(.a(new_n133), .b(new_n129), .o1(new_n136));
  xnrb03aa1n03x5               g041(.a(new_n136), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n03x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand42aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nano23aa1n06x5               g044(.a(new_n129), .b(new_n138), .c(new_n139), .d(new_n130), .out0(new_n140));
  and003aa1n02x5               g045(.a(new_n140), .b(new_n125), .c(new_n97), .o(new_n141));
  aoai13aa1n06x5               g046(.a(new_n141), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n142));
  oaoi03aa1n02x5               g047(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n143));
  aoi012aa1n02x5               g048(.a(new_n138), .b(new_n129), .c(new_n139), .o1(new_n144));
  aobi12aa1n12x5               g049(.a(new_n144), .b(new_n140), .c(new_n143), .out0(new_n145));
  xorc02aa1n12x5               g050(.a(\a[13] ), .b(\b[12] ), .out0(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n142), .c(new_n145), .out0(\s[13] ));
  orn002aa1n24x5               g052(.a(\a[13] ), .b(\b[12] ), .o(new_n148));
  aob012aa1n02x5               g053(.a(new_n146), .b(new_n142), .c(new_n145), .out0(new_n149));
  xorc02aa1n12x5               g054(.a(\a[14] ), .b(\b[13] ), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n149), .c(new_n148), .out0(\s[14] ));
  nanp02aa1n02x5               g056(.a(new_n150), .b(new_n146), .o1(new_n152));
  oaoi03aa1n12x5               g057(.a(\a[14] ), .b(\b[13] ), .c(new_n148), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n04x5               g059(.a(new_n154), .b(new_n152), .c(new_n142), .d(new_n145), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n04x5               g061(.a(\b[14] ), .b(\a[15] ), .o1(new_n157));
  nand42aa1d28x5               g062(.a(\b[14] ), .b(\a[15] ), .o1(new_n158));
  norp02aa1n04x5               g063(.a(\b[15] ), .b(\a[16] ), .o1(new_n159));
  nand02aa1d16x5               g064(.a(\b[15] ), .b(\a[16] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  aoai13aa1n02x5               g066(.a(new_n161), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n162));
  aoi112aa1n02x5               g067(.a(new_n157), .b(new_n161), .c(new_n155), .d(new_n158), .o1(new_n163));
  norb02aa1n02x7               g068(.a(new_n162), .b(new_n163), .out0(\s[16] ));
  nano23aa1n06x5               g069(.a(new_n157), .b(new_n159), .c(new_n160), .d(new_n158), .out0(new_n165));
  nand23aa1n04x5               g070(.a(new_n165), .b(new_n146), .c(new_n150), .o1(new_n166));
  nano32aa1n03x7               g071(.a(new_n166), .b(new_n140), .c(new_n125), .d(new_n97), .out0(new_n167));
  aoai13aa1n12x5               g072(.a(new_n167), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n168));
  tech160nm_fiao0012aa1n02p5x5 g073(.a(new_n159), .b(new_n157), .c(new_n160), .o(new_n169));
  aoi012aa1n06x5               g074(.a(new_n169), .b(new_n165), .c(new_n153), .o1(new_n170));
  inv040aa1n03x5               g075(.a(new_n170), .o1(new_n171));
  oab012aa1n12x5               g076(.a(new_n171), .b(new_n145), .c(new_n166), .out0(new_n172));
  nanp02aa1n09x5               g077(.a(new_n168), .b(new_n172), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g079(.a(\a[18] ), .o1(new_n175));
  inv000aa1d42x5               g080(.a(\a[17] ), .o1(new_n176));
  inv000aa1d42x5               g081(.a(\b[16] ), .o1(new_n177));
  oaoi03aa1n02x5               g082(.a(new_n176), .b(new_n177), .c(new_n173), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[17] ), .c(new_n175), .out0(\s[18] ));
  xroi22aa1d06x4               g084(.a(new_n176), .b(\b[16] ), .c(new_n175), .d(\b[17] ), .out0(new_n180));
  oai022aa1d24x5               g085(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n181));
  oaib12aa1n18x5               g086(.a(new_n181), .b(new_n175), .c(\b[17] ), .out0(new_n182));
  inv040aa1n08x5               g087(.a(new_n182), .o1(new_n183));
  aoi012aa1n12x5               g088(.a(new_n183), .b(new_n173), .c(new_n180), .o1(new_n184));
  nor042aa1d18x5               g089(.a(\b[18] ), .b(\a[19] ), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  nand02aa1n10x5               g091(.a(\b[18] ), .b(\a[19] ), .o1(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n184), .b(new_n187), .c(new_n186), .out0(\s[19] ));
  xnrc02aa1n02x5               g093(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g094(.a(new_n185), .b(new_n187), .out0(new_n190));
  nor042aa1n06x5               g095(.a(\b[19] ), .b(\a[20] ), .o1(new_n191));
  nand02aa1d16x5               g096(.a(\b[19] ), .b(\a[20] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  oaoi13aa1n06x5               g098(.a(new_n193), .b(new_n186), .c(new_n184), .d(new_n190), .o1(new_n194));
  nor042aa1n04x5               g099(.a(new_n184), .b(new_n190), .o1(new_n195));
  nano22aa1n03x5               g100(.a(new_n195), .b(new_n186), .c(new_n193), .out0(new_n196));
  norp02aa1n03x5               g101(.a(new_n194), .b(new_n196), .o1(\s[20] ));
  nano23aa1n09x5               g102(.a(new_n185), .b(new_n191), .c(new_n192), .d(new_n187), .out0(new_n198));
  nanp02aa1n02x5               g103(.a(new_n180), .b(new_n198), .o1(new_n199));
  nona23aa1d18x5               g104(.a(new_n192), .b(new_n187), .c(new_n185), .d(new_n191), .out0(new_n200));
  aoi012aa1d24x5               g105(.a(new_n191), .b(new_n185), .c(new_n192), .o1(new_n201));
  oai012aa1d24x5               g106(.a(new_n201), .b(new_n200), .c(new_n182), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n199), .c(new_n168), .d(new_n172), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g110(.a(\b[20] ), .b(\a[21] ), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[21] ), .b(\b[20] ), .out0(new_n207));
  xorc02aa1n02x5               g112(.a(\a[22] ), .b(\b[21] ), .out0(new_n208));
  aoai13aa1n03x5               g113(.a(new_n208), .b(new_n206), .c(new_n204), .d(new_n207), .o1(new_n209));
  aoi112aa1n02x5               g114(.a(new_n206), .b(new_n208), .c(new_n204), .d(new_n207), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n209), .b(new_n210), .out0(\s[22] ));
  inv000aa1d42x5               g116(.a(\a[21] ), .o1(new_n212));
  inv040aa1d32x5               g117(.a(\a[22] ), .o1(new_n213));
  xroi22aa1d06x4               g118(.a(new_n212), .b(\b[20] ), .c(new_n213), .d(\b[21] ), .out0(new_n214));
  nand23aa1n02x5               g119(.a(new_n214), .b(new_n180), .c(new_n198), .o1(new_n215));
  inv000aa1d42x5               g120(.a(\b[21] ), .o1(new_n216));
  oao003aa1n02x5               g121(.a(new_n213), .b(new_n216), .c(new_n206), .carry(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(new_n202), .c(new_n214), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n215), .c(new_n168), .d(new_n172), .o1(new_n219));
  xorb03aa1n02x5               g124(.a(new_n219), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g125(.a(\b[22] ), .b(\a[23] ), .o1(new_n221));
  tech160nm_fixorc02aa1n05x5   g126(.a(\a[23] ), .b(\b[22] ), .out0(new_n222));
  tech160nm_fixorc02aa1n02p5x5 g127(.a(\a[24] ), .b(\b[23] ), .out0(new_n223));
  aoai13aa1n03x5               g128(.a(new_n223), .b(new_n221), .c(new_n219), .d(new_n222), .o1(new_n224));
  aoi112aa1n02x5               g129(.a(new_n221), .b(new_n223), .c(new_n219), .d(new_n222), .o1(new_n225));
  norb02aa1n02x7               g130(.a(new_n224), .b(new_n225), .out0(\s[24] ));
  norb02aa1n02x5               g131(.a(new_n105), .b(new_n104), .out0(new_n227));
  norb02aa1n02x5               g132(.a(new_n107), .b(new_n106), .out0(new_n228));
  nanb03aa1n02x5               g133(.a(new_n103), .b(new_n228), .c(new_n227), .out0(new_n229));
  nano23aa1n03x7               g134(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n230));
  nona22aa1n02x4               g135(.a(new_n230), .b(new_n116), .c(new_n117), .out0(new_n231));
  aobi12aa1n06x5               g136(.a(new_n123), .b(new_n230), .c(new_n122), .out0(new_n232));
  aoai13aa1n04x5               g137(.a(new_n232), .b(new_n231), .c(new_n229), .d(new_n109), .o1(new_n233));
  tech160nm_fioai012aa1n03p5x5 g138(.a(new_n170), .b(new_n145), .c(new_n166), .o1(new_n234));
  and002aa1n06x5               g139(.a(new_n223), .b(new_n222), .o(new_n235));
  inv000aa1n02x5               g140(.a(new_n235), .o1(new_n236));
  nano32aa1n02x4               g141(.a(new_n236), .b(new_n214), .c(new_n180), .d(new_n198), .out0(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n233), .d(new_n167), .o1(new_n238));
  inv020aa1n03x5               g143(.a(new_n201), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n214), .b(new_n239), .c(new_n198), .d(new_n183), .o1(new_n240));
  inv000aa1n02x5               g145(.a(new_n217), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n242));
  oab012aa1n02x4               g147(.a(new_n242), .b(\a[24] ), .c(\b[23] ), .out0(new_n243));
  aoai13aa1n12x5               g148(.a(new_n243), .b(new_n236), .c(new_n240), .d(new_n241), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[24] ), .b(\a[25] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xnbna2aa1n03x5               g152(.a(new_n247), .b(new_n238), .c(new_n245), .out0(\s[25] ));
  nor042aa1n03x5               g153(.a(\b[24] ), .b(\a[25] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n247), .b(new_n244), .c(new_n173), .d(new_n237), .o1(new_n251));
  xnrc02aa1n12x5               g156(.a(\b[25] ), .b(\a[26] ), .out0(new_n252));
  tech160nm_fiaoi012aa1n05x5   g157(.a(new_n252), .b(new_n251), .c(new_n250), .o1(new_n253));
  nanp03aa1n06x5               g158(.a(new_n251), .b(new_n250), .c(new_n252), .o1(new_n254));
  norb02aa1n03x4               g159(.a(new_n254), .b(new_n253), .out0(\s[26] ));
  nor042aa1n06x5               g160(.a(new_n252), .b(new_n246), .o1(new_n256));
  nano22aa1n02x5               g161(.a(new_n215), .b(new_n235), .c(new_n256), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n234), .c(new_n233), .d(new_n167), .o1(new_n258));
  nanp02aa1n09x5               g163(.a(new_n244), .b(new_n256), .o1(new_n259));
  oao003aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .c(new_n250), .carry(new_n260));
  xorc02aa1n12x5               g165(.a(\a[27] ), .b(\b[26] ), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoi013aa1n06x4               g167(.a(new_n262), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n263));
  aobi12aa1n06x5               g168(.a(new_n257), .b(new_n168), .c(new_n172), .out0(new_n264));
  aoai13aa1n04x5               g169(.a(new_n235), .b(new_n217), .c(new_n202), .d(new_n214), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n256), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n260), .b(new_n266), .c(new_n265), .d(new_n243), .o1(new_n267));
  norp03aa1n02x5               g172(.a(new_n267), .b(new_n264), .c(new_n261), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n263), .b(new_n268), .o1(\s[27] ));
  norp02aa1n02x5               g174(.a(\b[26] ), .b(\a[27] ), .o1(new_n270));
  inv040aa1n03x5               g175(.a(new_n270), .o1(new_n271));
  oaih12aa1n02x5               g176(.a(new_n261), .b(new_n267), .c(new_n264), .o1(new_n272));
  xnrc02aa1n02x5               g177(.a(\b[27] ), .b(\a[28] ), .out0(new_n273));
  tech160nm_fiaoi012aa1n02p5x5 g178(.a(new_n273), .b(new_n272), .c(new_n271), .o1(new_n274));
  nano22aa1n03x5               g179(.a(new_n263), .b(new_n271), .c(new_n273), .out0(new_n275));
  norp02aa1n03x5               g180(.a(new_n274), .b(new_n275), .o1(\s[28] ));
  norb02aa1n02x5               g181(.a(new_n261), .b(new_n273), .out0(new_n277));
  oaih12aa1n02x5               g182(.a(new_n277), .b(new_n267), .c(new_n264), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[28] ), .b(\b[27] ), .c(new_n271), .carry(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[28] ), .b(\a[29] ), .out0(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n278), .c(new_n279), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n277), .o1(new_n282));
  aoi013aa1n03x5               g187(.a(new_n282), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n283));
  nano22aa1n03x5               g188(.a(new_n283), .b(new_n279), .c(new_n280), .out0(new_n284));
  norp02aa1n03x5               g189(.a(new_n281), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g190(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n06x5               g191(.a(new_n261), .b(new_n280), .c(new_n273), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n267), .c(new_n264), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n279), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n03p5x5 g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n287), .o1(new_n292));
  aoi013aa1n03x5               g197(.a(new_n292), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n290), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n291), .b(new_n294), .o1(\s[30] ));
  norb02aa1n02x5               g200(.a(new_n287), .b(new_n290), .out0(new_n296));
  inv000aa1n02x5               g201(.a(new_n296), .o1(new_n297));
  aoi013aa1n03x5               g202(.a(new_n297), .b(new_n259), .c(new_n258), .d(new_n260), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n300), .out0(new_n301));
  oaih12aa1n02x5               g206(.a(new_n296), .b(new_n267), .c(new_n264), .o1(new_n302));
  tech160nm_fiaoi012aa1n02p5x5 g207(.a(new_n300), .b(new_n302), .c(new_n299), .o1(new_n303));
  norp02aa1n03x5               g208(.a(new_n303), .b(new_n301), .o1(\s[31] ));
  xnrb03aa1n02x5               g209(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g210(.a(new_n104), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n228), .b(new_n100), .c(new_n102), .d(new_n101), .o1(new_n307));
  aoi012aa1n02x5               g212(.a(new_n106), .b(new_n306), .c(new_n105), .o1(new_n308));
  aoi022aa1n02x5               g213(.a(new_n110), .b(new_n306), .c(new_n307), .d(new_n308), .o1(\s[4] ));
  xorb03aa1n02x5               g214(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g215(.a(new_n119), .b(new_n120), .c(new_n110), .o1(new_n311));
  xnrb03aa1n02x5               g216(.a(new_n311), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g217(.a(\a[6] ), .b(\b[5] ), .c(new_n311), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g219(.a(new_n113), .b(new_n313), .c(new_n114), .o1(new_n315));
  xnrb03aa1n02x5               g220(.a(new_n315), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g221(.a(new_n233), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


