// Benchmark "adder" written by ABC on Wed Jul 17 21:56:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n348, new_n350, new_n353, new_n354,
    new_n356, new_n357;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d10x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1d24x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor042aa1n04x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  xnrc02aa1n03x5               g005(.a(\b[3] ), .b(\a[4] ), .out0(new_n101));
  nand42aa1n08x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb03aa1n12x5               g009(.a(new_n103), .b(new_n104), .c(new_n102), .out0(new_n105));
  nand02aa1n03x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  norb03aa1n03x5               g012(.a(new_n102), .b(new_n107), .c(new_n106), .out0(new_n108));
  inv020aa1n02x5               g013(.a(new_n108), .o1(new_n109));
  nona22aa1n06x5               g014(.a(new_n109), .b(new_n105), .c(new_n101), .out0(new_n110));
  inv000aa1n02x5               g015(.a(new_n103), .o1(new_n111));
  oao003aa1n09x5               g016(.a(\a[4] ), .b(\b[3] ), .c(new_n111), .carry(new_n112));
  nor042aa1d18x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  norb02aa1n03x5               g019(.a(new_n114), .b(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  nanp02aa1n06x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  norp02aa1n24x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  tech160nm_fixorc02aa1n03p5x5 g024(.a(\a[8] ), .b(\b[7] ), .out0(new_n120));
  nona23aa1n06x5               g025(.a(new_n120), .b(new_n115), .c(new_n116), .d(new_n119), .out0(new_n121));
  inv040aa1d32x5               g026(.a(\a[8] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[7] ), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(new_n122), .b(new_n123), .c(new_n113), .o1(new_n124));
  inv000aa1n03x5               g029(.a(new_n113), .o1(new_n125));
  oai112aa1n03x5               g030(.a(new_n125), .b(new_n114), .c(new_n123), .d(new_n122), .o1(new_n126));
  oaih22aa1d12x5               g031(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n127));
  oai112aa1n06x5               g032(.a(new_n127), .b(new_n117), .c(\b[7] ), .d(\a[8] ), .o1(new_n128));
  tech160nm_fioai012aa1n04x5   g033(.a(new_n124), .b(new_n128), .c(new_n126), .o1(new_n129));
  inv040aa1n02x5               g034(.a(new_n129), .o1(new_n130));
  aoai13aa1n12x5               g035(.a(new_n130), .b(new_n121), .c(new_n110), .d(new_n112), .o1(new_n131));
  xorc02aa1n12x5               g036(.a(\a[9] ), .b(\b[8] ), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n99), .b(new_n100), .c(new_n131), .d(new_n132), .o1(new_n133));
  oai013aa1n03x5               g038(.a(new_n112), .b(new_n108), .c(new_n105), .d(new_n101), .o1(new_n134));
  xorc02aa1n02x5               g039(.a(\a[5] ), .b(\b[4] ), .out0(new_n135));
  nanp02aa1n02x5               g040(.a(new_n135), .b(new_n115), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n118), .o1(new_n137));
  nano32aa1n03x7               g042(.a(new_n136), .b(new_n120), .c(new_n117), .d(new_n137), .out0(new_n138));
  aoai13aa1n02x5               g043(.a(new_n132), .b(new_n129), .c(new_n134), .d(new_n138), .o1(new_n139));
  norb03aa1n02x5               g044(.a(new_n98), .b(new_n97), .c(new_n100), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n139), .b(new_n140), .o1(new_n141));
  nanp02aa1n02x5               g046(.a(new_n133), .b(new_n141), .o1(\s[10] ));
  nand42aa1n08x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nor002aa1d32x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nanb03aa1n02x5               g049(.a(new_n144), .b(new_n98), .c(new_n143), .out0(new_n145));
  nanb02aa1n02x5               g050(.a(new_n145), .b(new_n141), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n144), .o1(new_n147));
  aoi022aa1n02x5               g052(.a(new_n141), .b(new_n98), .c(new_n147), .d(new_n143), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n146), .b(new_n148), .out0(\s[11] ));
  nor002aa1d32x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand02aa1d16x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  norb02aa1n06x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n150), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n144), .b(new_n153), .c(new_n151), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n147), .b(new_n145), .c(new_n139), .d(new_n140), .o1(new_n155));
  aoi022aa1n02x5               g060(.a(new_n146), .b(new_n154), .c(new_n155), .d(new_n152), .o1(\s[12] ));
  nanb02aa1n12x5               g061(.a(new_n144), .b(new_n143), .out0(new_n157));
  nona23aa1d24x5               g062(.a(new_n152), .b(new_n132), .c(new_n99), .d(new_n157), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n02x5               g064(.a(new_n159), .b(new_n129), .c(new_n134), .d(new_n138), .o1(new_n160));
  nanb03aa1n06x5               g065(.a(new_n150), .b(new_n151), .c(new_n143), .out0(new_n161));
  oai112aa1n06x5               g066(.a(new_n147), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n162));
  aoi012aa1n09x5               g067(.a(new_n150), .b(new_n144), .c(new_n151), .o1(new_n163));
  oai012aa1n18x5               g068(.a(new_n163), .b(new_n162), .c(new_n161), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nor042aa1n04x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  nanp02aa1n04x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n160), .c(new_n165), .out0(\s[13] ));
  nand02aa1n03x5               g074(.a(new_n160), .b(new_n165), .o1(new_n170));
  nor042aa1n03x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1n04x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(new_n166), .b(new_n173), .c(new_n170), .d(new_n168), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n173), .b(new_n166), .c(new_n170), .d(new_n167), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[14] ));
  nano23aa1n09x5               g081(.a(new_n166), .b(new_n171), .c(new_n172), .d(new_n167), .out0(new_n177));
  aoai13aa1n06x5               g082(.a(new_n177), .b(new_n164), .c(new_n131), .d(new_n159), .o1(new_n178));
  oai012aa1n12x5               g083(.a(new_n172), .b(new_n171), .c(new_n166), .o1(new_n179));
  xnrc02aa1n12x5               g084(.a(\b[14] ), .b(\a[15] ), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n178), .c(new_n179), .out0(\s[15] ));
  inv000aa1d42x5               g087(.a(new_n179), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n181), .b(new_n183), .c(new_n170), .d(new_n177), .o1(new_n184));
  xnrc02aa1n12x5               g089(.a(\b[15] ), .b(\a[16] ), .out0(new_n185));
  inv000aa1d42x5               g090(.a(new_n185), .o1(new_n186));
  nor042aa1n06x5               g091(.a(\b[14] ), .b(\a[15] ), .o1(new_n187));
  norb02aa1n02x5               g092(.a(new_n185), .b(new_n187), .out0(new_n188));
  inv000aa1d42x5               g093(.a(new_n187), .o1(new_n189));
  aoai13aa1n02x5               g094(.a(new_n189), .b(new_n180), .c(new_n178), .d(new_n179), .o1(new_n190));
  aoi022aa1n03x5               g095(.a(new_n190), .b(new_n186), .c(new_n184), .d(new_n188), .o1(\s[16] ));
  norp02aa1n24x5               g096(.a(new_n185), .b(new_n180), .o1(new_n192));
  nano22aa1d15x5               g097(.a(new_n158), .b(new_n177), .c(new_n192), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n129), .c(new_n134), .d(new_n138), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n192), .b(new_n183), .c(new_n164), .d(new_n177), .o1(new_n195));
  oao003aa1n02x5               g100(.a(\a[16] ), .b(\b[15] ), .c(new_n189), .carry(new_n196));
  nanp03aa1d12x5               g101(.a(new_n194), .b(new_n195), .c(new_n196), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  nano22aa1n02x4               g103(.a(new_n198), .b(new_n195), .c(new_n196), .out0(new_n199));
  aoi022aa1n02x5               g104(.a(new_n197), .b(new_n198), .c(new_n199), .d(new_n194), .o1(\s[17] ));
  inv000aa1d42x5               g105(.a(\a[17] ), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(\b[16] ), .b(new_n201), .out0(new_n202));
  inv000aa1n02x5               g107(.a(new_n192), .o1(new_n203));
  nano22aa1n02x4               g108(.a(new_n150), .b(new_n143), .c(new_n151), .out0(new_n204));
  oai012aa1n02x5               g109(.a(new_n98), .b(\b[10] ), .c(\a[11] ), .o1(new_n205));
  oab012aa1n04x5               g110(.a(new_n205), .b(new_n97), .c(new_n100), .out0(new_n206));
  inv020aa1n03x5               g111(.a(new_n163), .o1(new_n207));
  aoai13aa1n06x5               g112(.a(new_n177), .b(new_n207), .c(new_n206), .d(new_n204), .o1(new_n208));
  aoai13aa1n06x5               g113(.a(new_n196), .b(new_n203), .c(new_n208), .d(new_n179), .o1(new_n209));
  aoai13aa1n03x5               g114(.a(new_n198), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n210));
  norp02aa1n12x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nand02aa1d12x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  norb02aa1n06x4               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n210), .c(new_n202), .out0(\s[18] ));
  and002aa1n02x5               g119(.a(new_n198), .b(new_n213), .o(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n216));
  oaoi03aa1n02x5               g121(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  nor002aa1d32x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  nand42aa1n08x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  norb02aa1n12x5               g125(.a(new_n220), .b(new_n219), .out0(new_n221));
  xnbna2aa1n03x5               g126(.a(new_n221), .b(new_n216), .c(new_n218), .out0(\s[19] ));
  xnrc02aa1n02x5               g127(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g128(.a(new_n221), .b(new_n217), .c(new_n197), .d(new_n215), .o1(new_n224));
  nor002aa1d32x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand42aa1d28x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n06x4               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  inv000aa1d42x5               g132(.a(\a[19] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\b[18] ), .o1(new_n229));
  aboi22aa1n03x5               g134(.a(new_n225), .b(new_n226), .c(new_n228), .d(new_n229), .out0(new_n230));
  inv030aa1n06x5               g135(.a(new_n219), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n221), .o1(new_n232));
  aoai13aa1n02x5               g137(.a(new_n231), .b(new_n232), .c(new_n216), .d(new_n218), .o1(new_n233));
  aoi022aa1n03x5               g138(.a(new_n233), .b(new_n227), .c(new_n224), .d(new_n230), .o1(\s[20] ));
  nano32aa1n03x7               g139(.a(new_n232), .b(new_n198), .c(new_n227), .d(new_n213), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n236));
  nanb03aa1n09x5               g141(.a(new_n225), .b(new_n226), .c(new_n220), .out0(new_n237));
  nor042aa1n06x5               g142(.a(\b[16] ), .b(\a[17] ), .o1(new_n238));
  oai112aa1n06x5               g143(.a(new_n231), .b(new_n212), .c(new_n211), .d(new_n238), .o1(new_n239));
  aoi012aa1d18x5               g144(.a(new_n225), .b(new_n219), .c(new_n226), .o1(new_n240));
  oai012aa1d24x5               g145(.a(new_n240), .b(new_n239), .c(new_n237), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  nor042aa1d18x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  nand42aa1n10x5               g148(.a(\b[20] ), .b(\a[21] ), .o1(new_n244));
  norb02aa1n12x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  xnbna2aa1n03x5               g150(.a(new_n245), .b(new_n236), .c(new_n242), .out0(\s[21] ));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n241), .c(new_n197), .d(new_n235), .o1(new_n247));
  nor042aa1n06x5               g152(.a(\b[21] ), .b(\a[22] ), .o1(new_n248));
  nand42aa1n16x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  aoib12aa1n02x5               g155(.a(new_n243), .b(new_n249), .c(new_n248), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n243), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n245), .o1(new_n253));
  aoai13aa1n02x5               g158(.a(new_n252), .b(new_n253), .c(new_n236), .d(new_n242), .o1(new_n254));
  aoi022aa1n03x5               g159(.a(new_n254), .b(new_n250), .c(new_n247), .d(new_n251), .o1(\s[22] ));
  inv000aa1n02x5               g160(.a(new_n235), .o1(new_n256));
  nano22aa1n02x5               g161(.a(new_n256), .b(new_n245), .c(new_n250), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n258));
  nano23aa1d15x5               g163(.a(new_n243), .b(new_n248), .c(new_n249), .d(new_n244), .out0(new_n259));
  aoi012aa1n09x5               g164(.a(new_n248), .b(new_n243), .c(new_n249), .o1(new_n260));
  inv020aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  aoi012aa1d18x5               g166(.a(new_n261), .b(new_n241), .c(new_n259), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(new_n258), .b(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  aoi112aa1n02x5               g169(.a(new_n264), .b(new_n261), .c(new_n241), .d(new_n259), .o1(new_n265));
  aoi022aa1n02x5               g170(.a(new_n263), .b(new_n264), .c(new_n258), .d(new_n265), .o1(\s[23] ));
  inv000aa1d42x5               g171(.a(new_n262), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n264), .b(new_n267), .c(new_n197), .d(new_n257), .o1(new_n268));
  tech160nm_fixorc02aa1n02p5x5 g173(.a(\a[24] ), .b(\b[23] ), .out0(new_n269));
  nor042aa1n09x5               g174(.a(\b[22] ), .b(\a[23] ), .o1(new_n270));
  norp02aa1n02x5               g175(.a(new_n269), .b(new_n270), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n270), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n264), .o1(new_n273));
  aoai13aa1n03x5               g178(.a(new_n272), .b(new_n273), .c(new_n258), .d(new_n262), .o1(new_n274));
  aoi022aa1n03x5               g179(.a(new_n274), .b(new_n269), .c(new_n268), .d(new_n271), .o1(\s[24] ));
  and002aa1n12x5               g180(.a(new_n269), .b(new_n264), .o(new_n276));
  nano22aa1n02x5               g181(.a(new_n256), .b(new_n276), .c(new_n259), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n278));
  nano22aa1n02x4               g183(.a(new_n225), .b(new_n220), .c(new_n226), .out0(new_n279));
  oai012aa1n02x7               g184(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .o1(new_n280));
  oab012aa1n04x5               g185(.a(new_n280), .b(new_n238), .c(new_n211), .out0(new_n281));
  inv020aa1n02x5               g186(.a(new_n240), .o1(new_n282));
  aoai13aa1n04x5               g187(.a(new_n259), .b(new_n282), .c(new_n281), .d(new_n279), .o1(new_n283));
  inv000aa1n06x5               g188(.a(new_n276), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[24] ), .b(\b[23] ), .c(new_n272), .carry(new_n285));
  aoai13aa1n12x5               g190(.a(new_n285), .b(new_n284), .c(new_n283), .d(new_n260), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(new_n278), .b(new_n287), .o1(new_n288));
  xorc02aa1n12x5               g193(.a(\a[25] ), .b(\b[24] ), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n276), .b(new_n261), .c(new_n241), .d(new_n259), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n289), .o1(new_n291));
  and003aa1n02x5               g196(.a(new_n290), .b(new_n291), .c(new_n285), .o(new_n292));
  aoi022aa1n02x5               g197(.a(new_n288), .b(new_n289), .c(new_n278), .d(new_n292), .o1(\s[25] ));
  aoai13aa1n03x5               g198(.a(new_n289), .b(new_n286), .c(new_n197), .d(new_n277), .o1(new_n294));
  tech160nm_fixorc02aa1n02p5x5 g199(.a(\a[26] ), .b(\b[25] ), .out0(new_n295));
  nor042aa1n03x5               g200(.a(\b[24] ), .b(\a[25] ), .o1(new_n296));
  norp02aa1n02x5               g201(.a(new_n295), .b(new_n296), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n296), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n291), .c(new_n278), .d(new_n287), .o1(new_n299));
  aoi022aa1n03x5               g204(.a(new_n299), .b(new_n295), .c(new_n294), .d(new_n297), .o1(\s[26] ));
  and002aa1n12x5               g205(.a(new_n295), .b(new_n289), .o(new_n301));
  nano32aa1n03x7               g206(.a(new_n256), .b(new_n301), .c(new_n259), .d(new_n276), .out0(new_n302));
  aoai13aa1n06x5               g207(.a(new_n302), .b(new_n209), .c(new_n131), .d(new_n193), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[26] ), .b(\b[25] ), .c(new_n298), .carry(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  aoi012aa1d18x5               g210(.a(new_n305), .b(new_n286), .c(new_n301), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(new_n303), .b(new_n306), .o1(new_n307));
  xorc02aa1n12x5               g212(.a(\a[27] ), .b(\b[26] ), .out0(new_n308));
  aoi112aa1n02x5               g213(.a(new_n308), .b(new_n305), .c(new_n286), .d(new_n301), .o1(new_n309));
  aoi022aa1n02x5               g214(.a(new_n307), .b(new_n308), .c(new_n303), .d(new_n309), .o1(\s[27] ));
  inv000aa1d42x5               g215(.a(new_n301), .o1(new_n311));
  aoai13aa1n04x5               g216(.a(new_n304), .b(new_n311), .c(new_n290), .d(new_n285), .o1(new_n312));
  aoai13aa1n02x5               g217(.a(new_n308), .b(new_n312), .c(new_n197), .d(new_n302), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[28] ), .b(\b[27] ), .out0(new_n314));
  norp02aa1n02x5               g219(.a(\b[26] ), .b(\a[27] ), .o1(new_n315));
  norp02aa1n02x5               g220(.a(new_n314), .b(new_n315), .o1(new_n316));
  inv000aa1n03x5               g221(.a(new_n315), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n308), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n317), .b(new_n318), .c(new_n303), .d(new_n306), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n319), .b(new_n314), .c(new_n313), .d(new_n316), .o1(\s[28] ));
  and002aa1n02x5               g225(.a(new_n314), .b(new_n308), .o(new_n321));
  aoai13aa1n02x5               g226(.a(new_n321), .b(new_n312), .c(new_n197), .d(new_n302), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .out0(new_n323));
  oao003aa1n02x5               g228(.a(\a[28] ), .b(\b[27] ), .c(new_n317), .carry(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(new_n325));
  inv000aa1d42x5               g230(.a(new_n321), .o1(new_n326));
  aoai13aa1n03x5               g231(.a(new_n324), .b(new_n326), .c(new_n303), .d(new_n306), .o1(new_n327));
  aoi022aa1n03x5               g232(.a(new_n327), .b(new_n323), .c(new_n322), .d(new_n325), .o1(\s[29] ));
  xorb03aa1n02x5               g233(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g234(.a(new_n318), .b(new_n314), .c(new_n323), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n312), .c(new_n197), .d(new_n302), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .out0(new_n332));
  oao003aa1n02x5               g237(.a(\a[29] ), .b(\b[28] ), .c(new_n324), .carry(new_n333));
  norb02aa1n02x5               g238(.a(new_n333), .b(new_n332), .out0(new_n334));
  inv000aa1d42x5               g239(.a(new_n330), .o1(new_n335));
  aoai13aa1n03x5               g240(.a(new_n333), .b(new_n335), .c(new_n303), .d(new_n306), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n336), .b(new_n332), .c(new_n331), .d(new_n334), .o1(\s[30] ));
  nano32aa1n06x5               g242(.a(new_n318), .b(new_n332), .c(new_n314), .d(new_n323), .out0(new_n338));
  aoai13aa1n02x5               g243(.a(new_n338), .b(new_n312), .c(new_n197), .d(new_n302), .o1(new_n339));
  xorc02aa1n02x5               g244(.a(\a[31] ), .b(\b[30] ), .out0(new_n340));
  and002aa1n02x5               g245(.a(\b[29] ), .b(\a[30] ), .o(new_n341));
  oabi12aa1n02x5               g246(.a(new_n340), .b(\a[30] ), .c(\b[29] ), .out0(new_n342));
  oab012aa1n02x4               g247(.a(new_n342), .b(new_n333), .c(new_n341), .out0(new_n343));
  inv000aa1d42x5               g248(.a(new_n338), .o1(new_n344));
  oao003aa1n02x5               g249(.a(\a[30] ), .b(\b[29] ), .c(new_n333), .carry(new_n345));
  aoai13aa1n03x5               g250(.a(new_n345), .b(new_n344), .c(new_n303), .d(new_n306), .o1(new_n346));
  aoi022aa1n03x5               g251(.a(new_n346), .b(new_n340), .c(new_n339), .d(new_n343), .o1(\s[31] ));
  oai012aa1n02x5               g252(.a(new_n102), .b(new_n107), .c(new_n106), .o1(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n348), .b(new_n111), .c(new_n104), .out0(\s[3] ));
  oaoi03aa1n02x5               g254(.a(\a[3] ), .b(\b[2] ), .c(new_n348), .o1(new_n350));
  xorb03aa1n02x5               g255(.a(new_n350), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xnbna2aa1n03x5               g256(.a(new_n135), .b(new_n110), .c(new_n112), .out0(\s[5] ));
  orn002aa1n02x5               g257(.a(\a[5] ), .b(\b[4] ), .o(new_n353));
  aoai13aa1n06x5               g258(.a(new_n353), .b(new_n116), .c(new_n110), .d(new_n112), .o1(new_n354));
  xorb03aa1n02x5               g259(.a(new_n354), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g260(.a(new_n115), .b(new_n118), .c(new_n354), .d(new_n117), .o1(new_n356));
  aoi112aa1n02x5               g261(.a(new_n118), .b(new_n115), .c(new_n354), .d(new_n117), .o1(new_n357));
  norb02aa1n02x5               g262(.a(new_n356), .b(new_n357), .out0(\s[7] ));
  xnbna2aa1n03x5               g263(.a(new_n120), .b(new_n356), .c(new_n125), .out0(\s[8] ));
  xorb03aa1n02x5               g264(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


