// Benchmark "adder" written by ABC on Wed Jul 17 21:42:52 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n310,
    new_n313, new_n314, new_n316, new_n317, new_n318, new_n319, new_n321,
    new_n322, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor042aa1n03x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor042aa1d18x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nor042aa1n06x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n106));
  xnrc02aa1n02x5               g011(.a(\b[5] ), .b(\a[6] ), .out0(new_n107));
  xnrc02aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .out0(new_n108));
  nor043aa1n03x5               g013(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n109));
  nor002aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nor022aa1n08x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nona23aa1n03x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  nanp02aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nand02aa1n02x5               g020(.a(\b[0] ), .b(\a[1] ), .o1(new_n116));
  nor002aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  tech160nm_fioai012aa1n04x5   g022(.a(new_n115), .b(new_n117), .c(new_n116), .o1(new_n118));
  oai012aa1n02x5               g023(.a(new_n111), .b(new_n112), .c(new_n110), .o1(new_n119));
  oai012aa1n06x5               g024(.a(new_n119), .b(new_n114), .c(new_n118), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n102), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n104), .b(new_n103), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[5] ), .o1(new_n123));
  oai022aa1n02x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  oaib12aa1n06x5               g029(.a(new_n124), .b(new_n123), .c(\a[6] ), .out0(new_n125));
  oai112aa1n06x5               g030(.a(new_n121), .b(new_n122), .c(new_n106), .d(new_n125), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n126), .c(new_n120), .d(new_n109), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n99), .b(new_n128), .c(new_n101), .out0(\s[10] ));
  aoi012aa1n12x5               g034(.a(new_n126), .b(new_n120), .c(new_n109), .o1(new_n130));
  inv000aa1d42x5               g035(.a(new_n127), .o1(new_n131));
  oai112aa1n04x5               g036(.a(new_n99), .b(new_n101), .c(new_n130), .d(new_n131), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1d06x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1d27x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nona22aa1n02x4               g041(.a(new_n132), .b(new_n136), .c(new_n98), .out0(new_n137));
  aoib12aa1n02x5               g042(.a(new_n135), .b(new_n132), .c(new_n98), .out0(new_n138));
  norb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(\s[11] ));
  inv030aa1n06x5               g044(.a(new_n133), .o1(new_n140));
  nor002aa1n06x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand02aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n06x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  xnbna2aa1n03x5               g048(.a(new_n143), .b(new_n137), .c(new_n140), .out0(\s[12] ));
  nona23aa1n09x5               g049(.a(new_n142), .b(new_n134), .c(new_n133), .d(new_n141), .out0(new_n145));
  oabi12aa1n18x5               g050(.a(new_n98), .b(new_n100), .c(new_n97), .out0(new_n146));
  tech160nm_fioaoi03aa1n05x5   g051(.a(\a[12] ), .b(\b[11] ), .c(new_n140), .o1(new_n147));
  oabi12aa1n18x5               g052(.a(new_n147), .b(new_n145), .c(new_n146), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nand23aa1n06x5               g054(.a(new_n99), .b(new_n135), .c(new_n143), .o1(new_n150));
  oai012aa1n03x5               g055(.a(new_n149), .b(new_n128), .c(new_n150), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n02x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n03x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n02x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand02aa1d04x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nano23aa1n06x5               g063(.a(new_n153), .b(new_n157), .c(new_n158), .d(new_n154), .out0(new_n159));
  nona23aa1n02x4               g064(.a(new_n159), .b(new_n127), .c(new_n130), .d(new_n150), .out0(new_n160));
  nano23aa1n03x7               g065(.a(new_n133), .b(new_n141), .c(new_n142), .d(new_n134), .out0(new_n161));
  oab012aa1n03x5               g066(.a(new_n98), .b(new_n97), .c(new_n100), .out0(new_n162));
  aoai13aa1n06x5               g067(.a(new_n159), .b(new_n147), .c(new_n161), .d(new_n162), .o1(new_n163));
  aoi012aa1n09x5               g068(.a(new_n157), .b(new_n153), .c(new_n158), .o1(new_n164));
  nand02aa1d06x5               g069(.a(new_n163), .b(new_n164), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  nor042aa1n06x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n03x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n160), .c(new_n166), .out0(\s[15] ));
  inv000aa1d42x5               g075(.a(new_n167), .o1(new_n171));
  nor043aa1n03x5               g076(.a(new_n130), .b(new_n131), .c(new_n150), .o1(new_n172));
  aoai13aa1n03x5               g077(.a(new_n169), .b(new_n165), .c(new_n172), .d(new_n159), .o1(new_n173));
  nor002aa1n03x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nand02aa1n03x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n173), .c(new_n171), .out0(\s[16] ));
  nona23aa1d18x5               g082(.a(new_n175), .b(new_n168), .c(new_n167), .d(new_n174), .out0(new_n178));
  nano23aa1n06x5               g083(.a(new_n150), .b(new_n178), .c(new_n159), .d(new_n127), .out0(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n126), .c(new_n109), .d(new_n120), .o1(new_n180));
  inv000aa1d42x5               g085(.a(new_n164), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n178), .o1(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n181), .c(new_n148), .d(new_n159), .o1(new_n183));
  tech160nm_fiaoi012aa1n03p5x5 g088(.a(new_n174), .b(new_n167), .c(new_n175), .o1(new_n184));
  nanp03aa1d12x5               g089(.a(new_n180), .b(new_n183), .c(new_n184), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g091(.a(\a[18] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[16] ), .o1(new_n189));
  tech160nm_fioaoi03aa1n03p5x5 g094(.a(new_n188), .b(new_n189), .c(new_n185), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(new_n187), .out0(\s[18] ));
  norb02aa1n09x5               g096(.a(new_n179), .b(new_n130), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n184), .b(new_n178), .c(new_n163), .d(new_n164), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n188), .b(\b[16] ), .c(new_n187), .d(\b[17] ), .out0(new_n194));
  oai012aa1n02x5               g099(.a(new_n194), .b(new_n192), .c(new_n193), .o1(new_n195));
  oai022aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oaib12aa1n02x5               g101(.a(new_n196), .b(new_n187), .c(\b[17] ), .out0(new_n197));
  nor042aa1n12x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nanp02aa1n04x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g108(.a(new_n198), .o1(new_n204));
  nanp02aa1n02x5               g109(.a(new_n189), .b(new_n188), .o1(new_n205));
  oaoi03aa1n02x5               g110(.a(\a[18] ), .b(\b[17] ), .c(new_n205), .o1(new_n206));
  aoai13aa1n06x5               g111(.a(new_n201), .b(new_n206), .c(new_n185), .d(new_n194), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1n08x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  nand03aa1n02x5               g115(.a(new_n207), .b(new_n204), .c(new_n210), .o1(new_n211));
  aoi012aa1n03x5               g116(.a(new_n210), .b(new_n207), .c(new_n204), .o1(new_n212));
  norb02aa1n02x7               g117(.a(new_n211), .b(new_n212), .out0(\s[20] ));
  nano23aa1n09x5               g118(.a(new_n198), .b(new_n208), .c(new_n209), .d(new_n199), .out0(new_n214));
  nand02aa1d04x5               g119(.a(new_n194), .b(new_n214), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  nona23aa1n09x5               g121(.a(new_n209), .b(new_n199), .c(new_n198), .d(new_n208), .out0(new_n217));
  aoi012aa1d18x5               g122(.a(new_n208), .b(new_n198), .c(new_n209), .o1(new_n218));
  oai012aa1n09x5               g123(.a(new_n218), .b(new_n217), .c(new_n197), .o1(new_n219));
  oaoi13aa1n06x5               g124(.a(new_n219), .b(new_n216), .c(new_n192), .d(new_n193), .o1(new_n220));
  nor042aa1n06x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  inv000aa1n09x5               g126(.a(new_n221), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n220), .b(new_n223), .c(new_n222), .out0(\s[21] ));
  norb02aa1n02x5               g129(.a(new_n223), .b(new_n221), .out0(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n219), .c(new_n185), .d(new_n216), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[21] ), .b(\a[22] ), .out0(new_n227));
  nand23aa1n03x5               g132(.a(new_n226), .b(new_n222), .c(new_n227), .o1(new_n228));
  aoi012aa1n03x5               g133(.a(new_n227), .b(new_n226), .c(new_n222), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n228), .b(new_n229), .out0(\s[22] ));
  nano22aa1n03x7               g135(.a(new_n227), .b(new_n222), .c(new_n223), .out0(new_n231));
  and003aa1n02x5               g136(.a(new_n194), .b(new_n231), .c(new_n214), .o(new_n232));
  oai012aa1n02x5               g137(.a(new_n232), .b(new_n192), .c(new_n193), .o1(new_n233));
  oao003aa1n02x5               g138(.a(\a[22] ), .b(\b[21] ), .c(new_n222), .carry(new_n234));
  inv000aa1n02x5               g139(.a(new_n234), .o1(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(new_n219), .c(new_n231), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[22] ), .b(\a[23] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  xnbna2aa1n03x5               g143(.a(new_n238), .b(new_n233), .c(new_n236), .out0(\s[23] ));
  nor042aa1n03x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n236), .o1(new_n242));
  aoai13aa1n04x5               g147(.a(new_n238), .b(new_n242), .c(new_n185), .d(new_n232), .o1(new_n243));
  xnrc02aa1n02x5               g148(.a(\b[23] ), .b(\a[24] ), .out0(new_n244));
  nanp03aa1n03x5               g149(.a(new_n243), .b(new_n241), .c(new_n244), .o1(new_n245));
  aoi012aa1n02x7               g150(.a(new_n244), .b(new_n243), .c(new_n241), .o1(new_n246));
  norb02aa1n02x7               g151(.a(new_n245), .b(new_n246), .out0(\s[24] ));
  nor042aa1n02x5               g152(.a(new_n244), .b(new_n237), .o1(new_n248));
  nano22aa1n06x5               g153(.a(new_n215), .b(new_n231), .c(new_n248), .out0(new_n249));
  inv000aa1n02x5               g154(.a(new_n218), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n231), .b(new_n250), .c(new_n214), .d(new_n206), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n248), .o1(new_n252));
  oao003aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .c(new_n241), .carry(new_n253));
  aoai13aa1n04x5               g158(.a(new_n253), .b(new_n252), .c(new_n251), .d(new_n234), .o1(new_n254));
  oaoi13aa1n04x5               g159(.a(new_n254), .b(new_n249), .c(new_n192), .d(new_n193), .o1(new_n255));
  xnrc02aa1n12x5               g160(.a(\b[24] ), .b(\a[25] ), .out0(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  xnrc02aa1n03x5               g162(.a(new_n255), .b(new_n257), .out0(\s[25] ));
  nor042aa1n03x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n257), .b(new_n254), .c(new_n185), .d(new_n249), .o1(new_n261));
  tech160nm_fixnrc02aa1n04x5   g166(.a(\b[25] ), .b(\a[26] ), .out0(new_n262));
  nand23aa1n03x5               g167(.a(new_n261), .b(new_n260), .c(new_n262), .o1(new_n263));
  aoi012aa1n03x5               g168(.a(new_n262), .b(new_n261), .c(new_n260), .o1(new_n264));
  norb02aa1n03x4               g169(.a(new_n263), .b(new_n264), .out0(\s[26] ));
  nor042aa1n04x5               g170(.a(new_n262), .b(new_n256), .o1(new_n266));
  nano32aa1n03x7               g171(.a(new_n215), .b(new_n266), .c(new_n231), .d(new_n248), .out0(new_n267));
  tech160nm_fioai012aa1n05x5   g172(.a(new_n267), .b(new_n192), .c(new_n193), .o1(new_n268));
  oao003aa1n02x5               g173(.a(\a[26] ), .b(\b[25] ), .c(new_n260), .carry(new_n269));
  aobi12aa1n06x5               g174(.a(new_n269), .b(new_n254), .c(new_n266), .out0(new_n270));
  xorc02aa1n02x5               g175(.a(\a[27] ), .b(\b[26] ), .out0(new_n271));
  xnbna2aa1n03x5               g176(.a(new_n271), .b(new_n268), .c(new_n270), .out0(\s[27] ));
  norp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  inv040aa1n03x5               g178(.a(new_n273), .o1(new_n274));
  aobi12aa1n03x5               g179(.a(new_n271), .b(new_n268), .c(new_n270), .out0(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[27] ), .b(\a[28] ), .out0(new_n276));
  nano22aa1n03x5               g181(.a(new_n275), .b(new_n274), .c(new_n276), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n248), .b(new_n235), .c(new_n219), .d(new_n231), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n266), .o1(new_n279));
  aoai13aa1n04x5               g184(.a(new_n269), .b(new_n279), .c(new_n278), .d(new_n253), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n271), .b(new_n280), .c(new_n185), .d(new_n267), .o1(new_n281));
  aoi012aa1n03x5               g186(.a(new_n276), .b(new_n281), .c(new_n274), .o1(new_n282));
  norp02aa1n03x5               g187(.a(new_n282), .b(new_n277), .o1(\s[28] ));
  norb02aa1n02x5               g188(.a(new_n271), .b(new_n276), .out0(new_n284));
  aobi12aa1n03x5               g189(.a(new_n284), .b(new_n268), .c(new_n270), .out0(new_n285));
  oao003aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .c(new_n274), .carry(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[28] ), .b(\a[29] ), .out0(new_n287));
  nano22aa1n03x5               g192(.a(new_n285), .b(new_n286), .c(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n284), .b(new_n280), .c(new_n185), .d(new_n267), .o1(new_n289));
  aoi012aa1n03x5               g194(.a(new_n287), .b(new_n289), .c(new_n286), .o1(new_n290));
  norp02aa1n03x5               g195(.a(new_n290), .b(new_n288), .o1(\s[29] ));
  xorb03aa1n02x5               g196(.a(new_n116), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g197(.a(new_n271), .b(new_n287), .c(new_n276), .out0(new_n293));
  aobi12aa1n03x5               g198(.a(new_n293), .b(new_n268), .c(new_n270), .out0(new_n294));
  oao003aa1n02x5               g199(.a(\a[29] ), .b(\b[28] ), .c(new_n286), .carry(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[29] ), .b(\a[30] ), .out0(new_n296));
  nano22aa1n03x5               g201(.a(new_n294), .b(new_n295), .c(new_n296), .out0(new_n297));
  aoai13aa1n02x7               g202(.a(new_n293), .b(new_n280), .c(new_n185), .d(new_n267), .o1(new_n298));
  aoi012aa1n03x5               g203(.a(new_n296), .b(new_n298), .c(new_n295), .o1(new_n299));
  nor002aa1n02x5               g204(.a(new_n299), .b(new_n297), .o1(\s[30] ));
  norb02aa1n02x5               g205(.a(new_n293), .b(new_n296), .out0(new_n301));
  aobi12aa1n03x5               g206(.a(new_n301), .b(new_n268), .c(new_n270), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n295), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  nano22aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n304), .out0(new_n305));
  aoai13aa1n06x5               g210(.a(new_n301), .b(new_n280), .c(new_n185), .d(new_n267), .o1(new_n306));
  aoi012aa1n02x7               g211(.a(new_n304), .b(new_n306), .c(new_n303), .o1(new_n307));
  norp02aa1n03x5               g212(.a(new_n307), .b(new_n305), .o1(\s[31] ));
  xnrb03aa1n02x5               g213(.a(new_n118), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g214(.a(\a[3] ), .b(\b[2] ), .c(new_n118), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g216(.a(new_n120), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g217(.a(new_n108), .b(new_n120), .out0(new_n313));
  tech160nm_fioai012aa1n03p5x5 g218(.a(new_n313), .b(\b[4] ), .c(\a[5] ), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g220(.a(new_n104), .b(new_n105), .out0(new_n316));
  nanb02aa1n02x5               g221(.a(new_n107), .b(new_n314), .out0(new_n317));
  oaoi13aa1n06x5               g222(.a(new_n316), .b(new_n317), .c(\a[6] ), .d(\b[5] ), .o1(new_n318));
  oai112aa1n02x5               g223(.a(new_n317), .b(new_n316), .c(\b[5] ), .d(\a[6] ), .o1(new_n319));
  norb02aa1n02x5               g224(.a(new_n319), .b(new_n318), .out0(\s[7] ));
  nanb02aa1n02x5               g225(.a(new_n102), .b(new_n103), .out0(new_n321));
  oab012aa1n02x4               g226(.a(new_n321), .b(new_n318), .c(new_n104), .out0(new_n322));
  aoi112aa1n02x5               g227(.a(new_n318), .b(new_n104), .c(new_n121), .d(new_n103), .o1(new_n323));
  norp02aa1n02x5               g228(.a(new_n322), .b(new_n323), .o1(\s[8] ));
  xnrc02aa1n02x5               g229(.a(new_n130), .b(new_n127), .out0(\s[9] ));
endmodule


