// Benchmark "adder" written by ABC on Wed Jul 17 20:11:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n341, new_n344, new_n346, new_n347, new_n349;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nona23aa1n02x4               g008(.a(new_n102), .b(new_n101), .c(new_n103), .d(new_n100), .out0(new_n104));
  xnrc02aa1n02x5               g009(.a(\b[5] ), .b(\a[6] ), .out0(new_n105));
  xnrc02aa1n02x5               g010(.a(\b[4] ), .b(\a[5] ), .out0(new_n106));
  nor043aa1n03x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  and002aa1n06x5               g012(.a(\b[3] ), .b(\a[4] ), .o(new_n108));
  inv040aa1d32x5               g013(.a(\a[3] ), .o1(new_n109));
  inv040aa1n08x5               g014(.a(\b[2] ), .o1(new_n110));
  nand42aa1n02x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(new_n111), .b(new_n112), .o1(new_n113));
  nor042aa1n02x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  nand42aa1n08x5               g019(.a(\b[0] ), .b(\a[1] ), .o1(new_n115));
  nand02aa1n08x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  aoi012aa1n06x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  oa0022aa1n06x5               g022(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n118));
  oaoi13aa1n12x5               g023(.a(new_n108), .b(new_n118), .c(new_n117), .d(new_n113), .o1(new_n119));
  aoi112aa1n02x5               g024(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n120));
  norb02aa1n03x5               g025(.a(new_n101), .b(new_n100), .out0(new_n121));
  norb02aa1n06x4               g026(.a(new_n102), .b(new_n103), .out0(new_n122));
  norp02aa1n02x5               g027(.a(\b[5] ), .b(\a[6] ), .o1(new_n123));
  aoi112aa1n09x5               g028(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n124));
  oai112aa1n04x5               g029(.a(new_n122), .b(new_n121), .c(new_n124), .d(new_n123), .o1(new_n125));
  nona22aa1n06x5               g030(.a(new_n125), .b(new_n120), .c(new_n100), .out0(new_n126));
  xorc02aa1n02x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n126), .c(new_n119), .d(new_n107), .o1(new_n128));
  norp02aa1n12x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1d28x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n128), .c(new_n99), .out0(\s[10] ));
  inv020aa1n04x5               g037(.a(new_n130), .o1(new_n133));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand22aa1n12x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv000aa1n02x5               g040(.a(new_n135), .o1(new_n136));
  oai112aa1n06x5               g041(.a(new_n128), .b(new_n99), .c(\b[9] ), .d(\a[10] ), .o1(new_n137));
  nona32aa1n02x4               g042(.a(new_n137), .b(new_n136), .c(new_n134), .d(new_n133), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n134), .o1(new_n139));
  aoi022aa1n02x5               g044(.a(new_n137), .b(new_n130), .c(new_n139), .d(new_n135), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n138), .b(new_n140), .out0(\s[11] ));
  nor002aa1d24x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand02aa1d12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  aoi113aa1n02x5               g049(.a(new_n134), .b(new_n144), .c(new_n137), .d(new_n135), .e(new_n130), .o1(new_n145));
  aobi12aa1n02x7               g050(.a(new_n144), .b(new_n138), .c(new_n139), .out0(new_n146));
  norp02aa1n02x5               g051(.a(new_n146), .b(new_n145), .o1(\s[12] ));
  and002aa1n02x7               g052(.a(\b[8] ), .b(\a[9] ), .o(new_n148));
  aoi112aa1n09x5               g053(.a(new_n133), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n149));
  norb03aa1d15x5               g054(.a(new_n143), .b(new_n134), .c(new_n142), .out0(new_n150));
  nona23aa1d16x5               g055(.a(new_n149), .b(new_n150), .c(new_n136), .d(new_n148), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n06x5               g057(.a(new_n152), .b(new_n126), .c(new_n119), .d(new_n107), .o1(new_n153));
  nona23aa1n09x5               g058(.a(new_n143), .b(new_n135), .c(new_n134), .d(new_n142), .out0(new_n154));
  oaih12aa1n12x5               g059(.a(new_n143), .b(new_n142), .c(new_n134), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n130), .b(new_n129), .c(new_n97), .d(new_n98), .o1(new_n156));
  oai012aa1d24x5               g061(.a(new_n155), .b(new_n154), .c(new_n156), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nor002aa1d32x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(new_n161));
  xobna2aa1n03x5               g066(.a(new_n161), .b(new_n153), .c(new_n158), .out0(\s[13] ));
  inv000aa1d42x5               g067(.a(new_n159), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n161), .c(new_n153), .d(new_n158), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n04x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  tech160nm_finand02aa1n03p5x5 g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  oai012aa1n02x7               g072(.a(new_n167), .b(new_n166), .c(new_n159), .o1(new_n168));
  nona23aa1n02x5               g073(.a(new_n167), .b(new_n160), .c(new_n159), .d(new_n166), .out0(new_n169));
  aoai13aa1n04x5               g074(.a(new_n168), .b(new_n169), .c(new_n153), .d(new_n158), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand42aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  nor002aa1d24x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  nanp02aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  aoi122aa1n02x5               g083(.a(new_n172), .b(new_n178), .c(new_n177), .d(new_n170), .e(new_n175), .o1(new_n179));
  inv000aa1d42x5               g084(.a(new_n172), .o1(new_n180));
  nanp02aa1n02x5               g085(.a(new_n170), .b(new_n175), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n176), .b(new_n178), .out0(new_n182));
  aoi012aa1n02x5               g087(.a(new_n182), .b(new_n181), .c(new_n180), .o1(new_n183));
  norp02aa1n03x5               g088(.a(new_n183), .b(new_n179), .o1(\s[16] ));
  nano23aa1n02x5               g089(.a(new_n159), .b(new_n166), .c(new_n167), .d(new_n160), .out0(new_n185));
  nano23aa1n03x7               g090(.a(new_n172), .b(new_n176), .c(new_n178), .d(new_n173), .out0(new_n186));
  nano22aa1d15x5               g091(.a(new_n151), .b(new_n185), .c(new_n186), .out0(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n126), .c(new_n119), .d(new_n107), .o1(new_n188));
  nona23aa1n03x5               g093(.a(new_n178), .b(new_n173), .c(new_n172), .d(new_n176), .out0(new_n189));
  nor042aa1n02x5               g094(.a(new_n189), .b(new_n169), .o1(new_n190));
  aoi112aa1n02x5               g095(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n191));
  oai012aa1n02x7               g096(.a(new_n177), .b(new_n189), .c(new_n168), .o1(new_n192));
  aoi112aa1n09x5               g097(.a(new_n192), .b(new_n191), .c(new_n157), .d(new_n190), .o1(new_n193));
  nand02aa1d08x5               g098(.a(new_n188), .b(new_n193), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g100(.a(\a[17] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[16] ), .o1(new_n197));
  oaoi03aa1n03x5               g102(.a(new_n196), .b(new_n197), .c(new_n194), .o1(new_n198));
  xnrb03aa1n03x5               g103(.a(new_n198), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n02x5               g104(.a(new_n197), .b(new_n196), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  nor022aa1n08x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nanp02aa1n06x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nanb02aa1n06x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  nano22aa1n09x5               g109(.a(new_n204), .b(new_n200), .c(new_n201), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  aoai13aa1n12x5               g111(.a(new_n203), .b(new_n202), .c(new_n196), .d(new_n197), .o1(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n206), .c(new_n188), .d(new_n193), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n09x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nor042aa1n02x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoi112aa1n02x5               g121(.a(new_n216), .b(new_n211), .c(new_n208), .d(new_n212), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n211), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n212), .b(new_n211), .out0(new_n219));
  nanp02aa1n03x5               g124(.a(new_n208), .b(new_n219), .o1(new_n220));
  tech160nm_fiaoi012aa1n02p5x5 g125(.a(new_n215), .b(new_n220), .c(new_n218), .o1(new_n221));
  norp02aa1n03x5               g126(.a(new_n221), .b(new_n217), .o1(\s[20] ));
  nano23aa1n06x5               g127(.a(new_n211), .b(new_n213), .c(new_n214), .d(new_n212), .out0(new_n223));
  nanp02aa1n02x5               g128(.a(new_n205), .b(new_n223), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n207), .o1(new_n225));
  oaih12aa1n02x5               g130(.a(new_n214), .b(new_n213), .c(new_n211), .o1(new_n226));
  aobi12aa1n06x5               g131(.a(new_n226), .b(new_n223), .c(new_n225), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n188), .d(new_n193), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  aoi112aa1n03x4               g137(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n233));
  inv000aa1n02x5               g138(.a(new_n230), .o1(new_n234));
  nanp02aa1n03x5               g139(.a(new_n228), .b(new_n231), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n232), .o1(new_n236));
  tech160nm_fiaoi012aa1n03p5x5 g141(.a(new_n236), .b(new_n235), .c(new_n234), .o1(new_n237));
  nor042aa1n03x5               g142(.a(new_n237), .b(new_n233), .o1(\s[22] ));
  inv000aa1d42x5               g143(.a(\a[21] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(\a[22] ), .o1(new_n240));
  xroi22aa1d04x5               g145(.a(new_n239), .b(\b[20] ), .c(new_n240), .d(\b[21] ), .out0(new_n241));
  nand23aa1n03x5               g146(.a(new_n241), .b(new_n205), .c(new_n223), .o1(new_n242));
  nona23aa1n02x4               g147(.a(new_n214), .b(new_n212), .c(new_n211), .d(new_n213), .out0(new_n243));
  oai012aa1n06x5               g148(.a(new_n226), .b(new_n243), .c(new_n207), .o1(new_n244));
  tech160nm_fioaoi03aa1n03p5x5 g149(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .o1(new_n245));
  aoi012aa1n02x5               g150(.a(new_n245), .b(new_n244), .c(new_n241), .o1(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n242), .c(new_n188), .d(new_n193), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor022aa1n12x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  nanp02aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  nor042aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nand42aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  aoi112aa1n03x4               g158(.a(new_n249), .b(new_n253), .c(new_n247), .d(new_n250), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n249), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n250), .b(new_n249), .out0(new_n256));
  nanp02aa1n03x5               g161(.a(new_n247), .b(new_n256), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n253), .o1(new_n258));
  tech160nm_fiaoi012aa1n03p5x5 g163(.a(new_n258), .b(new_n257), .c(new_n255), .o1(new_n259));
  nor042aa1n03x5               g164(.a(new_n259), .b(new_n254), .o1(\s[24] ));
  nano23aa1n06x5               g165(.a(new_n249), .b(new_n251), .c(new_n252), .d(new_n250), .out0(new_n261));
  nanb03aa1n02x5               g166(.a(new_n224), .b(new_n261), .c(new_n241), .out0(new_n262));
  nona22aa1n02x4               g167(.a(new_n252), .b(new_n251), .c(new_n249), .out0(new_n263));
  aoi022aa1n06x5               g168(.a(new_n261), .b(new_n245), .c(new_n263), .d(new_n252), .o1(new_n264));
  inv020aa1n03x5               g169(.a(new_n264), .o1(new_n265));
  aoi013aa1n03x5               g170(.a(new_n265), .b(new_n244), .c(new_n241), .d(new_n261), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n266), .b(new_n262), .c(new_n188), .d(new_n193), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  tech160nm_fixorc02aa1n02p5x5 g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xorc02aa1n12x5               g175(.a(\a[26] ), .b(\b[25] ), .out0(new_n271));
  aoi112aa1n03x4               g176(.a(new_n269), .b(new_n271), .c(new_n267), .d(new_n270), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n269), .o1(new_n273));
  nand02aa1n02x5               g178(.a(new_n267), .b(new_n270), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n271), .o1(new_n275));
  tech160nm_fiaoi012aa1n02p5x5 g180(.a(new_n275), .b(new_n274), .c(new_n273), .o1(new_n276));
  nor002aa1n02x5               g181(.a(new_n276), .b(new_n272), .o1(\s[26] ));
  nano23aa1n02x4               g182(.a(new_n103), .b(new_n100), .c(new_n101), .d(new_n102), .out0(new_n278));
  nona22aa1n02x4               g183(.a(new_n278), .b(new_n105), .c(new_n106), .out0(new_n279));
  inv000aa1d42x5               g184(.a(new_n108), .o1(new_n280));
  xorc02aa1n02x5               g185(.a(\a[3] ), .b(\b[2] ), .out0(new_n281));
  nanp02aa1n02x5               g186(.a(new_n116), .b(new_n115), .o1(new_n282));
  oai012aa1n02x5               g187(.a(new_n282), .b(\b[1] ), .c(\a[2] ), .o1(new_n283));
  inv000aa1n02x5               g188(.a(new_n118), .o1(new_n284));
  aoai13aa1n02x5               g189(.a(new_n280), .b(new_n284), .c(new_n283), .d(new_n281), .o1(new_n285));
  inv000aa1d42x5               g190(.a(\a[5] ), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\b[4] ), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(new_n287), .b(new_n286), .o1(new_n288));
  oaoi03aa1n02x5               g193(.a(\a[6] ), .b(\b[5] ), .c(new_n288), .o1(new_n289));
  aoi112aa1n02x5               g194(.a(new_n120), .b(new_n100), .c(new_n278), .d(new_n289), .o1(new_n290));
  oai012aa1n02x7               g195(.a(new_n290), .b(new_n285), .c(new_n279), .o1(new_n291));
  nanp02aa1n02x5               g196(.a(new_n157), .b(new_n190), .o1(new_n292));
  nona22aa1n02x4               g197(.a(new_n292), .b(new_n192), .c(new_n191), .out0(new_n293));
  and002aa1n12x5               g198(.a(new_n271), .b(new_n270), .o(new_n294));
  nano22aa1n03x7               g199(.a(new_n242), .b(new_n294), .c(new_n261), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n293), .c(new_n291), .d(new_n187), .o1(new_n296));
  nano22aa1n03x7               g201(.a(new_n227), .b(new_n241), .c(new_n261), .out0(new_n297));
  oaoi03aa1n02x5               g202(.a(\a[26] ), .b(\b[25] ), .c(new_n273), .o1(new_n298));
  oaoi13aa1n09x5               g203(.a(new_n298), .b(new_n294), .c(new_n297), .d(new_n265), .o1(new_n299));
  nor042aa1n06x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  nanp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  norb02aa1n02x5               g206(.a(new_n301), .b(new_n300), .out0(new_n302));
  xnbna2aa1n03x5               g207(.a(new_n302), .b(new_n296), .c(new_n299), .out0(\s[27] ));
  inv000aa1d42x5               g208(.a(new_n300), .o1(new_n304));
  aobi12aa1n02x7               g209(.a(new_n302), .b(new_n296), .c(new_n299), .out0(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[27] ), .b(\a[28] ), .out0(new_n306));
  nano22aa1n02x4               g211(.a(new_n305), .b(new_n304), .c(new_n306), .out0(new_n307));
  nanp03aa1n02x5               g212(.a(new_n244), .b(new_n241), .c(new_n261), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n294), .o1(new_n309));
  inv000aa1n02x5               g214(.a(new_n298), .o1(new_n310));
  aoai13aa1n06x5               g215(.a(new_n310), .b(new_n309), .c(new_n308), .d(new_n264), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n302), .b(new_n311), .c(new_n194), .d(new_n295), .o1(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n306), .b(new_n312), .c(new_n304), .o1(new_n313));
  norp02aa1n03x5               g218(.a(new_n313), .b(new_n307), .o1(\s[28] ));
  xnrc02aa1n02x5               g219(.a(\b[28] ), .b(\a[29] ), .out0(new_n315));
  nano22aa1n02x4               g220(.a(new_n306), .b(new_n304), .c(new_n301), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n311), .c(new_n194), .d(new_n295), .o1(new_n317));
  oao003aa1n03x5               g222(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n315), .b(new_n317), .c(new_n318), .o1(new_n319));
  aobi12aa1n02x7               g224(.a(new_n316), .b(new_n296), .c(new_n299), .out0(new_n320));
  nano22aa1n02x4               g225(.a(new_n320), .b(new_n315), .c(new_n318), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n115), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g228(.a(new_n315), .b(new_n306), .c(new_n301), .d(new_n304), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n311), .c(new_n194), .d(new_n295), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[29] ), .b(\b[28] ), .c(new_n318), .carry(new_n326));
  xnrc02aa1n02x5               g231(.a(\b[29] ), .b(\a[30] ), .out0(new_n327));
  tech160nm_fiaoi012aa1n02p5x5 g232(.a(new_n327), .b(new_n325), .c(new_n326), .o1(new_n328));
  aobi12aa1n02x7               g233(.a(new_n324), .b(new_n296), .c(new_n299), .out0(new_n329));
  nano22aa1n02x4               g234(.a(new_n329), .b(new_n326), .c(new_n327), .out0(new_n330));
  norp02aa1n03x5               g235(.a(new_n328), .b(new_n330), .o1(\s[30] ));
  xnrc02aa1n02x5               g236(.a(\b[30] ), .b(\a[31] ), .out0(new_n332));
  norb03aa1n02x5               g237(.a(new_n316), .b(new_n315), .c(new_n327), .out0(new_n333));
  aobi12aa1n02x7               g238(.a(new_n333), .b(new_n296), .c(new_n299), .out0(new_n334));
  oao003aa1n02x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n326), .carry(new_n335));
  nano22aa1n02x4               g240(.a(new_n334), .b(new_n332), .c(new_n335), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n333), .b(new_n311), .c(new_n194), .d(new_n295), .o1(new_n337));
  tech160nm_fiaoi012aa1n02p5x5 g242(.a(new_n332), .b(new_n337), .c(new_n335), .o1(new_n338));
  norp02aa1n03x5               g243(.a(new_n338), .b(new_n336), .o1(\s[31] ));
  xnbna2aa1n03x5               g244(.a(new_n117), .b(new_n111), .c(new_n112), .out0(\s[3] ));
  oaoi03aa1n02x5               g245(.a(\a[3] ), .b(\b[2] ), .c(new_n117), .o1(new_n341));
  xorb03aa1n02x5               g246(.a(new_n341), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g247(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g248(.a(new_n286), .b(new_n287), .c(new_n119), .o1(new_n344));
  xnrb03aa1n02x5               g249(.a(new_n344), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi112aa1n02x5               g250(.a(new_n285), .b(new_n106), .c(\a[6] ), .d(\b[5] ), .o1(new_n346));
  norp02aa1n02x5               g251(.a(new_n346), .b(new_n289), .o1(new_n347));
  xnrc02aa1n02x5               g252(.a(new_n347), .b(new_n122), .out0(\s[7] ));
  oaoi13aa1n02x5               g253(.a(new_n103), .b(new_n102), .c(new_n346), .d(new_n289), .o1(new_n349));
  xnrc02aa1n02x5               g254(.a(new_n349), .b(new_n121), .out0(\s[8] ));
  xorb03aa1n02x5               g255(.a(new_n291), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


