// Benchmark "adder" written by ABC on Wed Jul 17 13:55:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n339, new_n340, new_n341, new_n343, new_n344, new_n345, new_n347,
    new_n348, new_n349, new_n351, new_n353, new_n354, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  orn002aa1n06x5               g002(.a(\a[2] ), .b(\b[1] ), .o(new_n98));
  nanp02aa1n04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  aob012aa1n06x5               g004(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(new_n100));
  nor002aa1n20x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanb02aa1d24x5               g007(.a(new_n101), .b(new_n102), .out0(new_n103));
  oab012aa1d18x5               g008(.a(new_n101), .b(\a[4] ), .c(\b[3] ), .out0(new_n104));
  aoai13aa1n06x5               g009(.a(new_n104), .b(new_n103), .c(new_n100), .d(new_n98), .o1(new_n105));
  nanp02aa1n06x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  inv040aa1d32x5               g011(.a(\a[5] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[4] ), .o1(new_n108));
  nand02aa1d28x5               g013(.a(new_n108), .b(new_n107), .o1(new_n109));
  oai112aa1n03x5               g014(.a(new_n109), .b(new_n106), .c(\b[5] ), .d(\a[6] ), .o1(new_n110));
  nand02aa1n03x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  oai012aa1n02x5               g016(.a(new_n111), .b(\b[7] ), .c(\a[8] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  aoi022aa1d24x5               g018(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n114));
  oai112aa1n03x5               g019(.a(new_n114), .b(new_n113), .c(\b[6] ), .d(\a[7] ), .o1(new_n115));
  nor003aa1n03x5               g020(.a(new_n115), .b(new_n110), .c(new_n112), .o1(new_n116));
  oaih22aa1n06x5               g021(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  nor002aa1n03x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  and002aa1n02x7               g023(.a(\b[6] ), .b(\a[7] ), .o(new_n119));
  aoi112aa1n03x5               g024(.a(new_n119), .b(new_n118), .c(\a[6] ), .d(\b[5] ), .o1(new_n120));
  tech160nm_fixorc02aa1n05x5   g025(.a(\a[8] ), .b(\b[7] ), .out0(new_n121));
  nanp03aa1n02x5               g026(.a(new_n120), .b(new_n121), .c(new_n117), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\a[7] ), .o1(new_n123));
  nanb02aa1n02x5               g028(.a(\b[6] ), .b(new_n123), .out0(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  nanb02aa1n02x5               g030(.a(new_n125), .b(new_n122), .out0(new_n126));
  xnrc02aa1n12x5               g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n126), .c(new_n105), .d(new_n116), .o1(new_n129));
  tech160nm_fixnrc02aa1n05x5   g034(.a(\b[9] ), .b(\a[10] ), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n129), .c(new_n97), .out0(\s[10] ));
  nanp02aa1n06x5               g037(.a(new_n116), .b(new_n105), .o1(new_n133));
  aoi013aa1n09x5               g038(.a(new_n125), .b(new_n120), .c(new_n121), .d(new_n117), .o1(new_n134));
  aoai13aa1n02x5               g039(.a(new_n97), .b(new_n127), .c(new_n133), .d(new_n134), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(new_n135), .b(new_n131), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  oaih22aa1d12x5               g042(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n138), .b(new_n137), .o1(new_n139));
  inv040aa1d32x5               g044(.a(\a[11] ), .o1(new_n140));
  inv040aa1d28x5               g045(.a(\b[10] ), .o1(new_n141));
  nanp02aa1n04x5               g046(.a(new_n141), .b(new_n140), .o1(new_n142));
  nanp02aa1n04x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nanp02aa1n02x5               g048(.a(new_n142), .b(new_n143), .o1(new_n144));
  xobna2aa1n03x5               g049(.a(new_n144), .b(new_n136), .c(new_n139), .out0(\s[11] ));
  tech160nm_fiao0012aa1n02p5x5 g050(.a(new_n144), .b(new_n136), .c(new_n139), .o(new_n146));
  nor042aa1n12x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand22aa1n12x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n03x4               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  aboi22aa1n03x5               g054(.a(new_n147), .b(new_n148), .c(new_n140), .d(new_n141), .out0(new_n150));
  aoai13aa1n02x5               g055(.a(new_n142), .b(new_n144), .c(new_n136), .d(new_n139), .o1(new_n151));
  aoi022aa1n02x5               g056(.a(new_n146), .b(new_n150), .c(new_n151), .d(new_n149), .o1(\s[12] ));
  nona23aa1n09x5               g057(.a(new_n131), .b(new_n149), .c(new_n127), .d(new_n144), .out0(new_n153));
  nanb03aa1n12x5               g058(.a(new_n147), .b(new_n148), .c(new_n143), .out0(new_n154));
  nanp03aa1d12x5               g059(.a(new_n138), .b(new_n142), .c(new_n137), .o1(new_n155));
  nor002aa1n02x5               g060(.a(\b[10] ), .b(\a[11] ), .o1(new_n156));
  aoi012aa1n09x5               g061(.a(new_n147), .b(new_n156), .c(new_n148), .o1(new_n157));
  oai012aa1d24x5               g062(.a(new_n157), .b(new_n155), .c(new_n154), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n06x5               g064(.a(new_n159), .b(new_n153), .c(new_n133), .d(new_n134), .o1(new_n160));
  nor002aa1d32x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nanp02aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  norp02aa1n02x5               g068(.a(new_n158), .b(new_n163), .o1(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n153), .c(new_n133), .d(new_n134), .o1(new_n165));
  aobi12aa1n02x5               g070(.a(new_n165), .b(new_n163), .c(new_n160), .out0(\s[13] ));
  inv000aa1d42x5               g071(.a(new_n161), .o1(new_n167));
  nanp02aa1n02x5               g072(.a(new_n160), .b(new_n163), .o1(new_n168));
  norp02aa1n12x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nanp02aa1n06x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n168), .c(new_n167), .out0(\s[14] ));
  nona23aa1d18x5               g077(.a(new_n170), .b(new_n162), .c(new_n161), .d(new_n169), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  oaoi03aa1n02x5               g079(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n175));
  nor002aa1n03x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  aoai13aa1n03x5               g083(.a(new_n178), .b(new_n175), .c(new_n160), .d(new_n174), .o1(new_n179));
  aoi112aa1n02x5               g084(.a(new_n178), .b(new_n175), .c(new_n160), .d(new_n174), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(\s[15] ));
  nor042aa1n03x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand02aa1n03x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  norp02aa1n02x5               g089(.a(new_n184), .b(new_n176), .o1(new_n185));
  oaih12aa1n02x5               g090(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(new_n186), .b(new_n184), .c(new_n179), .d(new_n185), .o1(\s[16] ));
  aoi012aa1n02x5               g092(.a(new_n103), .b(new_n100), .c(new_n98), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n104), .o1(new_n189));
  norb02aa1n02x5               g094(.a(new_n106), .b(new_n117), .out0(new_n190));
  oai012aa1n02x5               g095(.a(new_n113), .b(\b[6] ), .c(\a[7] ), .o1(new_n191));
  nona23aa1n02x4               g096(.a(new_n190), .b(new_n114), .c(new_n191), .d(new_n112), .out0(new_n192));
  oab012aa1n06x5               g097(.a(new_n192), .b(new_n188), .c(new_n189), .out0(new_n193));
  nona23aa1n02x4               g098(.a(new_n183), .b(new_n177), .c(new_n176), .d(new_n182), .out0(new_n194));
  nor042aa1n06x5               g099(.a(new_n194), .b(new_n173), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n153), .out0(new_n196));
  tech160nm_fioai012aa1n03p5x5 g101(.a(new_n196), .b(new_n193), .c(new_n126), .o1(new_n197));
  nona23aa1n02x4               g102(.a(new_n148), .b(new_n143), .c(new_n156), .d(new_n147), .out0(new_n198));
  nona32aa1n03x5               g103(.a(new_n195), .b(new_n198), .c(new_n130), .d(new_n127), .out0(new_n199));
  nanb03aa1n02x5               g104(.a(new_n182), .b(new_n183), .c(new_n177), .out0(new_n200));
  oai122aa1n02x7               g105(.a(new_n170), .b(new_n169), .c(new_n161), .d(\b[14] ), .e(\a[15] ), .o1(new_n201));
  aoi012aa1n02x5               g106(.a(new_n182), .b(new_n176), .c(new_n183), .o1(new_n202));
  oai012aa1n02x5               g107(.a(new_n202), .b(new_n201), .c(new_n200), .o1(new_n203));
  aoi012aa1n12x5               g108(.a(new_n203), .b(new_n158), .c(new_n195), .o1(new_n204));
  aoai13aa1n12x5               g109(.a(new_n204), .b(new_n199), .c(new_n133), .d(new_n134), .o1(new_n205));
  xorc02aa1n02x5               g110(.a(\a[17] ), .b(\b[16] ), .out0(new_n206));
  aoi112aa1n02x5               g111(.a(new_n206), .b(new_n203), .c(new_n158), .d(new_n195), .o1(new_n207));
  aoi022aa1n02x5               g112(.a(new_n205), .b(new_n206), .c(new_n197), .d(new_n207), .o1(\s[17] ));
  inv040aa1d32x5               g113(.a(\a[17] ), .o1(new_n209));
  inv040aa1d32x5               g114(.a(\b[16] ), .o1(new_n210));
  nand42aa1n02x5               g115(.a(new_n210), .b(new_n209), .o1(new_n211));
  nanp02aa1n03x5               g116(.a(new_n205), .b(new_n206), .o1(new_n212));
  nor002aa1d32x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  nand42aa1d28x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n212), .c(new_n211), .out0(\s[18] ));
  nanp02aa1n02x5               g121(.a(\b[16] ), .b(\a[17] ), .o1(new_n217));
  nano32aa1n03x7               g122(.a(new_n213), .b(new_n211), .c(new_n214), .d(new_n217), .out0(new_n218));
  aoai13aa1n12x5               g123(.a(new_n214), .b(new_n213), .c(new_n209), .d(new_n210), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  tech160nm_fixorc02aa1n04x5   g125(.a(\a[19] ), .b(\b[18] ), .out0(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n220), .c(new_n205), .d(new_n218), .o1(new_n222));
  aoi112aa1n02x5               g127(.a(new_n221), .b(new_n220), .c(new_n205), .d(new_n218), .o1(new_n223));
  norb02aa1n03x4               g128(.a(new_n222), .b(new_n223), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  xorc02aa1n02x5               g130(.a(\a[20] ), .b(\b[19] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(\a[19] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\b[18] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\a[20] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\b[19] ), .o1(new_n230));
  nanp02aa1n02x5               g135(.a(new_n230), .b(new_n229), .o1(new_n231));
  nanp02aa1n02x5               g136(.a(\b[19] ), .b(\a[20] ), .o1(new_n232));
  aoi022aa1n02x5               g137(.a(new_n231), .b(new_n232), .c(new_n228), .d(new_n227), .o1(new_n233));
  oaib12aa1n06x5               g138(.a(new_n222), .b(\b[18] ), .c(new_n227), .out0(new_n234));
  aoi022aa1n03x5               g139(.a(new_n234), .b(new_n226), .c(new_n222), .d(new_n233), .o1(\s[20] ));
  nand23aa1n04x5               g140(.a(new_n218), .b(new_n221), .c(new_n226), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nand02aa1d06x5               g142(.a(new_n205), .b(new_n237), .o1(new_n238));
  nor042aa1n02x5               g143(.a(\b[18] ), .b(\a[19] ), .o1(new_n239));
  oai112aa1n04x5               g144(.a(new_n231), .b(new_n232), .c(new_n228), .d(new_n227), .o1(new_n240));
  tech160nm_fioaoi03aa1n02p5x5 g145(.a(new_n229), .b(new_n230), .c(new_n239), .o1(new_n241));
  oai013aa1d12x5               g146(.a(new_n241), .b(new_n240), .c(new_n219), .d(new_n239), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[20] ), .b(\a[21] ), .out0(new_n244));
  xobna2aa1n03x5               g149(.a(new_n244), .b(new_n238), .c(new_n243), .out0(\s[21] ));
  tech160nm_fiao0012aa1n03p5x5 g150(.a(new_n244), .b(new_n238), .c(new_n243), .o(new_n246));
  tech160nm_fixorc02aa1n03p5x5 g151(.a(\a[22] ), .b(\b[21] ), .out0(new_n247));
  nor042aa1n09x5               g152(.a(\b[20] ), .b(\a[21] ), .o1(new_n248));
  norp02aa1n02x5               g153(.a(new_n247), .b(new_n248), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n248), .o1(new_n250));
  aoai13aa1n03x5               g155(.a(new_n250), .b(new_n244), .c(new_n238), .d(new_n243), .o1(new_n251));
  aoi022aa1n02x7               g156(.a(new_n246), .b(new_n249), .c(new_n251), .d(new_n247), .o1(\s[22] ));
  norb02aa1n06x4               g157(.a(new_n247), .b(new_n244), .out0(new_n253));
  nand22aa1n12x5               g158(.a(new_n242), .b(new_n253), .o1(new_n254));
  oao003aa1n12x5               g159(.a(\a[22] ), .b(\b[21] ), .c(new_n250), .carry(new_n255));
  nanp02aa1n24x5               g160(.a(new_n254), .b(new_n255), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  nand23aa1n03x5               g162(.a(new_n205), .b(new_n237), .c(new_n253), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n258), .c(new_n257), .out0(\s[23] ));
  aob012aa1n03x5               g165(.a(new_n259), .b(new_n258), .c(new_n257), .out0(new_n261));
  tech160nm_fixorc02aa1n03p5x5 g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  norp02aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  norp02aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  aoi013aa1n02x4               g169(.a(new_n256), .b(new_n205), .c(new_n237), .d(new_n253), .o1(new_n265));
  tech160nm_fioaoi03aa1n02p5x5 g170(.a(\a[23] ), .b(\b[22] ), .c(new_n265), .o1(new_n266));
  aoi022aa1n03x5               g171(.a(new_n266), .b(new_n262), .c(new_n261), .d(new_n264), .o1(\s[24] ));
  nano32aa1n02x4               g172(.a(new_n244), .b(new_n262), .c(new_n247), .d(new_n259), .out0(new_n268));
  nand23aa1n06x5               g173(.a(new_n205), .b(new_n237), .c(new_n268), .o1(new_n269));
  and002aa1n06x5               g174(.a(new_n262), .b(new_n259), .o(new_n270));
  inv000aa1d42x5               g175(.a(\a[24] ), .o1(new_n271));
  inv000aa1d42x5               g176(.a(\b[23] ), .o1(new_n272));
  oaoi03aa1n12x5               g177(.a(new_n271), .b(new_n272), .c(new_n263), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  tech160nm_fiaoi012aa1n05x5   g179(.a(new_n274), .b(new_n256), .c(new_n270), .o1(new_n275));
  nanp02aa1n06x5               g180(.a(new_n269), .b(new_n275), .o1(new_n276));
  nor002aa1n16x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  and002aa1n03x5               g182(.a(\b[24] ), .b(\a[25] ), .o(new_n278));
  nor042aa1n02x5               g183(.a(new_n278), .b(new_n277), .o1(new_n279));
  aoi112aa1n02x5               g184(.a(new_n279), .b(new_n274), .c(new_n256), .d(new_n270), .o1(new_n280));
  aoi022aa1n02x5               g185(.a(new_n276), .b(new_n279), .c(new_n269), .d(new_n280), .o1(\s[25] ));
  nanp02aa1n03x5               g186(.a(new_n276), .b(new_n279), .o1(new_n282));
  xorc02aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .out0(new_n283));
  norp02aa1n02x5               g188(.a(new_n283), .b(new_n277), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n277), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n278), .c(new_n269), .d(new_n275), .o1(new_n286));
  aoi022aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n282), .d(new_n284), .o1(\s[26] ));
  and002aa1n06x5               g192(.a(new_n283), .b(new_n279), .o(new_n288));
  aoai13aa1n12x5               g193(.a(new_n288), .b(new_n274), .c(new_n256), .d(new_n270), .o1(new_n289));
  nano32aa1n02x5               g194(.a(new_n236), .b(new_n288), .c(new_n253), .d(new_n270), .out0(new_n290));
  oao003aa1n02x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n285), .carry(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  aoi012aa1n09x5               g197(.a(new_n292), .b(new_n205), .c(new_n290), .o1(new_n293));
  nand42aa1n02x5               g198(.a(new_n293), .b(new_n289), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoi112aa1n02x5               g200(.a(new_n295), .b(new_n292), .c(new_n205), .d(new_n290), .o1(new_n296));
  aoi022aa1n02x7               g201(.a(new_n294), .b(new_n295), .c(new_n289), .d(new_n296), .o1(\s[27] ));
  inv000aa1d42x5               g202(.a(new_n255), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n270), .b(new_n298), .c(new_n242), .d(new_n253), .o1(new_n299));
  aobi12aa1n06x5               g204(.a(new_n288), .b(new_n299), .c(new_n273), .out0(new_n300));
  nanb03aa1n03x5               g205(.a(new_n236), .b(new_n268), .c(new_n288), .out0(new_n301));
  aoai13aa1n04x5               g206(.a(new_n291), .b(new_n301), .c(new_n197), .d(new_n204), .o1(new_n302));
  oaih12aa1n02x5               g207(.a(new_n295), .b(new_n302), .c(new_n300), .o1(new_n303));
  xorc02aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .out0(new_n304));
  norp02aa1n02x5               g209(.a(\b[26] ), .b(\a[27] ), .o1(new_n305));
  norp02aa1n02x5               g210(.a(new_n304), .b(new_n305), .o1(new_n306));
  inv000aa1n03x5               g211(.a(new_n305), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n295), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n307), .b(new_n308), .c(new_n293), .d(new_n289), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n303), .d(new_n306), .o1(\s[28] ));
  and002aa1n02x5               g215(.a(new_n304), .b(new_n295), .o(new_n311));
  oaih12aa1n02x5               g216(.a(new_n311), .b(new_n302), .c(new_n300), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .out0(new_n313));
  oao003aa1n02x5               g218(.a(\a[28] ), .b(\b[27] ), .c(new_n307), .carry(new_n314));
  norb02aa1n02x5               g219(.a(new_n314), .b(new_n313), .out0(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  aoai13aa1n02x7               g221(.a(new_n314), .b(new_n316), .c(new_n293), .d(new_n289), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n312), .d(new_n315), .o1(\s[29] ));
  xorb03aa1n02x5               g223(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g224(.a(new_n308), .b(new_n304), .c(new_n313), .out0(new_n320));
  oaih12aa1n02x5               g225(.a(new_n320), .b(new_n302), .c(new_n300), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[29] ), .b(\b[28] ), .c(new_n314), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  inv000aa1n02x5               g229(.a(new_n320), .o1(new_n325));
  aoai13aa1n03x5               g230(.a(new_n323), .b(new_n325), .c(new_n293), .d(new_n289), .o1(new_n326));
  aoi022aa1n03x5               g231(.a(new_n326), .b(new_n322), .c(new_n321), .d(new_n324), .o1(\s[30] ));
  nano32aa1n02x4               g232(.a(new_n308), .b(new_n322), .c(new_n304), .d(new_n313), .out0(new_n328));
  oaih12aa1n02x5               g233(.a(new_n328), .b(new_n302), .c(new_n300), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  and002aa1n02x5               g235(.a(\b[29] ), .b(\a[30] ), .o(new_n331));
  oabi12aa1n02x5               g236(.a(new_n330), .b(\a[30] ), .c(\b[29] ), .out0(new_n332));
  oab012aa1n02x4               g237(.a(new_n332), .b(new_n323), .c(new_n331), .out0(new_n333));
  inv000aa1n02x5               g238(.a(new_n328), .o1(new_n334));
  oao003aa1n02x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n323), .carry(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n334), .c(new_n293), .d(new_n289), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n336), .b(new_n330), .c(new_n329), .d(new_n333), .o1(\s[31] ));
  xobna2aa1n03x5               g242(.a(new_n103), .b(new_n100), .c(new_n98), .out0(\s[3] ));
  xorc02aa1n02x5               g243(.a(\a[4] ), .b(\b[3] ), .out0(new_n339));
  norp03aa1n02x5               g244(.a(new_n188), .b(new_n339), .c(new_n101), .o1(new_n340));
  aboi22aa1n03x5               g245(.a(new_n188), .b(new_n104), .c(\a[4] ), .d(\b[3] ), .out0(new_n341));
  oaoi13aa1n02x5               g246(.a(new_n340), .b(new_n341), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  inv000aa1d42x5               g247(.a(new_n109), .o1(new_n343));
  nano32aa1n02x4               g248(.a(new_n343), .b(new_n105), .c(new_n111), .d(new_n106), .out0(new_n344));
  aoi022aa1n02x5               g249(.a(new_n105), .b(new_n111), .c(new_n106), .d(new_n109), .o1(new_n345));
  norp02aa1n02x5               g250(.a(new_n344), .b(new_n345), .o1(\s[5] ));
  xorc02aa1n02x5               g251(.a(\a[6] ), .b(\b[5] ), .out0(new_n347));
  oai012aa1n02x5               g252(.a(new_n347), .b(new_n344), .c(new_n343), .o1(new_n348));
  aoi113aa1n02x5               g253(.a(new_n347), .b(new_n343), .c(new_n105), .d(new_n111), .e(new_n106), .o1(new_n349));
  norb02aa1n02x5               g254(.a(new_n348), .b(new_n349), .out0(\s[6] ));
  oai012aa1n02x5               g255(.a(new_n348), .b(\b[5] ), .c(\a[6] ), .o1(new_n351));
  xorb03aa1n02x5               g256(.a(new_n351), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nona22aa1n02x4               g257(.a(new_n351), .b(new_n119), .c(new_n118), .out0(new_n353));
  nanp02aa1n02x5               g258(.a(new_n353), .b(new_n124), .o1(new_n354));
  norp02aa1n02x5               g259(.a(new_n121), .b(new_n118), .o1(new_n355));
  aoi022aa1n02x5               g260(.a(new_n354), .b(new_n121), .c(new_n353), .d(new_n355), .o1(\s[8] ));
  xnbna2aa1n03x5               g261(.a(new_n128), .b(new_n133), .c(new_n134), .out0(\s[9] ));
endmodule


