// Benchmark "adder" written by ABC on Thu Jul 18 00:31:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n179, new_n180, new_n181,
    new_n182, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n311, new_n314, new_n316, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d32x5               g001(.a(\a[4] ), .o1(new_n97));
  inv000aa1d48x5               g002(.a(\b[3] ), .o1(new_n98));
  tech160nm_finand02aa1n03p5x5 g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand42aa1n03x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(new_n99), .b(new_n100), .o1(new_n101));
  tech160nm_fixnrc02aa1n02p5x5 g006(.a(\b[2] ), .b(\a[3] ), .out0(new_n102));
  nand42aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nand22aa1n12x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  nor042aa1n06x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  oaih12aa1n06x5               g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  aoi112aa1n02x5               g011(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n107));
  norb02aa1n02x7               g012(.a(new_n99), .b(new_n107), .out0(new_n108));
  oai013aa1n06x5               g013(.a(new_n108), .b(new_n102), .c(new_n106), .d(new_n101), .o1(new_n109));
  nor022aa1n04x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand22aa1n09x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor022aa1n08x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n09x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .out0(new_n115));
  nor042aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nanb02aa1n02x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  nor043aa1n02x5               g023(.a(new_n114), .b(new_n115), .c(new_n118), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[6] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[5] ), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(new_n120), .b(new_n121), .c(new_n116), .o1(new_n122));
  tech160nm_fiao0012aa1n02p5x5 g027(.a(new_n110), .b(new_n112), .c(new_n111), .o(new_n123));
  oabi12aa1n06x5               g028(.a(new_n123), .b(new_n114), .c(new_n122), .out0(new_n124));
  aoi012aa1n02x5               g029(.a(new_n124), .b(new_n109), .c(new_n119), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[9] ), .b(\b[8] ), .c(new_n125), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand02aa1d08x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nor042aa1n04x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nano23aa1n03x7               g036(.a(new_n128), .b(new_n130), .c(new_n131), .d(new_n129), .out0(new_n132));
  aoai13aa1n03x5               g037(.a(new_n132), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n133));
  oai012aa1n12x5               g038(.a(new_n129), .b(new_n130), .c(new_n128), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(new_n133), .b(new_n134), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n16x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand22aa1n12x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  aoi012aa1n02x5               g043(.a(new_n137), .b(new_n135), .c(new_n138), .o1(new_n139));
  xnrb03aa1n02x5               g044(.a(new_n139), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1n16x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand22aa1n12x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nona23aa1n09x5               g047(.a(new_n142), .b(new_n138), .c(new_n137), .d(new_n141), .out0(new_n143));
  ao0012aa1n03x7               g048(.a(new_n141), .b(new_n137), .c(new_n142), .o(new_n144));
  oabi12aa1n18x5               g049(.a(new_n144), .b(new_n143), .c(new_n134), .out0(new_n145));
  oab012aa1n06x5               g050(.a(new_n145), .b(new_n133), .c(new_n143), .out0(new_n146));
  xnrb03aa1n02x5               g051(.a(new_n146), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n03x5               g052(.a(\a[13] ), .b(\b[12] ), .c(new_n146), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n20x5               g054(.a(\b[14] ), .b(\a[15] ), .o1(new_n150));
  nand42aa1d28x5               g055(.a(\b[14] ), .b(\a[15] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  nano23aa1d12x5               g057(.a(new_n137), .b(new_n141), .c(new_n142), .d(new_n138), .out0(new_n153));
  xnrc02aa1n12x5               g058(.a(\b[12] ), .b(\a[13] ), .out0(new_n154));
  xnrc02aa1n12x5               g059(.a(\b[13] ), .b(\a[14] ), .out0(new_n155));
  nor042aa1n06x5               g060(.a(new_n155), .b(new_n154), .o1(new_n156));
  nano32aa1n03x7               g061(.a(new_n125), .b(new_n156), .c(new_n132), .d(new_n153), .out0(new_n157));
  inv000aa1d42x5               g062(.a(\a[14] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(\b[13] ), .o1(new_n159));
  norp02aa1n02x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  oaoi03aa1n02x5               g065(.a(new_n158), .b(new_n159), .c(new_n160), .o1(new_n161));
  aobi12aa1n12x5               g066(.a(new_n161), .b(new_n145), .c(new_n156), .out0(new_n162));
  oaib12aa1n06x5               g067(.a(new_n152), .b(new_n157), .c(new_n162), .out0(new_n163));
  norb03aa1n02x5               g068(.a(new_n162), .b(new_n157), .c(new_n152), .out0(new_n164));
  norb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(\s[15] ));
  inv000aa1d42x5               g070(.a(new_n150), .o1(new_n166));
  nor042aa1n04x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nand42aa1n16x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n163), .c(new_n166), .out0(\s[16] ));
  nano23aa1d15x5               g075(.a(new_n150), .b(new_n167), .c(new_n168), .d(new_n151), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n167), .b(new_n150), .c(new_n168), .o1(new_n173));
  inv000aa1n02x5               g078(.a(new_n156), .o1(new_n174));
  nano32aa1n03x7               g079(.a(new_n174), .b(new_n171), .c(new_n132), .d(new_n153), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n176));
  oai112aa1n06x5               g081(.a(new_n176), .b(new_n173), .c(new_n162), .d(new_n172), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g083(.a(\a[18] ), .o1(new_n179));
  inv040aa1d32x5               g084(.a(\a[17] ), .o1(new_n180));
  inv030aa1d32x5               g085(.a(\b[16] ), .o1(new_n181));
  oaoi03aa1n03x5               g086(.a(new_n180), .b(new_n181), .c(new_n177), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[17] ), .c(new_n179), .out0(\s[18] ));
  nand42aa1n02x5               g088(.a(new_n109), .b(new_n119), .o1(new_n184));
  nanb02aa1n06x5               g089(.a(new_n124), .b(new_n184), .out0(new_n185));
  inv000aa1n06x5               g090(.a(new_n134), .o1(new_n186));
  aoai13aa1n02x7               g091(.a(new_n156), .b(new_n144), .c(new_n153), .d(new_n186), .o1(new_n187));
  aoai13aa1n06x5               g092(.a(new_n173), .b(new_n172), .c(new_n187), .d(new_n161), .o1(new_n188));
  xroi22aa1d06x4               g093(.a(new_n180), .b(\b[16] ), .c(new_n179), .d(\b[17] ), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n188), .c(new_n185), .d(new_n175), .o1(new_n190));
  oai022aa1n04x7               g095(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n191));
  oaib12aa1n12x5               g096(.a(new_n191), .b(new_n179), .c(\b[17] ), .out0(new_n192));
  nor002aa1d32x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nand42aa1d28x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(new_n193), .b(new_n194), .out0(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n190), .c(new_n192), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g103(.a(new_n193), .o1(new_n199));
  tech160nm_fiaoi012aa1n02p5x5 g104(.a(new_n195), .b(new_n190), .c(new_n192), .o1(new_n200));
  nor002aa1n16x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand02aa1d24x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nanb02aa1n02x5               g107(.a(new_n201), .b(new_n202), .out0(new_n203));
  nano22aa1n03x5               g108(.a(new_n200), .b(new_n199), .c(new_n203), .out0(new_n204));
  nanp02aa1n02x5               g109(.a(new_n181), .b(new_n180), .o1(new_n205));
  oaoi03aa1n12x5               g110(.a(\a[18] ), .b(\b[17] ), .c(new_n205), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n196), .b(new_n206), .c(new_n177), .d(new_n189), .o1(new_n207));
  aoi012aa1n03x5               g112(.a(new_n203), .b(new_n207), .c(new_n199), .o1(new_n208));
  nor002aa1n02x5               g113(.a(new_n208), .b(new_n204), .o1(\s[20] ));
  nano23aa1n06x5               g114(.a(new_n193), .b(new_n201), .c(new_n202), .d(new_n194), .out0(new_n210));
  nand02aa1d04x5               g115(.a(new_n189), .b(new_n210), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n03x5               g117(.a(new_n212), .b(new_n188), .c(new_n185), .d(new_n175), .o1(new_n213));
  nona23aa1n09x5               g118(.a(new_n202), .b(new_n194), .c(new_n193), .d(new_n201), .out0(new_n214));
  aoi012aa1n09x5               g119(.a(new_n201), .b(new_n193), .c(new_n202), .o1(new_n215));
  oai012aa1d24x5               g120(.a(new_n215), .b(new_n214), .c(new_n192), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  xorc02aa1n02x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  xnbna2aa1n03x5               g123(.a(new_n218), .b(new_n213), .c(new_n217), .out0(\s[21] ));
  orn002aa1n24x5               g124(.a(\a[21] ), .b(\b[20] ), .o(new_n220));
  aobi12aa1n02x5               g125(.a(new_n218), .b(new_n213), .c(new_n217), .out0(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[21] ), .b(\a[22] ), .out0(new_n222));
  nano22aa1n02x4               g127(.a(new_n221), .b(new_n220), .c(new_n222), .out0(new_n223));
  aoai13aa1n03x5               g128(.a(new_n218), .b(new_n216), .c(new_n177), .d(new_n212), .o1(new_n224));
  tech160nm_fiaoi012aa1n02p5x5 g129(.a(new_n222), .b(new_n224), .c(new_n220), .o1(new_n225));
  nor002aa1n02x5               g130(.a(new_n225), .b(new_n223), .o1(\s[22] ));
  nand42aa1n03x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  nano22aa1d18x5               g132(.a(new_n222), .b(new_n220), .c(new_n227), .out0(new_n228));
  oaoi03aa1n09x5               g133(.a(\a[22] ), .b(\b[21] ), .c(new_n220), .o1(new_n229));
  aoi012aa1d18x5               g134(.a(new_n229), .b(new_n216), .c(new_n228), .o1(new_n230));
  and003aa1n02x5               g135(.a(new_n189), .b(new_n228), .c(new_n210), .o(new_n231));
  aoai13aa1n03x5               g136(.a(new_n231), .b(new_n188), .c(new_n185), .d(new_n175), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[22] ), .b(\a[23] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnbna2aa1n03x5               g139(.a(new_n234), .b(new_n232), .c(new_n230), .out0(\s[23] ));
  nor042aa1n06x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi012aa1n02x7               g142(.a(new_n233), .b(new_n232), .c(new_n230), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[23] ), .b(\a[24] ), .out0(new_n239));
  nano22aa1n02x4               g144(.a(new_n238), .b(new_n237), .c(new_n239), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n230), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n234), .b(new_n241), .c(new_n177), .d(new_n231), .o1(new_n242));
  aoi012aa1n03x5               g147(.a(new_n239), .b(new_n242), .c(new_n237), .o1(new_n243));
  nor002aa1n02x5               g148(.a(new_n243), .b(new_n240), .o1(\s[24] ));
  nor042aa1n03x5               g149(.a(new_n239), .b(new_n233), .o1(new_n245));
  nano22aa1n06x5               g150(.a(new_n211), .b(new_n228), .c(new_n245), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n188), .c(new_n185), .d(new_n175), .o1(new_n247));
  inv040aa1n02x5               g152(.a(new_n215), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n228), .b(new_n248), .c(new_n210), .d(new_n206), .o1(new_n249));
  inv020aa1n02x5               g154(.a(new_n229), .o1(new_n250));
  inv020aa1n02x5               g155(.a(new_n245), .o1(new_n251));
  oao003aa1n02x5               g156(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .carry(new_n252));
  aoai13aa1n12x5               g157(.a(new_n252), .b(new_n251), .c(new_n249), .d(new_n250), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[24] ), .b(\a[25] ), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  xnbna2aa1n03x5               g161(.a(new_n256), .b(new_n247), .c(new_n254), .out0(\s[25] ));
  nor042aa1n03x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  aoi012aa1n02x5               g164(.a(new_n255), .b(new_n247), .c(new_n254), .o1(new_n260));
  tech160nm_fixnrc02aa1n04x5   g165(.a(\b[25] ), .b(\a[26] ), .out0(new_n261));
  nano22aa1n02x4               g166(.a(new_n260), .b(new_n259), .c(new_n261), .out0(new_n262));
  aoai13aa1n03x5               g167(.a(new_n256), .b(new_n253), .c(new_n177), .d(new_n246), .o1(new_n263));
  tech160nm_fiaoi012aa1n02p5x5 g168(.a(new_n261), .b(new_n263), .c(new_n259), .o1(new_n264));
  nor002aa1n02x5               g169(.a(new_n264), .b(new_n262), .o1(\s[26] ));
  nor042aa1n09x5               g170(.a(new_n261), .b(new_n255), .o1(new_n266));
  nano32aa1n03x7               g171(.a(new_n211), .b(new_n266), .c(new_n228), .d(new_n245), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n188), .c(new_n185), .d(new_n175), .o1(new_n268));
  oao003aa1n02x5               g173(.a(\a[26] ), .b(\b[25] ), .c(new_n259), .carry(new_n269));
  aobi12aa1n12x5               g174(.a(new_n269), .b(new_n253), .c(new_n266), .out0(new_n270));
  norp02aa1n02x5               g175(.a(\b[26] ), .b(\a[27] ), .o1(new_n271));
  nanp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  norb02aa1n02x5               g177(.a(new_n272), .b(new_n271), .out0(new_n273));
  xnbna2aa1n06x5               g178(.a(new_n273), .b(new_n268), .c(new_n270), .out0(\s[27] ));
  inv000aa1n06x5               g179(.a(new_n271), .o1(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[27] ), .b(\a[28] ), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n245), .b(new_n229), .c(new_n216), .d(new_n228), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n266), .o1(new_n278));
  aoai13aa1n04x5               g183(.a(new_n269), .b(new_n278), .c(new_n277), .d(new_n252), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n272), .b(new_n279), .c(new_n177), .d(new_n267), .o1(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n276), .b(new_n280), .c(new_n275), .o1(new_n281));
  aobi12aa1n06x5               g186(.a(new_n272), .b(new_n268), .c(new_n270), .out0(new_n282));
  nano22aa1n03x7               g187(.a(new_n282), .b(new_n275), .c(new_n276), .out0(new_n283));
  nor002aa1n02x5               g188(.a(new_n281), .b(new_n283), .o1(\s[28] ));
  nano22aa1n02x4               g189(.a(new_n276), .b(new_n275), .c(new_n272), .out0(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n279), .c(new_n177), .d(new_n267), .o1(new_n286));
  oao003aa1n02x5               g191(.a(\a[28] ), .b(\b[27] ), .c(new_n275), .carry(new_n287));
  xnrc02aa1n02x5               g192(.a(\b[28] ), .b(\a[29] ), .out0(new_n288));
  tech160nm_fiaoi012aa1n02p5x5 g193(.a(new_n288), .b(new_n286), .c(new_n287), .o1(new_n289));
  aobi12aa1n06x5               g194(.a(new_n285), .b(new_n268), .c(new_n270), .out0(new_n290));
  nano22aa1n03x7               g195(.a(new_n290), .b(new_n287), .c(new_n288), .out0(new_n291));
  norp02aa1n03x5               g196(.a(new_n289), .b(new_n291), .o1(\s[29] ));
  xorb03aa1n02x5               g197(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g198(.a(new_n273), .b(new_n288), .c(new_n276), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n279), .c(new_n177), .d(new_n267), .o1(new_n295));
  oao003aa1n02x5               g200(.a(\a[29] ), .b(\b[28] ), .c(new_n287), .carry(new_n296));
  xnrc02aa1n02x5               g201(.a(\b[29] ), .b(\a[30] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n295), .c(new_n296), .o1(new_n298));
  aobi12aa1n06x5               g203(.a(new_n294), .b(new_n268), .c(new_n270), .out0(new_n299));
  nano22aa1n03x7               g204(.a(new_n299), .b(new_n296), .c(new_n297), .out0(new_n300));
  norp02aa1n03x5               g205(.a(new_n298), .b(new_n300), .o1(\s[30] ));
  norb03aa1n02x5               g206(.a(new_n285), .b(new_n297), .c(new_n288), .out0(new_n302));
  aobi12aa1n06x5               g207(.a(new_n302), .b(new_n268), .c(new_n270), .out0(new_n303));
  oao003aa1n02x5               g208(.a(\a[30] ), .b(\b[29] ), .c(new_n296), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[30] ), .b(\a[31] ), .out0(new_n305));
  nano22aa1n03x7               g210(.a(new_n303), .b(new_n304), .c(new_n305), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n302), .b(new_n279), .c(new_n177), .d(new_n267), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n305), .b(new_n307), .c(new_n304), .o1(new_n308));
  norp02aa1n03x5               g213(.a(new_n308), .b(new_n306), .o1(\s[31] ));
  xnrb03aa1n02x5               g214(.a(new_n106), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g215(.a(\a[3] ), .b(\b[2] ), .c(new_n106), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g217(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g218(.a(new_n117), .b(new_n109), .c(new_n116), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[5] ), .c(new_n120), .out0(\s[6] ));
  oaoi03aa1n02x5               g220(.a(\a[6] ), .b(\b[5] ), .c(new_n314), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g222(.a(new_n112), .b(new_n316), .c(new_n113), .o1(new_n318));
  xnrb03aa1n02x5               g223(.a(new_n318), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g224(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


