// Benchmark "adder" written by ABC on Wed Jul 17 21:08:29 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n329, new_n331, new_n333, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  xnrc02aa1n02x5               g003(.a(\b[2] ), .b(\a[3] ), .out0(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n03x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor002aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai012aa1n02x5               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  norp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb03aa1n02x5               g011(.a(new_n106), .b(new_n104), .c(new_n105), .out0(new_n107));
  oai012aa1n06x5               g012(.a(new_n107), .b(new_n99), .c(new_n103), .o1(new_n108));
  norp02aa1n12x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(new_n109), .o1(new_n110));
  aoi022aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n111));
  norp02aa1n04x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nor002aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nona23aa1n02x4               g019(.a(new_n106), .b(new_n114), .c(new_n113), .d(new_n112), .out0(new_n115));
  nor002aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  aoi012aa1n02x5               g021(.a(new_n116), .b(\a[5] ), .c(\b[4] ), .o1(new_n117));
  nano32aa1n03x7               g022(.a(new_n115), .b(new_n117), .c(new_n110), .d(new_n111), .out0(new_n118));
  nanb02aa1n02x5               g023(.a(new_n113), .b(new_n114), .out0(new_n119));
  oa0012aa1n09x5               g024(.a(new_n114), .b(new_n116), .c(new_n113), .o(new_n120));
  inv000aa1n02x5               g025(.a(new_n120), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  norb03aa1n03x5               g027(.a(new_n122), .b(new_n109), .c(new_n112), .out0(new_n123));
  nanp02aa1n02x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nanb03aa1n02x5               g029(.a(new_n116), .b(new_n124), .c(new_n122), .out0(new_n125));
  oai013aa1n03x5               g030(.a(new_n121), .b(new_n123), .c(new_n125), .d(new_n119), .o1(new_n126));
  nanp02aa1n02x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n97), .out0(new_n128));
  aoai13aa1n03x5               g033(.a(new_n128), .b(new_n126), .c(new_n108), .d(new_n118), .o1(new_n129));
  norp02aa1n02x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n03x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  xorc02aa1n06x5               g038(.a(\a[11] ), .b(\b[10] ), .out0(new_n134));
  inv030aa1n02x5               g039(.a(new_n134), .o1(new_n135));
  nona22aa1n02x4               g040(.a(new_n129), .b(new_n130), .c(new_n97), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n135), .b(new_n136), .c(new_n131), .out0(\s[11] ));
  inv000aa1d42x5               g042(.a(\a[11] ), .o1(new_n138));
  inv000aa1d42x5               g043(.a(\b[10] ), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n139), .b(new_n138), .o1(new_n140));
  nanp03aa1n03x5               g045(.a(new_n136), .b(new_n131), .c(new_n134), .o1(new_n141));
  xorc02aa1n02x5               g046(.a(\a[12] ), .b(\b[11] ), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n141), .c(new_n140), .out0(\s[12] ));
  nano32aa1n02x4               g048(.a(new_n135), .b(new_n142), .c(new_n128), .d(new_n132), .out0(new_n144));
  aoai13aa1n03x5               g049(.a(new_n144), .b(new_n126), .c(new_n108), .d(new_n118), .o1(new_n145));
  nanp02aa1n02x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  oaih22aa1d12x5               g051(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n147));
  oai022aa1n02x5               g052(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n148));
  aoi022aa1n06x5               g053(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n146), .b(new_n147), .c(new_n148), .d(new_n149), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n145), .b(new_n150), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n02x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  aoi012aa1n02x5               g063(.a(new_n157), .b(new_n153), .c(new_n158), .o1(new_n159));
  nona23aa1n03x5               g064(.a(new_n158), .b(new_n154), .c(new_n153), .d(new_n157), .out0(new_n160));
  aoai13aa1n02x7               g065(.a(new_n159), .b(new_n160), .c(new_n145), .d(new_n150), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  xorc02aa1n03x5               g068(.a(\a[15] ), .b(\b[14] ), .out0(new_n164));
  tech160nm_fixorc02aa1n02p5x5 g069(.a(\a[16] ), .b(\b[15] ), .out0(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n163), .c(new_n161), .d(new_n164), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n165), .b(new_n163), .c(new_n161), .d(new_n164), .o1(new_n167));
  norb02aa1n03x4               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  nanp03aa1n02x5               g073(.a(new_n134), .b(new_n128), .c(new_n132), .o1(new_n169));
  nano23aa1n02x4               g074(.a(new_n153), .b(new_n157), .c(new_n158), .d(new_n154), .out0(new_n170));
  nand02aa1n03x5               g075(.a(new_n165), .b(new_n164), .o1(new_n171));
  nano23aa1n06x5               g076(.a(new_n169), .b(new_n171), .c(new_n170), .d(new_n142), .out0(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n126), .c(new_n108), .d(new_n118), .o1(new_n173));
  inv000aa1n02x5               g078(.a(new_n171), .o1(new_n174));
  oai012aa1n02x5               g079(.a(new_n159), .b(new_n150), .c(new_n160), .o1(new_n175));
  inv000aa1d42x5               g080(.a(\a[16] ), .o1(new_n176));
  inv000aa1d42x5               g081(.a(\b[15] ), .o1(new_n177));
  tech160nm_fioaoi03aa1n04x5   g082(.a(new_n176), .b(new_n177), .c(new_n163), .o1(new_n178));
  inv000aa1n02x5               g083(.a(new_n178), .o1(new_n179));
  aoi012aa1n12x5               g084(.a(new_n179), .b(new_n175), .c(new_n174), .o1(new_n180));
  xorc02aa1n12x5               g085(.a(\a[17] ), .b(\b[16] ), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n173), .c(new_n180), .out0(\s[17] ));
  nor022aa1n16x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n118), .b(new_n108), .o1(new_n185));
  norp03aa1n02x5               g090(.a(new_n123), .b(new_n125), .c(new_n119), .o1(new_n186));
  nona22aa1n02x4               g091(.a(new_n185), .b(new_n120), .c(new_n186), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n147), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n149), .b(new_n130), .c(new_n97), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n189), .b(new_n188), .o1(new_n190));
  nanp03aa1n02x5               g095(.a(new_n190), .b(new_n170), .c(new_n146), .o1(new_n191));
  aoai13aa1n02x5               g096(.a(new_n178), .b(new_n171), .c(new_n191), .d(new_n159), .o1(new_n192));
  aoai13aa1n02x5               g097(.a(new_n181), .b(new_n192), .c(new_n187), .d(new_n172), .o1(new_n193));
  xnrc02aa1n02x5               g098(.a(\b[17] ), .b(\a[18] ), .out0(new_n194));
  xobna2aa1n03x5               g099(.a(new_n194), .b(new_n193), .c(new_n184), .out0(\s[18] ));
  inv000aa1d42x5               g100(.a(\a[17] ), .o1(new_n196));
  inv020aa1n04x5               g101(.a(\a[18] ), .o1(new_n197));
  xroi22aa1d06x4               g102(.a(new_n196), .b(\b[16] ), .c(new_n197), .d(\b[17] ), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  oaoi03aa1n02x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n184), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n199), .c(new_n173), .d(new_n180), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand42aa1n02x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  xnrc02aa1n12x5               g111(.a(\b[19] ), .b(\a[20] ), .out0(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  aoi112aa1n02x5               g113(.a(new_n205), .b(new_n208), .c(new_n202), .d(new_n206), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n205), .o1(new_n210));
  aoi012aa1n06x5               g115(.a(new_n126), .b(new_n108), .c(new_n118), .o1(new_n211));
  nona22aa1n02x4               g116(.a(new_n144), .b(new_n160), .c(new_n171), .out0(new_n212));
  oai012aa1n12x5               g117(.a(new_n180), .b(new_n212), .c(new_n211), .o1(new_n213));
  nanb02aa1n09x5               g118(.a(new_n205), .b(new_n206), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n200), .c(new_n213), .d(new_n198), .o1(new_n216));
  aoi012aa1n03x5               g121(.a(new_n207), .b(new_n216), .c(new_n210), .o1(new_n217));
  norp02aa1n03x5               g122(.a(new_n217), .b(new_n209), .o1(\s[20] ));
  nona23aa1d18x5               g123(.a(new_n208), .b(new_n181), .c(new_n194), .d(new_n214), .out0(new_n219));
  oaih22aa1n06x5               g124(.a(\a[19] ), .b(\b[18] ), .c(\b[19] ), .d(\a[20] ), .o1(new_n220));
  nanp02aa1n02x5               g125(.a(\b[17] ), .b(\a[18] ), .o1(new_n221));
  oai022aa1n02x5               g126(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n222));
  nanp03aa1n02x5               g127(.a(new_n222), .b(new_n221), .c(new_n206), .o1(new_n223));
  aboi22aa1n03x5               g128(.a(new_n220), .b(new_n223), .c(\a[20] ), .d(\b[19] ), .out0(new_n224));
  inv000aa1n02x5               g129(.a(new_n224), .o1(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n219), .c(new_n173), .d(new_n180), .o1(new_n226));
  xorb03aa1n02x5               g131(.a(new_n226), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  nanb02aa1d36x5               g133(.a(\b[20] ), .b(new_n228), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoi112aa1n03x4               g138(.a(new_n230), .b(new_n233), .c(new_n226), .d(new_n231), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n219), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n231), .b(new_n224), .c(new_n213), .d(new_n235), .o1(new_n236));
  tech160nm_fiaoi012aa1n05x5   g141(.a(new_n232), .b(new_n236), .c(new_n229), .o1(new_n237));
  norp02aa1n02x5               g142(.a(new_n237), .b(new_n234), .o1(\s[22] ));
  nanp02aa1n02x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  nano22aa1n03x7               g144(.a(new_n232), .b(new_n229), .c(new_n239), .out0(new_n240));
  nona23aa1d18x5               g145(.a(new_n198), .b(new_n240), .c(new_n207), .d(new_n214), .out0(new_n241));
  oab012aa1n02x4               g146(.a(new_n183), .b(\a[18] ), .c(\b[17] ), .out0(new_n242));
  nano22aa1n03x7               g147(.a(new_n242), .b(new_n221), .c(new_n206), .out0(new_n243));
  nanp02aa1n02x5               g148(.a(\b[19] ), .b(\a[20] ), .o1(new_n244));
  nano32aa1n03x7               g149(.a(new_n232), .b(new_n239), .c(new_n229), .d(new_n244), .out0(new_n245));
  oaoi03aa1n02x5               g150(.a(\a[22] ), .b(\b[21] ), .c(new_n229), .o1(new_n246));
  oaoi13aa1n12x5               g151(.a(new_n246), .b(new_n245), .c(new_n243), .d(new_n220), .o1(new_n247));
  aoai13aa1n04x5               g152(.a(new_n247), .b(new_n241), .c(new_n173), .d(new_n180), .o1(new_n248));
  xorb03aa1n02x5               g153(.a(new_n248), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  xorc02aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .out0(new_n251));
  xorc02aa1n12x5               g156(.a(\a[24] ), .b(\b[23] ), .out0(new_n252));
  aoi112aa1n03x4               g157(.a(new_n250), .b(new_n252), .c(new_n248), .d(new_n251), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n250), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n241), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n247), .o1(new_n256));
  aoai13aa1n02x7               g161(.a(new_n251), .b(new_n256), .c(new_n213), .d(new_n255), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n252), .o1(new_n258));
  tech160nm_fiaoi012aa1n02p5x5 g163(.a(new_n258), .b(new_n257), .c(new_n254), .o1(new_n259));
  norp02aa1n02x5               g164(.a(new_n259), .b(new_n253), .o1(\s[24] ));
  nano32aa1n03x7               g165(.a(new_n219), .b(new_n252), .c(new_n240), .d(new_n251), .out0(new_n261));
  inv000aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  tech160nm_fioai012aa1n03p5x5 g167(.a(new_n245), .b(new_n243), .c(new_n220), .o1(new_n263));
  inv030aa1n02x5               g168(.a(new_n246), .o1(new_n264));
  nand22aa1n03x5               g169(.a(new_n252), .b(new_n251), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n254), .carry(new_n266));
  aoai13aa1n12x5               g171(.a(new_n266), .b(new_n265), .c(new_n263), .d(new_n264), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  aoai13aa1n04x5               g173(.a(new_n268), .b(new_n262), .c(new_n173), .d(new_n180), .o1(new_n269));
  xorb03aa1n02x5               g174(.a(new_n269), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  xorc02aa1n02x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xorc02aa1n12x5               g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  aoi112aa1n02x5               g178(.a(new_n271), .b(new_n273), .c(new_n269), .d(new_n272), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n271), .o1(new_n275));
  aoai13aa1n02x5               g180(.a(new_n272), .b(new_n267), .c(new_n213), .d(new_n261), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n273), .o1(new_n277));
  tech160nm_fiaoi012aa1n02p5x5 g182(.a(new_n277), .b(new_n276), .c(new_n275), .o1(new_n278));
  norp02aa1n02x5               g183(.a(new_n278), .b(new_n274), .o1(\s[26] ));
  inv000aa1n02x5               g184(.a(new_n265), .o1(new_n280));
  and002aa1n02x5               g185(.a(new_n273), .b(new_n272), .o(new_n281));
  nano22aa1n12x5               g186(.a(new_n241), .b(new_n280), .c(new_n281), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n192), .c(new_n187), .d(new_n172), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .c(new_n275), .carry(new_n284));
  aobi12aa1n09x5               g189(.a(new_n284), .b(new_n267), .c(new_n281), .out0(new_n285));
  xorc02aa1n02x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n285), .out0(\s[27] ));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv040aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  aobi12aa1n02x7               g194(.a(new_n286), .b(new_n283), .c(new_n285), .out0(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  nano22aa1n03x5               g196(.a(new_n290), .b(new_n289), .c(new_n291), .out0(new_n292));
  nanb02aa1n02x5               g197(.a(new_n220), .b(new_n223), .out0(new_n293));
  aoai13aa1n02x5               g198(.a(new_n280), .b(new_n246), .c(new_n293), .d(new_n245), .o1(new_n294));
  inv000aa1n02x5               g199(.a(new_n281), .o1(new_n295));
  aoai13aa1n02x5               g200(.a(new_n284), .b(new_n295), .c(new_n294), .d(new_n266), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n286), .b(new_n296), .c(new_n213), .d(new_n282), .o1(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n291), .b(new_n297), .c(new_n289), .o1(new_n298));
  norp02aa1n03x5               g203(.a(new_n298), .b(new_n292), .o1(\s[28] ));
  xnrc02aa1n02x5               g204(.a(\b[28] ), .b(\a[29] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n286), .b(new_n291), .out0(new_n301));
  aobi12aa1n02x7               g206(.a(new_n301), .b(new_n283), .c(new_n285), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n303));
  nano22aa1n03x5               g208(.a(new_n302), .b(new_n300), .c(new_n303), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n301), .b(new_n296), .c(new_n213), .d(new_n282), .o1(new_n305));
  tech160nm_fiaoi012aa1n02p5x5 g210(.a(new_n300), .b(new_n305), .c(new_n303), .o1(new_n306));
  norp02aa1n03x5               g211(.a(new_n306), .b(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g213(.a(new_n286), .b(new_n300), .c(new_n291), .out0(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n296), .c(new_n213), .d(new_n282), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .out0(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n312), .b(new_n310), .c(new_n311), .o1(new_n313));
  aobi12aa1n02x7               g218(.a(new_n309), .b(new_n283), .c(new_n285), .out0(new_n314));
  nano22aa1n03x5               g219(.a(new_n314), .b(new_n311), .c(new_n312), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n313), .b(new_n315), .o1(\s[30] ));
  norb02aa1n02x5               g221(.a(new_n309), .b(new_n312), .out0(new_n317));
  aobi12aa1n02x7               g222(.a(new_n317), .b(new_n283), .c(new_n285), .out0(new_n318));
  oao003aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n319));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n320), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n317), .b(new_n296), .c(new_n213), .d(new_n282), .o1(new_n322));
  tech160nm_fiaoi012aa1n02p5x5 g227(.a(new_n320), .b(new_n322), .c(new_n319), .o1(new_n323));
  norp02aa1n03x5               g228(.a(new_n323), .b(new_n321), .o1(\s[31] ));
  xnrb03aa1n02x5               g229(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanb02aa1n02x5               g230(.a(new_n105), .b(new_n106), .out0(new_n326));
  oaoi03aa1n02x5               g231(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n327));
  aob012aa1n02x5               g232(.a(new_n108), .b(new_n327), .c(new_n326), .out0(\s[4] ));
  xorc02aa1n02x5               g233(.a(\a[5] ), .b(\b[4] ), .out0(new_n329));
  xobna2aa1n03x5               g234(.a(new_n329), .b(new_n108), .c(new_n106), .out0(\s[5] ));
  aoi013aa1n02x4               g235(.a(new_n112), .b(new_n108), .c(new_n106), .d(new_n329), .o1(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n331), .b(new_n110), .c(new_n122), .out0(\s[6] ));
  oaoi03aa1n03x5               g237(.a(\a[6] ), .b(\b[5] ), .c(new_n331), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g239(.a(new_n116), .b(new_n333), .c(new_n124), .o1(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g241(.a(new_n211), .b(new_n127), .c(new_n98), .out0(\s[9] ));
endmodule


