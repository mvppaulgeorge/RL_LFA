// Benchmark "adder" written by ABC on Wed Jul 17 17:32:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n360, new_n362, new_n364, new_n365, new_n368, new_n370,
    new_n371, new_n372, new_n374;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n12x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n03x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand02aa1d20x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n04x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norb03aa1n12x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  xnrc02aa1n12x5               g007(.a(\b[3] ), .b(\a[4] ), .out0(new_n103));
  nand42aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nor042aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb03aa1n12x5               g010(.a(new_n105), .b(new_n100), .c(new_n104), .out0(new_n106));
  nor042aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  aob012aa1n03x5               g012(.a(new_n105), .b(\b[3] ), .c(\a[4] ), .out0(new_n108));
  norb02aa1n06x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  oai013aa1n06x5               g014(.a(new_n109), .b(new_n102), .c(new_n106), .d(new_n103), .o1(new_n110));
  nor002aa1d32x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand42aa1n06x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n06x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nona23aa1n02x4               g019(.a(new_n113), .b(new_n112), .c(new_n114), .d(new_n111), .out0(new_n115));
  tech160nm_fixorc02aa1n03p5x5 g020(.a(\a[7] ), .b(\b[6] ), .out0(new_n116));
  nor002aa1d32x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand42aa1n08x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanb02aa1d24x5               g023(.a(new_n117), .b(new_n118), .out0(new_n119));
  norb03aa1n03x5               g024(.a(new_n116), .b(new_n115), .c(new_n119), .out0(new_n120));
  nanp02aa1n04x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  oai112aa1n06x5               g026(.a(new_n118), .b(new_n121), .c(new_n117), .d(new_n111), .o1(new_n122));
  oab012aa1n03x5               g027(.a(new_n114), .b(\a[7] ), .c(\b[6] ), .out0(new_n123));
  aoi022aa1n09x5               g028(.a(new_n122), .b(new_n123), .c(\b[7] ), .d(\a[8] ), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n110), .d(new_n120), .o1(new_n126));
  nor042aa1n04x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nanp02aa1n09x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n06x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  inv000aa1n03x5               g035(.a(new_n102), .o1(new_n131));
  nona22aa1n12x5               g036(.a(new_n131), .b(new_n106), .c(new_n103), .out0(new_n132));
  norb02aa1n03x4               g037(.a(new_n112), .b(new_n111), .out0(new_n133));
  nanb02aa1n06x5               g038(.a(new_n114), .b(new_n113), .out0(new_n134));
  nona23aa1n06x5               g039(.a(new_n116), .b(new_n133), .c(new_n119), .d(new_n134), .out0(new_n135));
  inv040aa1n06x5               g040(.a(new_n124), .o1(new_n136));
  aoai13aa1n12x5               g041(.a(new_n136), .b(new_n135), .c(new_n132), .d(new_n109), .o1(new_n137));
  aoai13aa1n06x5               g042(.a(new_n129), .b(new_n97), .c(new_n137), .d(new_n125), .o1(new_n138));
  oai012aa1n02x5               g043(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n139));
  nand42aa1n08x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nor042aa1n06x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nanb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xobna2aa1n03x5               g047(.a(new_n142), .b(new_n138), .c(new_n139), .out0(\s[11] ));
  norb02aa1n02x5               g048(.a(new_n139), .b(new_n142), .out0(new_n144));
  nanp02aa1n03x5               g049(.a(new_n138), .b(new_n144), .o1(new_n145));
  orn002aa1n02x5               g050(.a(\a[12] ), .b(\b[11] ), .o(new_n146));
  nand02aa1d08x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  aoi022aa1n03x5               g052(.a(new_n145), .b(new_n140), .c(new_n147), .d(new_n146), .o1(new_n148));
  nor042aa1n04x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nano22aa1n02x4               g054(.a(new_n149), .b(new_n140), .c(new_n147), .out0(new_n150));
  aoi012aa1n02x7               g055(.a(new_n148), .b(new_n145), .c(new_n150), .o1(\s[12] ));
  nano23aa1n06x5               g056(.a(new_n149), .b(new_n141), .c(new_n147), .d(new_n140), .out0(new_n152));
  and003aa1n02x5               g057(.a(new_n152), .b(new_n129), .c(new_n125), .o(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n124), .c(new_n110), .d(new_n120), .o1(new_n154));
  norb03aa1n12x5               g059(.a(new_n147), .b(new_n141), .c(new_n149), .out0(new_n155));
  nand42aa1n02x5               g060(.a(new_n140), .b(new_n128), .o1(new_n156));
  oab012aa1n09x5               g061(.a(new_n156), .b(new_n97), .c(new_n127), .out0(new_n157));
  tech160nm_fiaoi012aa1n05x5   g062(.a(new_n149), .b(new_n141), .c(new_n147), .o1(new_n158));
  inv030aa1n04x5               g063(.a(new_n158), .o1(new_n159));
  aoi012aa1d24x5               g064(.a(new_n159), .b(new_n157), .c(new_n155), .o1(new_n160));
  nand22aa1n03x5               g065(.a(new_n154), .b(new_n160), .o1(new_n161));
  nand42aa1n04x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nor042aa1n06x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  aoi112aa1n02x5               g069(.a(new_n159), .b(new_n164), .c(new_n157), .d(new_n155), .o1(new_n165));
  aoi022aa1n02x5               g070(.a(new_n161), .b(new_n164), .c(new_n154), .d(new_n165), .o1(\s[13] ));
  inv000aa1n06x5               g071(.a(new_n163), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n160), .o1(new_n168));
  aoai13aa1n06x5               g073(.a(new_n164), .b(new_n168), .c(new_n137), .d(new_n153), .o1(new_n169));
  norp02aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand42aa1n06x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  nona23aa1n02x4               g077(.a(new_n169), .b(new_n171), .c(new_n170), .d(new_n163), .out0(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n172), .c(new_n167), .d(new_n169), .o1(\s[14] ));
  nano23aa1n06x5               g079(.a(new_n170), .b(new_n163), .c(new_n171), .d(new_n162), .out0(new_n175));
  tech160nm_fioaoi03aa1n04x5   g080(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n176));
  nand42aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nor002aa1n12x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n176), .c(new_n161), .d(new_n175), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n176), .c(new_n161), .d(new_n175), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(\s[15] ));
  inv000aa1d42x5               g087(.a(new_n178), .o1(new_n183));
  nor002aa1n04x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand02aa1n08x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  norb03aa1n02x5               g091(.a(new_n185), .b(new_n178), .c(new_n184), .out0(new_n187));
  tech160nm_finand02aa1n05x5   g092(.a(new_n180), .b(new_n187), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n186), .c(new_n183), .d(new_n180), .o1(\s[16] ));
  nor042aa1d18x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nand42aa1n04x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  norb02aa1n03x5               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  nano23aa1n06x5               g097(.a(new_n184), .b(new_n178), .c(new_n185), .d(new_n177), .out0(new_n193));
  nand02aa1d04x5               g098(.a(new_n193), .b(new_n175), .o1(new_n194));
  nano32aa1n09x5               g099(.a(new_n194), .b(new_n152), .c(new_n129), .d(new_n125), .out0(new_n195));
  aoai13aa1n06x5               g100(.a(new_n195), .b(new_n124), .c(new_n110), .d(new_n120), .o1(new_n196));
  oai112aa1n02x5               g101(.a(new_n146), .b(new_n147), .c(\b[10] ), .d(\a[11] ), .o1(new_n197));
  aoi022aa1n02x5               g102(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n198));
  oai012aa1n02x5               g103(.a(new_n198), .b(new_n127), .c(new_n97), .o1(new_n199));
  nona23aa1n02x4               g104(.a(new_n162), .b(new_n171), .c(new_n170), .d(new_n163), .out0(new_n200));
  oaoi13aa1n04x5               g105(.a(new_n200), .b(new_n158), .c(new_n197), .d(new_n199), .o1(new_n201));
  aoi012aa1d18x5               g106(.a(new_n184), .b(new_n178), .c(new_n185), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  oaoi13aa1n04x5               g108(.a(new_n203), .b(new_n193), .c(new_n201), .d(new_n176), .o1(new_n204));
  oai012aa1n02x5               g109(.a(new_n193), .b(new_n201), .c(new_n176), .o1(new_n205));
  oai022aa1n02x5               g110(.a(\a[16] ), .b(\b[15] ), .c(\b[16] ), .d(\a[17] ), .o1(new_n206));
  aoi122aa1n02x5               g111(.a(new_n206), .b(\b[16] ), .c(\a[17] ), .d(new_n178), .e(new_n185), .o1(new_n207));
  nanp03aa1n02x5               g112(.a(new_n196), .b(new_n205), .c(new_n207), .o1(new_n208));
  aoai13aa1n02x5               g113(.a(new_n208), .b(new_n192), .c(new_n204), .d(new_n196), .o1(\s[17] ));
  nor042aa1d18x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nand02aa1d28x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  nanb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  nanp02aa1n02x5               g117(.a(new_n208), .b(new_n191), .o1(new_n213));
  nano22aa1n02x4               g118(.a(new_n210), .b(new_n191), .c(new_n211), .out0(new_n214));
  aoi022aa1n02x5               g119(.a(new_n213), .b(new_n212), .c(new_n208), .d(new_n214), .o1(\s[18] ));
  inv000aa1n02x5               g120(.a(new_n176), .o1(new_n216));
  inv000aa1n02x5               g121(.a(new_n193), .o1(new_n217));
  aoai13aa1n12x5               g122(.a(new_n175), .b(new_n159), .c(new_n157), .d(new_n155), .o1(new_n218));
  aoai13aa1n12x5               g123(.a(new_n202), .b(new_n217), .c(new_n218), .d(new_n216), .o1(new_n219));
  nano23aa1n02x4               g124(.a(new_n190), .b(new_n210), .c(new_n211), .d(new_n191), .out0(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n219), .c(new_n137), .d(new_n195), .o1(new_n221));
  oa0012aa1n02x5               g126(.a(new_n211), .b(new_n210), .c(new_n190), .o(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  nand02aa1n12x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  nor002aa1d32x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  norb02aa1n12x5               g130(.a(new_n224), .b(new_n225), .out0(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n221), .c(new_n223), .out0(\s[19] ));
  xnrc02aa1n02x5               g132(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g133(.a(new_n225), .o1(new_n229));
  nand02aa1d06x5               g134(.a(new_n204), .b(new_n196), .o1(new_n230));
  aoai13aa1n03x5               g135(.a(new_n226), .b(new_n222), .c(new_n230), .d(new_n220), .o1(new_n231));
  nor002aa1n16x5               g136(.a(\b[19] ), .b(\a[20] ), .o1(new_n232));
  nand02aa1d28x5               g137(.a(\b[19] ), .b(\a[20] ), .o1(new_n233));
  norb02aa1n03x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  inv030aa1n03x5               g139(.a(new_n226), .o1(new_n235));
  norb03aa1n09x5               g140(.a(new_n233), .b(new_n225), .c(new_n232), .out0(new_n236));
  aoai13aa1n02x7               g141(.a(new_n236), .b(new_n235), .c(new_n221), .d(new_n223), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n234), .c(new_n231), .d(new_n229), .o1(\s[20] ));
  nano23aa1n09x5               g143(.a(new_n235), .b(new_n212), .c(new_n234), .d(new_n192), .out0(new_n239));
  aoai13aa1n03x5               g144(.a(new_n239), .b(new_n219), .c(new_n137), .d(new_n195), .o1(new_n240));
  nona22aa1n09x5               g145(.a(new_n233), .b(new_n232), .c(new_n225), .out0(new_n241));
  oai112aa1n06x5               g146(.a(new_n211), .b(new_n224), .c(new_n210), .d(new_n190), .o1(new_n242));
  aoi012aa1n12x5               g147(.a(new_n232), .b(new_n225), .c(new_n233), .o1(new_n243));
  oai012aa1n18x5               g148(.a(new_n243), .b(new_n242), .c(new_n241), .o1(new_n244));
  nand42aa1n04x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  nor042aa1d18x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  norb02aa1n03x5               g151(.a(new_n245), .b(new_n246), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n244), .c(new_n230), .d(new_n239), .o1(new_n248));
  nand22aa1n03x5               g153(.a(new_n224), .b(new_n211), .o1(new_n249));
  oab012aa1n03x5               g154(.a(new_n249), .b(new_n190), .c(new_n210), .out0(new_n250));
  inv000aa1n06x5               g155(.a(new_n243), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(new_n251), .b(new_n247), .c(new_n250), .d(new_n236), .o1(new_n252));
  aobi12aa1n03x7               g157(.a(new_n248), .b(new_n252), .c(new_n240), .out0(\s[21] ));
  inv000aa1d42x5               g158(.a(new_n246), .o1(new_n254));
  nor002aa1n12x5               g159(.a(\b[21] ), .b(\a[22] ), .o1(new_n255));
  nand42aa1n16x5               g160(.a(\b[21] ), .b(\a[22] ), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n244), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n247), .o1(new_n259));
  norb03aa1n02x5               g164(.a(new_n256), .b(new_n246), .c(new_n255), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n259), .c(new_n240), .d(new_n258), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n257), .c(new_n248), .d(new_n254), .o1(\s[22] ));
  inv000aa1n02x5               g167(.a(new_n239), .o1(new_n263));
  nano22aa1n02x4               g168(.a(new_n263), .b(new_n247), .c(new_n257), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n264), .b(new_n219), .c(new_n137), .d(new_n195), .o1(new_n265));
  nano23aa1d15x5               g170(.a(new_n255), .b(new_n246), .c(new_n256), .d(new_n245), .out0(new_n266));
  aoi012aa1d24x5               g171(.a(new_n255), .b(new_n246), .c(new_n256), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  aoi012aa1n02x5               g173(.a(new_n268), .b(new_n244), .c(new_n266), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(new_n265), .b(new_n269), .o1(new_n270));
  nor042aa1n02x5               g175(.a(\b[22] ), .b(\a[23] ), .o1(new_n271));
  and002aa1n12x5               g176(.a(\b[22] ), .b(\a[23] ), .o(new_n272));
  nor042aa1n06x5               g177(.a(new_n272), .b(new_n271), .o1(new_n273));
  aoi112aa1n02x5               g178(.a(new_n273), .b(new_n268), .c(new_n244), .d(new_n266), .o1(new_n274));
  aoi022aa1n02x5               g179(.a(new_n270), .b(new_n273), .c(new_n265), .d(new_n274), .o1(\s[23] ));
  aoai13aa1n06x5               g180(.a(new_n266), .b(new_n251), .c(new_n250), .d(new_n236), .o1(new_n276));
  aoi112aa1n02x5               g181(.a(new_n255), .b(new_n271), .c(new_n246), .d(new_n256), .o1(new_n277));
  nanp02aa1n03x5               g182(.a(new_n276), .b(new_n277), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[24] ), .b(\b[23] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n272), .c(new_n265), .d(new_n279), .o1(new_n281));
  orn002aa1n02x5               g186(.a(new_n280), .b(new_n272), .o(new_n282));
  aoai13aa1n03x5               g187(.a(new_n281), .b(new_n282), .c(new_n279), .d(new_n265), .o1(\s[24] ));
  nano32aa1n02x5               g188(.a(new_n263), .b(new_n280), .c(new_n266), .d(new_n273), .out0(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n219), .c(new_n137), .d(new_n195), .o1(new_n285));
  and002aa1n02x5               g190(.a(new_n280), .b(new_n273), .o(new_n286));
  inv000aa1n02x5               g191(.a(new_n286), .o1(new_n287));
  orn002aa1n02x5               g192(.a(\a[23] ), .b(\b[22] ), .o(new_n288));
  oao003aa1n02x5               g193(.a(\a[24] ), .b(\b[23] ), .c(new_n288), .carry(new_n289));
  aoai13aa1n12x5               g194(.a(new_n289), .b(new_n287), .c(new_n276), .d(new_n267), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[25] ), .b(\b[24] ), .out0(new_n291));
  aoai13aa1n06x5               g196(.a(new_n291), .b(new_n290), .c(new_n230), .d(new_n284), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n286), .b(new_n268), .c(new_n244), .d(new_n266), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n291), .o1(new_n294));
  and003aa1n02x5               g199(.a(new_n293), .b(new_n294), .c(new_n289), .o(new_n295));
  aobi12aa1n03x7               g200(.a(new_n292), .b(new_n295), .c(new_n285), .out0(\s[25] ));
  nor042aa1n03x5               g201(.a(\b[24] ), .b(\a[25] ), .o1(new_n297));
  inv000aa1n02x5               g202(.a(new_n297), .o1(new_n298));
  norp02aa1n02x5               g203(.a(\b[25] ), .b(\a[26] ), .o1(new_n299));
  and002aa1n03x5               g204(.a(\b[25] ), .b(\a[26] ), .o(new_n300));
  nor002aa1n02x5               g205(.a(new_n300), .b(new_n299), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n290), .o1(new_n302));
  norp03aa1n02x5               g207(.a(new_n300), .b(new_n299), .c(new_n297), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n294), .c(new_n285), .d(new_n302), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n292), .d(new_n298), .o1(\s[26] ));
  and002aa1n12x5               g210(.a(new_n291), .b(new_n301), .o(new_n306));
  nano32aa1n03x7               g211(.a(new_n263), .b(new_n306), .c(new_n266), .d(new_n286), .out0(new_n307));
  aoai13aa1n06x5               g212(.a(new_n307), .b(new_n219), .c(new_n137), .d(new_n195), .o1(new_n308));
  oab012aa1n02x4               g213(.a(new_n299), .b(new_n298), .c(new_n300), .out0(new_n309));
  inv000aa1n02x5               g214(.a(new_n309), .o1(new_n310));
  aoi012aa1n12x5               g215(.a(new_n310), .b(new_n290), .c(new_n306), .o1(new_n311));
  nanp02aa1n02x5               g216(.a(new_n308), .b(new_n311), .o1(new_n312));
  nor042aa1n04x5               g217(.a(\b[26] ), .b(\a[27] ), .o1(new_n313));
  and002aa1n12x5               g218(.a(\b[26] ), .b(\a[27] ), .o(new_n314));
  nor042aa1n03x5               g219(.a(new_n314), .b(new_n313), .o1(new_n315));
  aoi112aa1n02x5               g220(.a(new_n315), .b(new_n310), .c(new_n290), .d(new_n306), .o1(new_n316));
  aoi022aa1n02x5               g221(.a(new_n312), .b(new_n315), .c(new_n308), .d(new_n316), .o1(\s[27] ));
  inv000aa1d42x5               g222(.a(new_n306), .o1(new_n318));
  aoai13aa1n04x5               g223(.a(new_n309), .b(new_n318), .c(new_n293), .d(new_n289), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n314), .o1(new_n320));
  aoai13aa1n02x5               g225(.a(new_n320), .b(new_n319), .c(new_n230), .d(new_n307), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[28] ), .b(\b[27] ), .out0(new_n322));
  norp02aa1n02x5               g227(.a(new_n322), .b(new_n313), .o1(new_n323));
  inv000aa1d42x5               g228(.a(new_n313), .o1(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n314), .c(new_n308), .d(new_n311), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n325), .b(new_n322), .c(new_n321), .d(new_n323), .o1(\s[28] ));
  and002aa1n06x5               g231(.a(new_n322), .b(new_n315), .o(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n319), .c(new_n230), .d(new_n307), .o1(new_n328));
  inv020aa1n02x5               g233(.a(new_n327), .o1(new_n329));
  oao003aa1n02x5               g234(.a(\a[28] ), .b(\b[27] ), .c(new_n324), .carry(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n329), .c(new_n308), .d(new_n311), .o1(new_n331));
  xorc02aa1n02x5               g236(.a(\a[29] ), .b(\b[28] ), .out0(new_n332));
  norb02aa1n02x5               g237(.a(new_n330), .b(new_n332), .out0(new_n333));
  aoi022aa1n03x5               g238(.a(new_n331), .b(new_n332), .c(new_n328), .d(new_n333), .o1(\s[29] ));
  xorb03aa1n02x5               g239(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g240(.a(new_n322), .b(new_n332), .c(new_n315), .o(new_n336));
  aoai13aa1n02x5               g241(.a(new_n336), .b(new_n319), .c(new_n230), .d(new_n307), .o1(new_n337));
  inv000aa1d42x5               g242(.a(new_n336), .o1(new_n338));
  inv000aa1d42x5               g243(.a(\b[28] ), .o1(new_n339));
  inv000aa1d42x5               g244(.a(\a[29] ), .o1(new_n340));
  oaib12aa1n02x5               g245(.a(new_n330), .b(\b[28] ), .c(new_n340), .out0(new_n341));
  oaib12aa1n02x5               g246(.a(new_n341), .b(new_n339), .c(\a[29] ), .out0(new_n342));
  aoai13aa1n03x5               g247(.a(new_n342), .b(new_n338), .c(new_n308), .d(new_n311), .o1(new_n343));
  xorc02aa1n02x5               g248(.a(\a[30] ), .b(\b[29] ), .out0(new_n344));
  oaoi13aa1n02x5               g249(.a(new_n344), .b(new_n341), .c(new_n340), .d(new_n339), .o1(new_n345));
  aoi022aa1n03x5               g250(.a(new_n343), .b(new_n344), .c(new_n337), .d(new_n345), .o1(\s[30] ));
  nano22aa1n03x7               g251(.a(new_n329), .b(new_n332), .c(new_n344), .out0(new_n347));
  aoai13aa1n02x5               g252(.a(new_n347), .b(new_n319), .c(new_n230), .d(new_n307), .o1(new_n348));
  inv000aa1d42x5               g253(.a(new_n347), .o1(new_n349));
  norp02aa1n02x5               g254(.a(\b[29] ), .b(\a[30] ), .o1(new_n350));
  aoi022aa1n02x5               g255(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n351));
  aoi012aa1n02x5               g256(.a(new_n350), .b(new_n341), .c(new_n351), .o1(new_n352));
  aoai13aa1n03x5               g257(.a(new_n352), .b(new_n349), .c(new_n308), .d(new_n311), .o1(new_n353));
  nanb02aa1n02x5               g258(.a(\b[30] ), .b(\a[31] ), .out0(new_n354));
  nanb02aa1n02x5               g259(.a(\a[31] ), .b(\b[30] ), .out0(new_n355));
  nanp02aa1n02x5               g260(.a(new_n355), .b(new_n354), .o1(new_n356));
  oai112aa1n02x5               g261(.a(new_n354), .b(new_n355), .c(\b[29] ), .d(\a[30] ), .o1(new_n357));
  aoi012aa1n02x5               g262(.a(new_n357), .b(new_n341), .c(new_n351), .o1(new_n358));
  aoi022aa1n03x5               g263(.a(new_n353), .b(new_n356), .c(new_n348), .d(new_n358), .o1(\s[31] ));
  norb02aa1n02x5               g264(.a(new_n104), .b(new_n105), .out0(new_n360));
  xobna2aa1n03x5               g265(.a(new_n360), .b(new_n131), .c(new_n100), .out0(\s[3] ));
  aoai13aa1n02x5               g266(.a(new_n360), .b(new_n102), .c(\a[2] ), .d(\b[1] ), .o1(new_n362));
  xnbna2aa1n03x5               g267(.a(new_n103), .b(new_n362), .c(new_n104), .out0(\s[4] ));
  nano23aa1n02x4               g268(.a(new_n107), .b(new_n111), .c(new_n108), .d(new_n112), .out0(new_n364));
  oai013aa1n03x5               g269(.a(new_n364), .b(new_n103), .c(new_n102), .d(new_n106), .o1(new_n365));
  aoai13aa1n02x5               g270(.a(new_n365), .b(new_n133), .c(new_n132), .d(new_n109), .o1(\s[5] ));
  xnbna2aa1n03x5               g271(.a(new_n119), .b(new_n365), .c(new_n112), .out0(\s[6] ));
  tech160nm_fiao0012aa1n03p5x5 g272(.a(new_n119), .b(new_n365), .c(new_n112), .o(new_n368));
  xobna2aa1n03x5               g273(.a(new_n116), .b(new_n368), .c(new_n118), .out0(\s[7] ));
  aob012aa1n03x5               g274(.a(new_n116), .b(new_n368), .c(new_n118), .out0(new_n370));
  nanp02aa1n02x5               g275(.a(new_n370), .b(new_n121), .o1(new_n371));
  nano22aa1n02x4               g276(.a(new_n114), .b(new_n113), .c(new_n121), .out0(new_n372));
  aoi022aa1n02x5               g277(.a(new_n371), .b(new_n134), .c(new_n370), .d(new_n372), .o1(\s[8] ));
  aoi112aa1n02x5               g278(.a(new_n125), .b(new_n124), .c(new_n110), .d(new_n120), .o1(new_n374));
  aoi012aa1n02x5               g279(.a(new_n374), .b(new_n137), .c(new_n125), .o1(\s[9] ));
endmodule


