// Benchmark "adder" written by ABC on Thu Jul 18 08:49:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n304, new_n305, new_n306, new_n309, new_n311, new_n313;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nanp02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n09x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nor002aa1d24x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1d06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  aoi012aa1d18x5               g012(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n108));
  oaih12aa1n12x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  tech160nm_fixnrc02aa1n02p5x5 g014(.a(\b[5] ), .b(\a[6] ), .out0(new_n110));
  norp02aa1n09x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand22aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  xnrc02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  nor043aa1n06x5               g021(.a(new_n115), .b(new_n116), .c(new_n110), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\a[5] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[4] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n119), .b(new_n118), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[6] ), .b(\b[5] ), .c(new_n120), .o1(new_n121));
  aoi012aa1n02x5               g026(.a(new_n111), .b(new_n113), .c(new_n112), .o1(new_n122));
  oaib12aa1n06x5               g027(.a(new_n122), .b(new_n115), .c(new_n121), .out0(new_n123));
  xorc02aa1n12x5               g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n97), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  nor002aa1d32x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  inv040aa1n04x5               g032(.a(new_n127), .o1(new_n128));
  nand42aa1d28x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  tech160nm_fiao0012aa1n03p5x5 g034(.a(new_n123), .b(new_n109), .c(new_n117), .o(new_n130));
  oai022aa1d24x5               g035(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  aob012aa1d18x5               g036(.a(new_n131), .b(\b[9] ), .c(\a[10] ), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  aoi013aa1n06x4               g038(.a(new_n133), .b(new_n130), .c(new_n124), .d(new_n97), .o1(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n128), .c(new_n129), .out0(\s[11] ));
  nanb02aa1n02x5               g040(.a(new_n127), .b(new_n129), .out0(new_n136));
  nor042aa1d18x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand42aa1n16x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(new_n139));
  oaoi13aa1n02x7               g044(.a(new_n139), .b(new_n128), .c(new_n134), .d(new_n136), .o1(new_n140));
  oai112aa1n02x5               g045(.a(new_n128), .b(new_n139), .c(new_n134), .d(new_n136), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(\s[12] ));
  nano23aa1d15x5               g047(.a(new_n127), .b(new_n137), .c(new_n138), .d(new_n129), .out0(new_n143));
  nand23aa1d12x5               g048(.a(new_n143), .b(new_n97), .c(new_n124), .o1(new_n144));
  inv000aa1d42x5               g049(.a(new_n144), .o1(new_n145));
  aoai13aa1n06x5               g050(.a(new_n145), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n146));
  nona23aa1n09x5               g051(.a(new_n138), .b(new_n129), .c(new_n127), .d(new_n137), .out0(new_n147));
  oaoi03aa1n09x5               g052(.a(\a[12] ), .b(\b[11] ), .c(new_n128), .o1(new_n148));
  oabi12aa1n18x5               g053(.a(new_n148), .b(new_n147), .c(new_n132), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nor002aa1n20x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nand42aa1n04x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n146), .c(new_n150), .out0(\s[13] ));
  inv000aa1d42x5               g059(.a(new_n151), .o1(new_n155));
  aob012aa1n02x5               g060(.a(new_n153), .b(new_n146), .c(new_n150), .out0(new_n156));
  nor022aa1n08x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand42aa1n04x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  norb02aa1n02x5               g063(.a(new_n158), .b(new_n157), .out0(new_n159));
  xnbna2aa1n03x5               g064(.a(new_n159), .b(new_n156), .c(new_n155), .out0(\s[14] ));
  nona23aa1n02x5               g065(.a(new_n158), .b(new_n152), .c(new_n151), .d(new_n157), .out0(new_n161));
  oaih12aa1n02x5               g066(.a(new_n158), .b(new_n157), .c(new_n151), .o1(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n161), .c(new_n146), .d(new_n150), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  tech160nm_fixorc02aa1n03p5x5 g070(.a(\a[15] ), .b(\b[14] ), .out0(new_n166));
  xnrc02aa1n12x5               g071(.a(\b[15] ), .b(\a[16] ), .out0(new_n167));
  inv040aa1d30x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n165), .b(new_n168), .c(new_n163), .d(new_n166), .o1(new_n170));
  norb02aa1n03x4               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nano23aa1n06x5               g076(.a(new_n151), .b(new_n157), .c(new_n158), .d(new_n152), .out0(new_n172));
  nano32aa1d12x5               g077(.a(new_n144), .b(new_n168), .c(new_n172), .d(new_n166), .out0(new_n173));
  aoai13aa1n12x5               g078(.a(new_n173), .b(new_n123), .c(new_n109), .d(new_n117), .o1(new_n174));
  xnrc02aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .out0(new_n175));
  nor003aa1n03x5               g080(.a(new_n161), .b(new_n175), .c(new_n167), .o1(new_n176));
  nor043aa1n02x5               g081(.a(new_n167), .b(new_n175), .c(new_n162), .o1(new_n177));
  aob012aa1n02x5               g082(.a(new_n165), .b(\b[15] ), .c(\a[16] ), .out0(new_n178));
  oai012aa1n02x5               g083(.a(new_n178), .b(\b[15] ), .c(\a[16] ), .o1(new_n179));
  aoi112aa1n09x5               g084(.a(new_n179), .b(new_n177), .c(new_n149), .d(new_n176), .o1(new_n180));
  nand02aa1d08x5               g085(.a(new_n174), .b(new_n180), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g087(.a(\a[18] ), .o1(new_n183));
  inv040aa1d32x5               g088(.a(\a[17] ), .o1(new_n184));
  inv000aa1d42x5               g089(.a(\b[16] ), .o1(new_n185));
  oaoi03aa1n02x5               g090(.a(new_n184), .b(new_n185), .c(new_n181), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[17] ), .c(new_n183), .out0(\s[18] ));
  xroi22aa1d04x5               g092(.a(new_n184), .b(\b[16] ), .c(new_n183), .d(\b[17] ), .out0(new_n188));
  nanp02aa1n02x5               g093(.a(new_n185), .b(new_n184), .o1(new_n189));
  oaoi03aa1n12x5               g094(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n190));
  aoi012aa1n12x5               g095(.a(new_n190), .b(new_n181), .c(new_n188), .o1(new_n191));
  nor042aa1n09x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  nand42aa1n04x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n191), .b(new_n194), .c(new_n193), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g101(.a(new_n192), .b(new_n194), .out0(new_n197));
  nor002aa1n04x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nand42aa1n06x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  oaoi13aa1n02x7               g105(.a(new_n200), .b(new_n193), .c(new_n191), .d(new_n197), .o1(new_n201));
  nor042aa1n03x5               g106(.a(new_n191), .b(new_n197), .o1(new_n202));
  nano22aa1n03x5               g107(.a(new_n202), .b(new_n193), .c(new_n200), .out0(new_n203));
  norp02aa1n03x5               g108(.a(new_n201), .b(new_n203), .o1(\s[20] ));
  nano23aa1n03x7               g109(.a(new_n192), .b(new_n198), .c(new_n199), .d(new_n194), .out0(new_n205));
  nanp02aa1n02x5               g110(.a(new_n188), .b(new_n205), .o1(new_n206));
  oai022aa1n02x5               g111(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n207));
  oaib12aa1n09x5               g112(.a(new_n207), .b(new_n183), .c(\b[17] ), .out0(new_n208));
  nona23aa1n09x5               g113(.a(new_n199), .b(new_n194), .c(new_n192), .d(new_n198), .out0(new_n209));
  aoi012aa1n09x5               g114(.a(new_n198), .b(new_n192), .c(new_n199), .o1(new_n210));
  oai012aa1n18x5               g115(.a(new_n210), .b(new_n209), .c(new_n208), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n206), .c(new_n174), .d(new_n180), .o1(new_n213));
  xorb03aa1n02x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  xorc02aa1n02x5               g121(.a(\a[22] ), .b(\b[21] ), .out0(new_n217));
  aoai13aa1n03x5               g122(.a(new_n217), .b(new_n215), .c(new_n213), .d(new_n216), .o1(new_n218));
  aoi112aa1n02x5               g123(.a(new_n215), .b(new_n217), .c(new_n213), .d(new_n216), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n218), .b(new_n219), .out0(\s[22] ));
  inv000aa1d42x5               g125(.a(\a[21] ), .o1(new_n221));
  inv040aa1d32x5               g126(.a(\a[22] ), .o1(new_n222));
  xroi22aa1d06x4               g127(.a(new_n221), .b(\b[20] ), .c(new_n222), .d(\b[21] ), .out0(new_n223));
  nanp03aa1n02x5               g128(.a(new_n223), .b(new_n188), .c(new_n205), .o1(new_n224));
  inv000aa1d42x5               g129(.a(\b[21] ), .o1(new_n225));
  oao003aa1n02x5               g130(.a(new_n222), .b(new_n225), .c(new_n215), .carry(new_n226));
  aoi012aa1n02x5               g131(.a(new_n226), .b(new_n211), .c(new_n223), .o1(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n174), .d(new_n180), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g134(.a(\b[22] ), .b(\a[23] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[23] ), .b(\b[22] ), .out0(new_n231));
  xorc02aa1n02x5               g136(.a(\a[24] ), .b(\b[23] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n230), .c(new_n228), .d(new_n231), .o1(new_n233));
  aoi112aa1n02x5               g138(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n233), .b(new_n234), .out0(\s[24] ));
  inv000aa1d42x5               g140(.a(\a[23] ), .o1(new_n236));
  inv040aa1d32x5               g141(.a(\a[24] ), .o1(new_n237));
  xroi22aa1d06x4               g142(.a(new_n236), .b(\b[22] ), .c(new_n237), .d(\b[23] ), .out0(new_n238));
  nano22aa1n02x4               g143(.a(new_n206), .b(new_n223), .c(new_n238), .out0(new_n239));
  inv000aa1n03x5               g144(.a(new_n210), .o1(new_n240));
  aoai13aa1n06x5               g145(.a(new_n223), .b(new_n240), .c(new_n205), .d(new_n190), .o1(new_n241));
  inv000aa1n02x5               g146(.a(new_n226), .o1(new_n242));
  inv000aa1n02x5               g147(.a(new_n238), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n244));
  aoib12aa1n02x5               g149(.a(new_n244), .b(new_n237), .c(\b[23] ), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n242), .o1(new_n246));
  xorc02aa1n02x5               g151(.a(\a[25] ), .b(\b[24] ), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n246), .c(new_n181), .d(new_n239), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n247), .b(new_n246), .c(new_n181), .d(new_n239), .o1(new_n249));
  norb02aa1n03x4               g154(.a(new_n248), .b(new_n249), .out0(\s[25] ));
  nor042aa1n03x5               g155(.a(\b[24] ), .b(\a[25] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[26] ), .b(\b[25] ), .out0(new_n253));
  aobi12aa1n06x5               g158(.a(new_n253), .b(new_n248), .c(new_n252), .out0(new_n254));
  nona22aa1n02x5               g159(.a(new_n248), .b(new_n253), .c(new_n251), .out0(new_n255));
  norb02aa1n03x4               g160(.a(new_n255), .b(new_n254), .out0(\s[26] ));
  inv000aa1d42x5               g161(.a(\a[25] ), .o1(new_n257));
  inv020aa1n04x5               g162(.a(\a[26] ), .o1(new_n258));
  xroi22aa1d06x4               g163(.a(new_n257), .b(\b[24] ), .c(new_n258), .d(\b[25] ), .out0(new_n259));
  nano32aa1n03x7               g164(.a(new_n206), .b(new_n259), .c(new_n223), .d(new_n238), .out0(new_n260));
  nand02aa1d06x5               g165(.a(new_n181), .b(new_n260), .o1(new_n261));
  oao003aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .c(new_n252), .carry(new_n262));
  aobi12aa1n06x5               g167(.a(new_n262), .b(new_n246), .c(new_n259), .out0(new_n263));
  xorc02aa1n02x5               g168(.a(\a[27] ), .b(\b[26] ), .out0(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n263), .c(new_n261), .out0(\s[27] ));
  norp02aa1n02x5               g170(.a(\b[26] ), .b(\a[27] ), .o1(new_n266));
  inv040aa1n03x5               g171(.a(new_n266), .o1(new_n267));
  aobi12aa1n06x5               g172(.a(new_n260), .b(new_n174), .c(new_n180), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n238), .b(new_n226), .c(new_n211), .d(new_n223), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n259), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n262), .b(new_n270), .c(new_n269), .d(new_n245), .o1(new_n271));
  oaih12aa1n02x5               g176(.a(new_n264), .b(new_n271), .c(new_n268), .o1(new_n272));
  xnrc02aa1n02x5               g177(.a(\b[27] ), .b(\a[28] ), .out0(new_n273));
  tech160nm_fiaoi012aa1n02p5x5 g178(.a(new_n273), .b(new_n272), .c(new_n267), .o1(new_n274));
  aobi12aa1n06x5               g179(.a(new_n264), .b(new_n263), .c(new_n261), .out0(new_n275));
  nano22aa1n03x7               g180(.a(new_n275), .b(new_n267), .c(new_n273), .out0(new_n276));
  norp02aa1n03x5               g181(.a(new_n274), .b(new_n276), .o1(\s[28] ));
  norb02aa1n02x5               g182(.a(new_n264), .b(new_n273), .out0(new_n278));
  oaih12aa1n02x5               g183(.a(new_n278), .b(new_n271), .c(new_n268), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[28] ), .b(\b[27] ), .c(new_n267), .carry(new_n280));
  xnrc02aa1n02x5               g185(.a(\b[28] ), .b(\a[29] ), .out0(new_n281));
  tech160nm_fiaoi012aa1n02p5x5 g186(.a(new_n281), .b(new_n279), .c(new_n280), .o1(new_n282));
  aobi12aa1n06x5               g187(.a(new_n278), .b(new_n263), .c(new_n261), .out0(new_n283));
  nano22aa1n03x7               g188(.a(new_n283), .b(new_n280), .c(new_n281), .out0(new_n284));
  norp02aa1n03x5               g189(.a(new_n282), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g190(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g191(.a(new_n264), .b(new_n281), .c(new_n273), .out0(new_n287));
  oaih12aa1n02x5               g192(.a(new_n287), .b(new_n271), .c(new_n268), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n280), .carry(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  tech160nm_fiaoi012aa1n02p5x5 g195(.a(new_n290), .b(new_n288), .c(new_n289), .o1(new_n291));
  aobi12aa1n06x5               g196(.a(new_n287), .b(new_n263), .c(new_n261), .out0(new_n292));
  nano22aa1n03x7               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  norp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[30] ));
  norb02aa1n02x5               g199(.a(new_n287), .b(new_n290), .out0(new_n295));
  aobi12aa1n06x5               g200(.a(new_n295), .b(new_n263), .c(new_n261), .out0(new_n296));
  oao003aa1n02x5               g201(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[30] ), .b(\a[31] ), .out0(new_n298));
  nano22aa1n03x7               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  oaih12aa1n02x5               g204(.a(new_n295), .b(new_n271), .c(new_n268), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  norp02aa1n03x5               g206(.a(new_n301), .b(new_n299), .o1(\s[31] ));
  xnrb03aa1n02x5               g207(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g208(.a(new_n103), .o1(new_n304));
  nona22aa1n02x4               g209(.a(new_n106), .b(new_n102), .c(new_n105), .out0(new_n305));
  aoi012aa1n02x5               g210(.a(new_n105), .b(new_n304), .c(new_n104), .o1(new_n306));
  aoi022aa1n02x5               g211(.a(new_n109), .b(new_n304), .c(new_n305), .d(new_n306), .o1(\s[4] ));
  xorb03aa1n02x5               g212(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g213(.a(new_n118), .b(new_n119), .c(new_n109), .o1(new_n309));
  xnrb03aa1n02x5               g214(.a(new_n309), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n02x5               g215(.a(\a[6] ), .b(\b[5] ), .c(new_n309), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g217(.a(new_n113), .b(new_n311), .c(new_n114), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g219(.a(new_n130), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


