// Benchmark "adder" written by ABC on Thu Jul 18 09:18:28 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n305, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n323,
    new_n325, new_n328, new_n329, new_n331, new_n332, new_n333, new_n335,
    new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d32x5               g001(.a(\a[10] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[9] ), .o1(new_n98));
  nand02aa1n06x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand02aa1d08x5               g004(.a(\b[9] ), .b(\a[10] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(new_n99), .b(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(new_n101), .o1(new_n102));
  orn002aa1n24x5               g007(.a(\a[9] ), .b(\b[8] ), .o(new_n103));
  nand42aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n08x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor002aa1n12x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  oai012aa1n02x7               g011(.a(new_n104), .b(new_n106), .c(new_n105), .o1(new_n107));
  norb02aa1n06x5               g012(.a(new_n104), .b(new_n105), .out0(new_n108));
  nand42aa1n08x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  norb02aa1n03x5               g014(.a(new_n109), .b(new_n106), .out0(new_n110));
  nor042aa1n02x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  aoi022aa1d24x5               g016(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n112));
  oai112aa1n06x5               g017(.a(new_n108), .b(new_n110), .c(new_n111), .d(new_n112), .o1(new_n113));
  nanp02aa1n06x5               g018(.a(new_n113), .b(new_n107), .o1(new_n114));
  nand42aa1d28x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor002aa1d24x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  tech160nm_fixnrc02aa1n04x5   g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  nor022aa1n04x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nanp02aa1n04x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  nor022aa1n16x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nand42aa1n03x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  nona23aa1n09x5               g027(.a(new_n122), .b(new_n120), .c(new_n119), .d(new_n121), .out0(new_n123));
  nor043aa1n04x5               g028(.a(new_n123), .b(new_n118), .c(new_n117), .o1(new_n124));
  inv040aa1d32x5               g029(.a(\a[5] ), .o1(new_n125));
  inv040aa1d28x5               g030(.a(\b[4] ), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n115), .b(new_n116), .c(new_n126), .d(new_n125), .o1(new_n127));
  oai012aa1n02x5               g032(.a(new_n120), .b(new_n121), .c(new_n119), .o1(new_n128));
  oai012aa1n12x5               g033(.a(new_n128), .b(new_n123), .c(new_n127), .o1(new_n129));
  nand02aa1d24x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nand42aa1d28x5               g035(.a(new_n103), .b(new_n130), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  aoai13aa1n06x5               g037(.a(new_n132), .b(new_n129), .c(new_n114), .d(new_n124), .o1(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n102), .b(new_n133), .c(new_n103), .out0(\s[10] ));
  nanp03aa1n02x5               g039(.a(new_n133), .b(new_n102), .c(new_n103), .o1(new_n135));
  nor002aa1n16x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand42aa1d28x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanb02aa1n03x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n135), .c(new_n100), .out0(\s[11] ));
  aoi013aa1n02x4               g044(.a(new_n136), .b(new_n135), .c(new_n100), .d(new_n137), .o1(new_n140));
  xnrb03aa1n02x5               g045(.a(new_n140), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n06x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand42aa1n10x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nano23aa1d15x5               g048(.a(new_n136), .b(new_n142), .c(new_n143), .d(new_n137), .out0(new_n144));
  nona22aa1d36x5               g049(.a(new_n144), .b(new_n131), .c(new_n101), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  aoai13aa1n02x5               g051(.a(new_n146), .b(new_n129), .c(new_n114), .d(new_n124), .o1(new_n147));
  nanb02aa1n02x5               g052(.a(new_n142), .b(new_n143), .out0(new_n148));
  oai022aa1n02x5               g053(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n149));
  nano23aa1n06x5               g054(.a(new_n148), .b(new_n138), .c(new_n149), .d(new_n100), .out0(new_n150));
  oa0012aa1n02x5               g055(.a(new_n143), .b(new_n142), .c(new_n136), .o(new_n151));
  norp02aa1n02x5               g056(.a(new_n150), .b(new_n151), .o1(new_n152));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n03x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  xnbna2aa1n03x5               g060(.a(new_n155), .b(new_n147), .c(new_n152), .out0(\s[13] ));
  inv000aa1d42x5               g061(.a(new_n153), .o1(new_n157));
  nanb02aa1n02x5               g062(.a(new_n153), .b(new_n154), .out0(new_n158));
  aoai13aa1n02x5               g063(.a(new_n157), .b(new_n158), .c(new_n147), .d(new_n152), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nanp02aa1n03x5               g065(.a(new_n147), .b(new_n152), .o1(new_n161));
  inv040aa1d32x5               g066(.a(\a[14] ), .o1(new_n162));
  inv040aa1d28x5               g067(.a(\b[13] ), .o1(new_n163));
  nand02aa1d12x5               g068(.a(new_n163), .b(new_n162), .o1(new_n164));
  nanp02aa1n12x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand02aa1d06x5               g070(.a(new_n164), .b(new_n165), .o1(new_n166));
  nona22aa1n02x4               g071(.a(new_n161), .b(new_n158), .c(new_n166), .out0(new_n167));
  oaoi03aa1n12x5               g072(.a(new_n162), .b(new_n163), .c(new_n153), .o1(new_n168));
  nor002aa1d32x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand42aa1n04x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n167), .c(new_n168), .out0(\s[15] ));
  inv000aa1d42x5               g077(.a(new_n166), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n168), .o1(new_n174));
  aoi013aa1n02x4               g079(.a(new_n174), .b(new_n161), .c(new_n155), .d(new_n173), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n169), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n171), .o1(new_n177));
  nor022aa1n06x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand42aa1n03x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  oaoi13aa1n02x7               g086(.a(new_n181), .b(new_n176), .c(new_n175), .d(new_n177), .o1(new_n182));
  aoi012aa1n02x5               g087(.a(new_n177), .b(new_n167), .c(new_n168), .o1(new_n183));
  nano22aa1n02x4               g088(.a(new_n183), .b(new_n176), .c(new_n181), .out0(new_n184));
  norp02aa1n02x5               g089(.a(new_n182), .b(new_n184), .o1(\s[16] ));
  nano23aa1n02x4               g090(.a(new_n169), .b(new_n178), .c(new_n179), .d(new_n170), .out0(new_n186));
  nona22aa1n03x5               g091(.a(new_n186), .b(new_n158), .c(new_n166), .out0(new_n187));
  nor042aa1n06x5               g092(.a(new_n187), .b(new_n145), .o1(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n129), .c(new_n114), .d(new_n124), .o1(new_n189));
  nona23aa1n02x5               g094(.a(new_n179), .b(new_n170), .c(new_n169), .d(new_n178), .out0(new_n190));
  nano32aa1n02x5               g095(.a(new_n190), .b(new_n155), .c(new_n164), .d(new_n165), .out0(new_n191));
  oaoi03aa1n02x5               g096(.a(\a[16] ), .b(\b[15] ), .c(new_n176), .o1(new_n192));
  oabi12aa1n03x5               g097(.a(new_n192), .b(new_n190), .c(new_n168), .out0(new_n193));
  oaoi13aa1n09x5               g098(.a(new_n193), .b(new_n191), .c(new_n150), .d(new_n151), .o1(new_n194));
  xorc02aa1n06x5               g099(.a(\a[17] ), .b(\b[16] ), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n189), .c(new_n194), .out0(\s[17] ));
  inv000aa1d42x5               g101(.a(\a[17] ), .o1(new_n197));
  inv000aa1d48x5               g102(.a(\b[16] ), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(new_n198), .b(new_n197), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n195), .o1(new_n200));
  aoai13aa1n02x5               g105(.a(new_n199), .b(new_n200), .c(new_n189), .d(new_n194), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n06x5               g107(.a(new_n189), .b(new_n194), .o1(new_n203));
  nor042aa1d18x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nand42aa1n06x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nanb02aa1n03x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  nona22aa1n03x5               g111(.a(new_n203), .b(new_n200), .c(new_n206), .out0(new_n207));
  aoai13aa1n12x5               g112(.a(new_n205), .b(new_n204), .c(new_n197), .d(new_n198), .o1(new_n208));
  nor042aa1n06x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand42aa1n08x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n207), .c(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g118(.a(new_n209), .o1(new_n214));
  aoi112aa1n03x4               g119(.a(new_n206), .b(new_n200), .c(new_n189), .d(new_n194), .o1(new_n215));
  inv040aa1n03x5               g120(.a(new_n208), .o1(new_n216));
  oai012aa1n02x5               g121(.a(new_n211), .b(new_n215), .c(new_n216), .o1(new_n217));
  nor042aa1n02x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand42aa1n06x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nanb02aa1n02x5               g124(.a(new_n218), .b(new_n219), .out0(new_n220));
  tech160nm_fiaoi012aa1n02p5x5 g125(.a(new_n220), .b(new_n217), .c(new_n214), .o1(new_n221));
  aobi12aa1n06x5               g126(.a(new_n211), .b(new_n207), .c(new_n208), .out0(new_n222));
  nano22aa1n03x7               g127(.a(new_n222), .b(new_n214), .c(new_n220), .out0(new_n223));
  norp02aa1n02x5               g128(.a(new_n221), .b(new_n223), .o1(\s[20] ));
  inv000aa1d42x5               g129(.a(new_n206), .o1(new_n225));
  nano23aa1n09x5               g130(.a(new_n209), .b(new_n218), .c(new_n219), .d(new_n210), .out0(new_n226));
  nand03aa1n06x5               g131(.a(new_n226), .b(new_n225), .c(new_n195), .o1(new_n227));
  aoi012aa1n06x5               g132(.a(new_n227), .b(new_n189), .c(new_n194), .o1(new_n228));
  nona23aa1n09x5               g133(.a(new_n219), .b(new_n210), .c(new_n209), .d(new_n218), .out0(new_n229));
  oaoi03aa1n09x5               g134(.a(\a[20] ), .b(\b[19] ), .c(new_n214), .o1(new_n230));
  inv040aa1n03x5               g135(.a(new_n230), .o1(new_n231));
  oai012aa1n12x5               g136(.a(new_n231), .b(new_n229), .c(new_n208), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[20] ), .b(\a[21] ), .out0(new_n233));
  oabi12aa1n06x5               g138(.a(new_n233), .b(new_n228), .c(new_n232), .out0(new_n234));
  norb03aa1n02x5               g139(.a(new_n233), .b(new_n228), .c(new_n232), .out0(new_n235));
  norb02aa1n02x5               g140(.a(new_n234), .b(new_n235), .out0(\s[21] ));
  orn002aa1n24x5               g141(.a(\a[21] ), .b(\b[20] ), .o(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[21] ), .b(\a[22] ), .out0(new_n238));
  tech160nm_fiaoi012aa1n02p5x5 g143(.a(new_n238), .b(new_n234), .c(new_n237), .o1(new_n239));
  nanp03aa1n03x5               g144(.a(new_n234), .b(new_n237), .c(new_n238), .o1(new_n240));
  norb02aa1n03x4               g145(.a(new_n240), .b(new_n239), .out0(\s[22] ));
  nor042aa1n04x5               g146(.a(new_n238), .b(new_n233), .o1(new_n242));
  oaoi03aa1n09x5               g147(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .o1(new_n243));
  aoi012aa1d18x5               g148(.a(new_n243), .b(new_n232), .c(new_n242), .o1(new_n244));
  nona32aa1n03x5               g149(.a(new_n203), .b(new_n238), .c(new_n233), .d(new_n227), .out0(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[22] ), .b(\a[23] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xnbna2aa1n03x5               g152(.a(new_n247), .b(new_n245), .c(new_n244), .out0(\s[23] ));
  orn002aa1n24x5               g153(.a(\a[23] ), .b(\b[22] ), .o(new_n249));
  inv000aa1d42x5               g154(.a(new_n244), .o1(new_n250));
  aoai13aa1n03x5               g155(.a(new_n247), .b(new_n250), .c(new_n228), .d(new_n242), .o1(new_n251));
  xnrc02aa1n12x5               g156(.a(\b[23] ), .b(\a[24] ), .out0(new_n252));
  aoi012aa1n03x5               g157(.a(new_n252), .b(new_n251), .c(new_n249), .o1(new_n253));
  tech160nm_fiaoi012aa1n04x5   g158(.a(new_n246), .b(new_n245), .c(new_n244), .o1(new_n254));
  nano22aa1n03x7               g159(.a(new_n254), .b(new_n249), .c(new_n252), .out0(new_n255));
  nor002aa1n02x5               g160(.a(new_n253), .b(new_n255), .o1(\s[24] ));
  aoai13aa1n06x5               g161(.a(new_n242), .b(new_n230), .c(new_n226), .d(new_n216), .o1(new_n257));
  inv000aa1n04x5               g162(.a(new_n243), .o1(new_n258));
  nor042aa1n02x5               g163(.a(new_n252), .b(new_n246), .o1(new_n259));
  inv000aa1n03x5               g164(.a(new_n259), .o1(new_n260));
  tech160nm_fioaoi03aa1n02p5x5 g165(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .o1(new_n261));
  inv000aa1n03x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n12x5               g167(.a(new_n262), .b(new_n260), .c(new_n257), .d(new_n258), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  nanp02aa1n02x5               g169(.a(new_n259), .b(new_n242), .o1(new_n265));
  nona22aa1n03x5               g170(.a(new_n203), .b(new_n227), .c(new_n265), .out0(new_n266));
  xnrc02aa1n12x5               g171(.a(\b[24] ), .b(\a[25] ), .out0(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  xnbna2aa1n03x5               g173(.a(new_n268), .b(new_n266), .c(new_n264), .out0(\s[25] ));
  nor042aa1n03x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoi112aa1n03x4               g176(.a(new_n265), .b(new_n227), .c(new_n189), .d(new_n194), .o1(new_n272));
  oai012aa1n02x7               g177(.a(new_n268), .b(new_n272), .c(new_n263), .o1(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[25] ), .b(\a[26] ), .out0(new_n274));
  tech160nm_fiaoi012aa1n02p5x5 g179(.a(new_n274), .b(new_n273), .c(new_n271), .o1(new_n275));
  tech160nm_fiaoi012aa1n05x5   g180(.a(new_n267), .b(new_n266), .c(new_n264), .o1(new_n276));
  nano22aa1n03x7               g181(.a(new_n276), .b(new_n271), .c(new_n274), .out0(new_n277));
  nor002aa1n02x5               g182(.a(new_n275), .b(new_n277), .o1(\s[26] ));
  xorc02aa1n02x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  nor042aa1n04x5               g184(.a(new_n274), .b(new_n267), .o1(new_n280));
  oao003aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n281));
  aobi12aa1n12x5               g186(.a(new_n281), .b(new_n263), .c(new_n280), .out0(new_n282));
  inv000aa1d42x5               g187(.a(new_n280), .o1(new_n283));
  nona32aa1n09x5               g188(.a(new_n203), .b(new_n283), .c(new_n265), .d(new_n227), .out0(new_n284));
  xnbna2aa1n03x5               g189(.a(new_n279), .b(new_n282), .c(new_n284), .out0(\s[27] ));
  norp02aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  inv040aa1n03x5               g191(.a(new_n286), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n259), .b(new_n243), .c(new_n232), .d(new_n242), .o1(new_n288));
  aoai13aa1n04x5               g193(.a(new_n281), .b(new_n283), .c(new_n288), .d(new_n262), .o1(new_n289));
  nano22aa1n02x4               g194(.a(new_n283), .b(new_n242), .c(new_n259), .out0(new_n290));
  aoai13aa1n03x5               g195(.a(new_n279), .b(new_n289), .c(new_n228), .d(new_n290), .o1(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .out0(new_n292));
  aoi012aa1n02x7               g197(.a(new_n292), .b(new_n291), .c(new_n287), .o1(new_n293));
  aobi12aa1n02x7               g198(.a(new_n279), .b(new_n282), .c(new_n284), .out0(new_n294));
  nano22aa1n03x5               g199(.a(new_n294), .b(new_n287), .c(new_n292), .out0(new_n295));
  nor002aa1n02x5               g200(.a(new_n293), .b(new_n295), .o1(\s[28] ));
  xnrc02aa1n02x5               g201(.a(\b[28] ), .b(\a[29] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n279), .b(new_n292), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n289), .c(new_n228), .d(new_n290), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n300));
  aoi012aa1n03x5               g205(.a(new_n297), .b(new_n299), .c(new_n300), .o1(new_n301));
  aobi12aa1n03x5               g206(.a(new_n298), .b(new_n282), .c(new_n284), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n297), .c(new_n300), .out0(new_n303));
  nor002aa1n02x5               g208(.a(new_n301), .b(new_n303), .o1(\s[29] ));
  nanp02aa1n02x5               g209(.a(\b[0] ), .b(\a[1] ), .o1(new_n305));
  xorb03aa1n02x5               g210(.a(new_n305), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g211(.a(\b[29] ), .b(\a[30] ), .out0(new_n307));
  norb03aa1n02x5               g212(.a(new_n279), .b(new_n297), .c(new_n292), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n289), .c(new_n228), .d(new_n290), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n310));
  aoi012aa1n03x5               g215(.a(new_n307), .b(new_n309), .c(new_n310), .o1(new_n311));
  aobi12aa1n03x5               g216(.a(new_n308), .b(new_n282), .c(new_n284), .out0(new_n312));
  nano22aa1n03x5               g217(.a(new_n312), .b(new_n307), .c(new_n310), .out0(new_n313));
  nor002aa1n02x5               g218(.a(new_n311), .b(new_n313), .o1(\s[30] ));
  norb02aa1n02x5               g219(.a(new_n308), .b(new_n307), .out0(new_n315));
  aobi12aa1n06x5               g220(.a(new_n315), .b(new_n282), .c(new_n284), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n310), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  nano22aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n318), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n315), .b(new_n289), .c(new_n228), .d(new_n290), .o1(new_n320));
  aoi012aa1n03x5               g225(.a(new_n318), .b(new_n320), .c(new_n317), .o1(new_n321));
  norp02aa1n03x5               g226(.a(new_n321), .b(new_n319), .o1(\s[31] ));
  norp02aa1n02x5               g227(.a(new_n112), .b(new_n111), .o1(new_n323));
  xnrb03aa1n02x5               g228(.a(new_n323), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi13aa1n02x5               g229(.a(new_n106), .b(new_n109), .c(new_n112), .d(new_n111), .o1(new_n325));
  xnrc02aa1n02x5               g230(.a(new_n325), .b(new_n108), .out0(\s[4] ));
  xobna2aa1n03x5               g231(.a(new_n118), .b(new_n113), .c(new_n107), .out0(\s[5] ));
  nanp02aa1n02x5               g232(.a(new_n126), .b(new_n125), .o1(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n118), .c(new_n113), .d(new_n107), .o1(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g235(.a(new_n127), .o1(new_n331));
  aoi112aa1n02x5               g236(.a(new_n117), .b(new_n118), .c(new_n113), .d(new_n107), .o1(new_n332));
  norp02aa1n02x5               g237(.a(new_n332), .b(new_n331), .o1(new_n333));
  xnrb03aa1n02x5               g238(.a(new_n333), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi13aa1n02x5               g239(.a(new_n121), .b(new_n122), .c(new_n332), .d(new_n331), .o1(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  aoi112aa1n02x5               g241(.a(new_n132), .b(new_n129), .c(new_n114), .d(new_n124), .o1(new_n337));
  norb02aa1n02x5               g242(.a(new_n133), .b(new_n337), .out0(\s[9] ));
endmodule


