// Benchmark "adder" written by ABC on Wed Jul 17 17:25:13 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n325, new_n328, new_n330, new_n331, new_n333, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n06x5               g001(.a(\b[3] ), .b(\a[4] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  tech160nm_finor002aa1n05x5   g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  ao0012aa1n03x7               g004(.a(new_n97), .b(new_n99), .c(new_n98), .o(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[1] ), .o1(new_n102));
  nand22aa1n03x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  tech160nm_fioaoi03aa1n03p5x5 g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  nand42aa1n16x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n02x4               g010(.a(new_n105), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n106));
  oabi12aa1n06x5               g011(.a(new_n100), .b(new_n106), .c(new_n104), .out0(new_n107));
  nand02aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor002aa1n20x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand02aa1d24x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor002aa1d32x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n02x4               g016(.a(new_n110), .b(new_n108), .c(new_n111), .d(new_n109), .out0(new_n112));
  tech160nm_fixorc02aa1n02p5x5 g017(.a(\a[5] ), .b(\b[4] ), .out0(new_n113));
  tech160nm_fixorc02aa1n04x5   g018(.a(\a[6] ), .b(\b[5] ), .out0(new_n114));
  nano22aa1n03x7               g019(.a(new_n112), .b(new_n113), .c(new_n114), .out0(new_n115));
  inv000aa1d42x5               g020(.a(new_n110), .o1(new_n116));
  orn002aa1n12x5               g021(.a(\a[6] ), .b(\b[5] ), .o(new_n117));
  norp02aa1n02x5               g022(.a(new_n111), .b(new_n109), .o1(new_n118));
  nanp02aa1n03x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nona22aa1n03x5               g024(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .out0(new_n120));
  aoai13aa1n06x5               g025(.a(new_n118), .b(new_n116), .c(new_n120), .d(new_n117), .o1(new_n121));
  nand42aa1n04x5               g026(.a(new_n121), .b(new_n108), .o1(new_n122));
  inv040aa1n02x5               g027(.a(new_n122), .o1(new_n123));
  nor002aa1d32x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nanp02aa1n04x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n06x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n123), .c(new_n107), .d(new_n115), .o1(new_n127));
  nor002aa1d32x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand02aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n15x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  oaoi13aa1n04x5               g036(.a(new_n131), .b(new_n127), .c(\a[9] ), .d(\b[8] ), .o1(new_n132));
  oao003aa1n03x5               g037(.a(new_n101), .b(new_n102), .c(new_n103), .carry(new_n133));
  nano23aa1n03x5               g038(.a(new_n97), .b(new_n99), .c(new_n105), .d(new_n98), .out0(new_n134));
  tech160nm_fiaoi012aa1n05x5   g039(.a(new_n100), .b(new_n134), .c(new_n133), .o1(new_n135));
  nanb02aa1n06x5               g040(.a(new_n109), .b(new_n108), .out0(new_n136));
  nanb02aa1d24x5               g041(.a(new_n111), .b(new_n110), .out0(new_n137));
  nona23aa1n09x5               g042(.a(new_n113), .b(new_n114), .c(new_n137), .d(new_n136), .out0(new_n138));
  oai012aa1n02x5               g043(.a(new_n122), .b(new_n135), .c(new_n138), .o1(new_n139));
  aoi112aa1n02x5               g044(.a(new_n130), .b(new_n124), .c(new_n139), .d(new_n125), .o1(new_n140));
  norp02aa1n02x5               g045(.a(new_n132), .b(new_n140), .o1(\s[10] ));
  oai012aa1n12x5               g046(.a(new_n129), .b(new_n128), .c(new_n124), .o1(new_n142));
  inv020aa1n04x5               g047(.a(new_n142), .o1(new_n143));
  nand02aa1d28x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nor002aa1d32x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n144), .b(new_n145), .out0(new_n146));
  oabi12aa1n02x5               g051(.a(new_n146), .b(new_n132), .c(new_n143), .out0(new_n147));
  nano22aa1n03x5               g052(.a(new_n132), .b(new_n142), .c(new_n146), .out0(new_n148));
  nanb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(\s[11] ));
  nor002aa1d24x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand02aa1d16x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  aoai13aa1n02x7               g057(.a(new_n152), .b(new_n148), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  nona22aa1n03x5               g058(.a(new_n144), .b(new_n148), .c(new_n152), .out0(new_n154));
  nanp02aa1n03x5               g059(.a(new_n154), .b(new_n153), .o1(\s[12] ));
  nona23aa1d24x5               g060(.a(new_n144), .b(new_n151), .c(new_n150), .d(new_n145), .out0(new_n156));
  nano22aa1d15x5               g061(.a(new_n156), .b(new_n126), .c(new_n130), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n123), .c(new_n107), .d(new_n115), .o1(new_n158));
  oa0012aa1n03x5               g063(.a(new_n151), .b(new_n150), .c(new_n145), .o(new_n159));
  oabi12aa1n18x5               g064(.a(new_n159), .b(new_n142), .c(new_n156), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  nand42aa1d28x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nor002aa1n16x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanb02aa1n03x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  xobna2aa1n03x5               g069(.a(new_n164), .b(new_n158), .c(new_n161), .out0(\s[13] ));
  nanp02aa1n02x5               g070(.a(new_n158), .b(new_n161), .o1(new_n166));
  nor002aa1n12x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand42aa1n20x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nanb02aa1n03x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n163), .c(new_n166), .d(new_n162), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n169), .b(new_n163), .c(new_n166), .d(new_n162), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(\s[14] ));
  nano23aa1d15x5               g077(.a(new_n167), .b(new_n163), .c(new_n168), .d(new_n162), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  oai012aa1n12x5               g079(.a(new_n168), .b(new_n167), .c(new_n163), .o1(new_n175));
  aoai13aa1n04x5               g080(.a(new_n175), .b(new_n174), .c(new_n158), .d(new_n161), .o1(new_n176));
  xorb03aa1n02x5               g081(.a(new_n176), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nand42aa1n06x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nor002aa1d24x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nor022aa1n16x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanp02aa1n06x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  aoai13aa1n02x5               g087(.a(new_n182), .b(new_n179), .c(new_n176), .d(new_n178), .o1(new_n183));
  aoi112aa1n03x5               g088(.a(new_n182), .b(new_n179), .c(new_n176), .d(new_n178), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n184), .b(new_n183), .out0(\s[16] ));
  nano23aa1n03x7               g090(.a(new_n150), .b(new_n145), .c(new_n151), .d(new_n144), .out0(new_n186));
  nano23aa1n03x7               g091(.a(new_n180), .b(new_n179), .c(new_n181), .d(new_n178), .out0(new_n187));
  nand42aa1n02x5               g092(.a(new_n187), .b(new_n173), .o1(new_n188));
  nano32aa1n02x5               g093(.a(new_n188), .b(new_n186), .c(new_n130), .d(new_n126), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n123), .c(new_n107), .d(new_n115), .o1(new_n190));
  oai012aa1n02x5               g095(.a(new_n181), .b(new_n180), .c(new_n179), .o1(new_n191));
  inv000aa1d42x5               g096(.a(new_n175), .o1(new_n192));
  aoai13aa1n09x5               g097(.a(new_n187), .b(new_n192), .c(new_n160), .d(new_n173), .o1(new_n193));
  nand23aa1n06x5               g098(.a(new_n190), .b(new_n193), .c(new_n191), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1n09x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nona23aa1n09x5               g102(.a(new_n178), .b(new_n181), .c(new_n180), .d(new_n179), .out0(new_n198));
  nona32aa1n03x5               g103(.a(new_n157), .b(new_n198), .c(new_n169), .d(new_n164), .out0(new_n199));
  oaoi13aa1n09x5               g104(.a(new_n199), .b(new_n122), .c(new_n135), .d(new_n138), .o1(new_n200));
  aoai13aa1n04x5               g105(.a(new_n173), .b(new_n159), .c(new_n186), .d(new_n143), .o1(new_n201));
  aoai13aa1n06x5               g106(.a(new_n191), .b(new_n198), .c(new_n201), .d(new_n175), .o1(new_n202));
  oai013aa1n02x4               g107(.a(new_n197), .b(new_n202), .c(new_n200), .d(new_n196), .o1(new_n203));
  xnrb03aa1n02x5               g108(.a(new_n203), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor002aa1n04x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nand22aa1n04x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nano23aa1n06x5               g111(.a(new_n196), .b(new_n205), .c(new_n206), .d(new_n197), .out0(new_n207));
  oaih12aa1n02x5               g112(.a(new_n207), .b(new_n202), .c(new_n200), .o1(new_n208));
  tech160nm_fiaoi012aa1n04x5   g113(.a(new_n205), .b(new_n196), .c(new_n206), .o1(new_n209));
  nand02aa1n04x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nor042aa1n04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  norb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n208), .c(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g119(.a(new_n208), .b(new_n209), .o1(new_n215));
  nor042aa1n02x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nanp02aa1n06x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nanb02aa1n02x5               g122(.a(new_n216), .b(new_n217), .out0(new_n218));
  aoai13aa1n03x5               g123(.a(new_n218), .b(new_n211), .c(new_n215), .d(new_n212), .o1(new_n219));
  inv020aa1n03x5               g124(.a(new_n209), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n212), .b(new_n220), .c(new_n194), .d(new_n207), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n218), .c(new_n211), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n219), .b(new_n222), .o1(\s[20] ));
  nor042aa1n03x5               g128(.a(new_n202), .b(new_n200), .o1(new_n224));
  nano23aa1n06x5               g129(.a(new_n216), .b(new_n211), .c(new_n217), .d(new_n210), .out0(new_n225));
  nand02aa1d06x5               g130(.a(new_n225), .b(new_n207), .o1(new_n226));
  nona23aa1n09x5               g131(.a(new_n210), .b(new_n217), .c(new_n216), .d(new_n211), .out0(new_n227));
  aoi012aa1n02x7               g132(.a(new_n216), .b(new_n211), .c(new_n217), .o1(new_n228));
  oai012aa1n06x5               g133(.a(new_n228), .b(new_n227), .c(new_n209), .o1(new_n229));
  oabi12aa1n06x5               g134(.a(new_n229), .b(new_n224), .c(new_n226), .out0(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[21] ), .b(\b[20] ), .out0(new_n233));
  xorc02aa1n02x5               g138(.a(\a[22] ), .b(\b[21] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n226), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n233), .b(new_n229), .c(new_n194), .d(new_n237), .o1(new_n238));
  nona22aa1n02x4               g143(.a(new_n238), .b(new_n235), .c(new_n232), .out0(new_n239));
  nanp02aa1n03x5               g144(.a(new_n236), .b(new_n239), .o1(\s[22] ));
  inv020aa1n03x5               g145(.a(new_n228), .o1(new_n241));
  inv000aa1d42x5               g146(.a(\a[21] ), .o1(new_n242));
  inv040aa1d32x5               g147(.a(\a[22] ), .o1(new_n243));
  xroi22aa1d06x4               g148(.a(new_n242), .b(\b[20] ), .c(new_n243), .d(\b[21] ), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n241), .c(new_n225), .d(new_n220), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\b[21] ), .o1(new_n246));
  oaoi03aa1n12x5               g151(.a(new_n243), .b(new_n246), .c(new_n232), .o1(new_n247));
  nanp02aa1n02x5               g152(.a(new_n245), .b(new_n247), .o1(new_n248));
  inv020aa1d32x5               g153(.a(new_n248), .o1(new_n249));
  oai112aa1n03x5               g154(.a(new_n237), .b(new_n244), .c(new_n202), .d(new_n200), .o1(new_n250));
  xnrc02aa1n12x5               g155(.a(\b[22] ), .b(\a[23] ), .out0(new_n251));
  xobna2aa1n03x5               g156(.a(new_n251), .b(new_n250), .c(new_n249), .out0(\s[23] ));
  and002aa1n02x5               g157(.a(\b[22] ), .b(\a[23] ), .o(new_n253));
  xorc02aa1n12x5               g158(.a(\a[24] ), .b(\b[23] ), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n247), .o1(new_n256));
  norp02aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  aoi112aa1n02x5               g162(.a(new_n257), .b(new_n256), .c(new_n229), .d(new_n244), .o1(new_n258));
  aoai13aa1n02x7               g163(.a(new_n255), .b(new_n253), .c(new_n250), .d(new_n258), .o1(new_n259));
  aoi112aa1n02x7               g164(.a(new_n255), .b(new_n253), .c(new_n250), .d(new_n258), .o1(new_n260));
  norb02aa1n03x4               g165(.a(new_n259), .b(new_n260), .out0(\s[24] ));
  norb02aa1n09x5               g166(.a(new_n254), .b(new_n251), .out0(new_n262));
  inv030aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  nano32aa1n02x4               g168(.a(new_n263), .b(new_n244), .c(new_n225), .d(new_n207), .out0(new_n264));
  oaih12aa1n02x5               g169(.a(new_n264), .b(new_n202), .c(new_n200), .o1(new_n265));
  aoi112aa1n02x5               g170(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n266));
  oab012aa1n02x4               g171(.a(new_n266), .b(\a[24] ), .c(\b[23] ), .out0(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n263), .c(new_n245), .d(new_n247), .o1(new_n268));
  nanb02aa1n03x5               g173(.a(new_n268), .b(new_n265), .out0(new_n269));
  xorb03aa1n02x5               g174(.a(new_n269), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g175(.a(\b[24] ), .b(\a[25] ), .o1(new_n271));
  tech160nm_fixorc02aa1n03p5x5 g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  xorc02aa1n12x5               g177(.a(\a[26] ), .b(\b[25] ), .out0(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n02x5               g179(.a(new_n274), .b(new_n271), .c(new_n269), .d(new_n272), .o1(new_n275));
  aoai13aa1n03x5               g180(.a(new_n272), .b(new_n268), .c(new_n194), .d(new_n264), .o1(new_n276));
  nona22aa1n03x5               g181(.a(new_n276), .b(new_n274), .c(new_n271), .out0(new_n277));
  nanp02aa1n02x5               g182(.a(new_n275), .b(new_n277), .o1(\s[26] ));
  and002aa1n12x5               g183(.a(new_n273), .b(new_n272), .o(new_n279));
  nano32aa1n03x7               g184(.a(new_n226), .b(new_n279), .c(new_n244), .d(new_n262), .out0(new_n280));
  oai012aa1n06x5               g185(.a(new_n280), .b(new_n202), .c(new_n200), .o1(new_n281));
  orn002aa1n02x5               g186(.a(\a[25] ), .b(\b[24] ), .o(new_n282));
  oao003aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .c(new_n282), .carry(new_n283));
  aobi12aa1n06x5               g188(.a(new_n283), .b(new_n268), .c(new_n279), .out0(new_n284));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(\b[26] ), .b(\a[27] ), .o1(new_n286));
  norb02aa1n02x5               g191(.a(new_n286), .b(new_n285), .out0(new_n287));
  xnbna2aa1n03x5               g192(.a(new_n287), .b(new_n284), .c(new_n281), .out0(\s[27] ));
  inv000aa1n06x5               g193(.a(new_n285), .o1(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[27] ), .b(\a[28] ), .out0(new_n290));
  aobi12aa1n02x7               g195(.a(new_n286), .b(new_n284), .c(new_n281), .out0(new_n291));
  nano22aa1n03x5               g196(.a(new_n291), .b(new_n289), .c(new_n290), .out0(new_n292));
  aoai13aa1n04x5               g197(.a(new_n262), .b(new_n256), .c(new_n229), .d(new_n244), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n279), .o1(new_n294));
  aoai13aa1n06x5               g199(.a(new_n283), .b(new_n294), .c(new_n293), .d(new_n267), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n286), .b(new_n295), .c(new_n194), .d(new_n280), .o1(new_n296));
  tech160nm_fiaoi012aa1n02p5x5 g201(.a(new_n290), .b(new_n296), .c(new_n289), .o1(new_n297));
  norp02aa1n03x5               g202(.a(new_n297), .b(new_n292), .o1(\s[28] ));
  nano22aa1n02x4               g203(.a(new_n290), .b(new_n289), .c(new_n286), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n295), .c(new_n194), .d(new_n280), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[28] ), .b(\a[29] ), .out0(new_n302));
  aoi012aa1n02x7               g207(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n303));
  aobi12aa1n02x7               g208(.a(new_n299), .b(new_n284), .c(new_n281), .out0(new_n304));
  nano22aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n302), .out0(new_n305));
  norp02aa1n03x5               g210(.a(new_n303), .b(new_n305), .o1(\s[29] ));
  xorb03aa1n02x5               g211(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g212(.a(new_n287), .b(new_n302), .c(new_n290), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n295), .c(new_n194), .d(new_n280), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .carry(new_n310));
  xnrc02aa1n02x5               g215(.a(\b[29] ), .b(\a[30] ), .out0(new_n311));
  aoi012aa1n03x5               g216(.a(new_n311), .b(new_n309), .c(new_n310), .o1(new_n312));
  aobi12aa1n06x5               g217(.a(new_n308), .b(new_n284), .c(new_n281), .out0(new_n313));
  nano22aa1n03x5               g218(.a(new_n313), .b(new_n310), .c(new_n311), .out0(new_n314));
  nor002aa1n02x5               g219(.a(new_n312), .b(new_n314), .o1(\s[30] ));
  norb03aa1n02x5               g220(.a(new_n299), .b(new_n311), .c(new_n302), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n295), .c(new_n194), .d(new_n280), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n310), .carry(new_n318));
  xnrc02aa1n02x5               g223(.a(\b[30] ), .b(\a[31] ), .out0(new_n319));
  tech160nm_fiaoi012aa1n02p5x5 g224(.a(new_n319), .b(new_n317), .c(new_n318), .o1(new_n320));
  aobi12aa1n02x7               g225(.a(new_n316), .b(new_n284), .c(new_n281), .out0(new_n321));
  nano22aa1n03x5               g226(.a(new_n321), .b(new_n318), .c(new_n319), .out0(new_n322));
  norp02aa1n03x5               g227(.a(new_n320), .b(new_n322), .o1(\s[31] ));
  xnrb03aa1n02x5               g228(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g229(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oao003aa1n03x5               g232(.a(\a[5] ), .b(\b[4] ), .c(new_n135), .carry(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n117), .c(new_n119), .out0(\s[6] ));
  inv000aa1d42x5               g234(.a(new_n137), .o1(new_n330));
  aob012aa1n03x5               g235(.a(new_n119), .b(new_n328), .c(new_n117), .out0(new_n331));
  xnrc02aa1n02x5               g236(.a(new_n331), .b(new_n330), .out0(\s[7] ));
  aoai13aa1n02x5               g237(.a(new_n136), .b(new_n116), .c(new_n331), .d(new_n330), .o1(new_n333));
  aoi112aa1n02x5               g238(.a(new_n136), .b(new_n116), .c(new_n331), .d(new_n330), .o1(new_n334));
  norb02aa1n03x4               g239(.a(new_n333), .b(new_n334), .out0(\s[8] ));
  xorb03aa1n02x5               g240(.a(new_n139), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


