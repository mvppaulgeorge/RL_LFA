// Benchmark "adder" written by ABC on Wed Jul 17 14:43:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n328, new_n329, new_n332, new_n334,
    new_n335, new_n336, new_n338, new_n340;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n06x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  inv040aa1d32x5               g004(.a(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[8] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  and002aa1n12x5               g007(.a(\b[0] ), .b(\a[1] ), .o(new_n103));
  oaoi03aa1n09x5               g008(.a(\a[2] ), .b(\b[1] ), .c(new_n103), .o1(new_n104));
  nor002aa1n03x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nand42aa1n10x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  norb02aa1n03x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  norp02aa1n12x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand42aa1n10x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  norb02aa1d21x5               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  nand23aa1n06x5               g015(.a(new_n104), .b(new_n107), .c(new_n110), .o1(new_n111));
  aoi012aa1n06x5               g016(.a(new_n105), .b(new_n108), .c(new_n106), .o1(new_n112));
  nand42aa1d28x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor042aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor042aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n24x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1d15x5               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  tech160nm_fixorc02aa1n05x5   g022(.a(\a[6] ), .b(\b[5] ), .out0(new_n118));
  xorc02aa1n12x5               g023(.a(\a[5] ), .b(\b[4] ), .out0(new_n119));
  nand23aa1n06x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  nor042aa1d18x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  inv030aa1n06x5               g026(.a(new_n121), .o1(new_n122));
  oaoi03aa1n12x5               g027(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n123));
  oai022aa1n02x5               g028(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n124));
  aoi022aa1n09x5               g029(.a(new_n117), .b(new_n123), .c(new_n113), .d(new_n124), .o1(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n120), .c(new_n111), .d(new_n112), .o1(new_n126));
  xnrc02aa1n12x5               g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(new_n126), .b(new_n128), .o1(new_n129));
  xobna2aa1n03x5               g034(.a(new_n99), .b(new_n129), .c(new_n102), .out0(\s[10] ));
  norp02aa1n02x5               g035(.a(new_n127), .b(new_n99), .o1(new_n131));
  oaoi03aa1n02x5               g036(.a(\a[10] ), .b(\b[9] ), .c(new_n102), .o1(new_n132));
  nor002aa1d24x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1n06x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n133), .b(new_n134), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  aoai13aa1n03x5               g041(.a(new_n136), .b(new_n132), .c(new_n126), .d(new_n131), .o1(new_n137));
  aoi112aa1n02x5               g042(.a(new_n136), .b(new_n132), .c(new_n126), .d(new_n131), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n137), .b(new_n138), .out0(\s[11] ));
  inv020aa1n04x5               g044(.a(new_n133), .o1(new_n140));
  nor022aa1n16x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1n06x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  xobna2aa1n03x5               g048(.a(new_n143), .b(new_n137), .c(new_n140), .out0(\s[12] ));
  nano23aa1n09x5               g049(.a(new_n133), .b(new_n141), .c(new_n142), .d(new_n134), .out0(new_n145));
  nona22aa1n09x5               g050(.a(new_n145), .b(new_n127), .c(new_n99), .out0(new_n146));
  nanb02aa1n06x5               g051(.a(new_n146), .b(new_n126), .out0(new_n147));
  aoai13aa1n06x5               g052(.a(new_n98), .b(new_n97), .c(new_n100), .d(new_n101), .o1(new_n148));
  nona23aa1d18x5               g053(.a(new_n142), .b(new_n134), .c(new_n133), .d(new_n141), .out0(new_n149));
  oaoi03aa1n09x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n140), .o1(new_n150));
  oabi12aa1n18x5               g055(.a(new_n150), .b(new_n149), .c(new_n148), .out0(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nor042aa1n04x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1n08x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(new_n155));
  xobna2aa1n03x5               g060(.a(new_n155), .b(new_n147), .c(new_n152), .out0(\s[13] ));
  nand22aa1n03x5               g061(.a(new_n147), .b(new_n152), .o1(new_n157));
  tech160nm_fiaoi012aa1n05x5   g062(.a(new_n153), .b(new_n157), .c(new_n154), .o1(new_n158));
  xnrb03aa1n03x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n06x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nano23aa1d15x5               g066(.a(new_n153), .b(new_n160), .c(new_n161), .d(new_n154), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  tech160nm_fioai012aa1n04x5   g068(.a(new_n161), .b(new_n160), .c(new_n153), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n163), .c(new_n147), .d(new_n152), .o1(new_n165));
  nor042aa1n06x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nand42aa1n08x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  inv020aa1n02x5               g074(.a(new_n164), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n169), .b(new_n170), .c(new_n157), .d(new_n162), .o1(new_n171));
  aoi012aa1n02x5               g076(.a(new_n171), .b(new_n165), .c(new_n169), .o1(\s[15] ));
  nor002aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand42aa1n08x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n166), .c(new_n165), .d(new_n169), .o1(new_n176));
  nand42aa1n04x5               g081(.a(new_n165), .b(new_n169), .o1(new_n177));
  nona22aa1n02x4               g082(.a(new_n177), .b(new_n175), .c(new_n166), .out0(new_n178));
  nanp02aa1n03x5               g083(.a(new_n178), .b(new_n176), .o1(\s[16] ));
  inv040aa1d32x5               g084(.a(\a[17] ), .o1(new_n180));
  nano23aa1d15x5               g085(.a(new_n166), .b(new_n173), .c(new_n174), .d(new_n167), .out0(new_n181));
  nano22aa1n12x5               g086(.a(new_n146), .b(new_n162), .c(new_n181), .out0(new_n182));
  inv000aa1d42x5               g087(.a(new_n181), .o1(new_n183));
  aoai13aa1n06x5               g088(.a(new_n162), .b(new_n150), .c(new_n145), .d(new_n132), .o1(new_n184));
  aoi012aa1n06x5               g089(.a(new_n183), .b(new_n184), .c(new_n164), .o1(new_n185));
  aoi012aa1n02x7               g090(.a(new_n173), .b(new_n166), .c(new_n174), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n186), .o1(new_n187));
  aoi112aa1n09x5               g092(.a(new_n185), .b(new_n187), .c(new_n126), .d(new_n182), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(new_n180), .out0(\s[17] ));
  inv030aa1n24x5               g094(.a(\b[16] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n190), .b(new_n180), .o1(new_n191));
  aoai13aa1n04x5               g096(.a(new_n186), .b(new_n183), .c(new_n184), .d(new_n164), .o1(new_n192));
  tech160nm_fixorc02aa1n03p5x5 g097(.a(\a[17] ), .b(\b[16] ), .out0(new_n193));
  aoai13aa1n03x5               g098(.a(new_n193), .b(new_n192), .c(new_n126), .d(new_n182), .o1(new_n194));
  norp02aa1n12x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nand02aa1n06x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nanb02aa1n12x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  xobna2aa1n03x5               g102(.a(new_n197), .b(new_n194), .c(new_n191), .out0(\s[18] ));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  xroi22aa1d06x4               g104(.a(new_n180), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n200));
  inv000aa1n02x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n196), .b(new_n195), .c(new_n180), .d(new_n190), .o1(new_n202));
  tech160nm_fioai012aa1n05x5   g107(.a(new_n202), .b(new_n188), .c(new_n201), .o1(new_n203));
  nor002aa1d32x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanp02aa1n04x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  norb02aa1n06x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  nanp02aa1n06x5               g111(.a(new_n126), .b(new_n182), .o1(new_n207));
  aoai13aa1n09x5               g112(.a(new_n181), .b(new_n170), .c(new_n151), .d(new_n162), .o1(new_n208));
  nand23aa1d12x5               g113(.a(new_n207), .b(new_n208), .c(new_n186), .o1(new_n209));
  oaoi03aa1n03x5               g114(.a(\a[18] ), .b(\b[17] ), .c(new_n191), .o1(new_n210));
  aoi112aa1n02x5               g115(.a(new_n206), .b(new_n210), .c(new_n209), .d(new_n200), .o1(new_n211));
  tech160nm_fiaoi012aa1n02p5x5 g116(.a(new_n211), .b(new_n203), .c(new_n206), .o1(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n16x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand22aa1n12x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nanb02aa1n03x5               g120(.a(new_n214), .b(new_n215), .out0(new_n216));
  aoai13aa1n02x7               g121(.a(new_n216), .b(new_n204), .c(new_n203), .d(new_n206), .o1(new_n217));
  aoai13aa1n04x5               g122(.a(new_n206), .b(new_n210), .c(new_n209), .d(new_n200), .o1(new_n218));
  nona22aa1n03x5               g123(.a(new_n218), .b(new_n216), .c(new_n204), .out0(new_n219));
  nanp02aa1n03x5               g124(.a(new_n217), .b(new_n219), .o1(\s[20] ));
  nona23aa1d18x5               g125(.a(new_n206), .b(new_n193), .c(new_n216), .d(new_n197), .out0(new_n221));
  nona23aa1n09x5               g126(.a(new_n215), .b(new_n205), .c(new_n204), .d(new_n214), .out0(new_n222));
  ao0012aa1n03x7               g127(.a(new_n214), .b(new_n204), .c(new_n215), .o(new_n223));
  oabi12aa1n18x5               g128(.a(new_n223), .b(new_n222), .c(new_n202), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  tech160nm_fioai012aa1n04x5   g130(.a(new_n225), .b(new_n188), .c(new_n221), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n221), .o1(new_n229));
  aoi112aa1n03x4               g134(.a(new_n228), .b(new_n224), .c(new_n209), .d(new_n229), .o1(new_n230));
  aoi012aa1n02x5               g135(.a(new_n230), .b(new_n226), .c(new_n228), .o1(\s[21] ));
  nor002aa1n03x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[21] ), .b(\a[22] ), .out0(new_n233));
  aoai13aa1n03x5               g138(.a(new_n233), .b(new_n232), .c(new_n226), .d(new_n228), .o1(new_n234));
  aoai13aa1n04x5               g139(.a(new_n228), .b(new_n224), .c(new_n209), .d(new_n229), .o1(new_n235));
  nona22aa1n03x5               g140(.a(new_n235), .b(new_n233), .c(new_n232), .out0(new_n236));
  nanp02aa1n03x5               g141(.a(new_n234), .b(new_n236), .o1(\s[22] ));
  nano23aa1n03x7               g142(.a(new_n204), .b(new_n214), .c(new_n215), .d(new_n205), .out0(new_n238));
  nor042aa1n06x5               g143(.a(new_n233), .b(new_n227), .o1(new_n239));
  nano22aa1n03x7               g144(.a(new_n201), .b(new_n239), .c(new_n238), .out0(new_n240));
  inv000aa1n02x5               g145(.a(new_n240), .o1(new_n241));
  inv000aa1d42x5               g146(.a(\a[22] ), .o1(new_n242));
  inv000aa1d42x5               g147(.a(\b[21] ), .o1(new_n243));
  oaoi03aa1n12x5               g148(.a(new_n242), .b(new_n243), .c(new_n232), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  aoi012aa1d18x5               g150(.a(new_n245), .b(new_n224), .c(new_n239), .o1(new_n246));
  tech160nm_fioai012aa1n04x5   g151(.a(new_n246), .b(new_n188), .c(new_n241), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[23] ), .b(\b[22] ), .out0(new_n248));
  inv000aa1d42x5               g153(.a(new_n246), .o1(new_n249));
  aoi112aa1n03x4               g154(.a(new_n248), .b(new_n249), .c(new_n209), .d(new_n240), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n250), .b(new_n247), .c(new_n248), .o1(\s[23] ));
  norp02aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  xnrc02aa1n12x5               g157(.a(\b[23] ), .b(\a[24] ), .out0(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n252), .c(new_n247), .d(new_n248), .o1(new_n254));
  aoai13aa1n04x5               g159(.a(new_n248), .b(new_n249), .c(new_n209), .d(new_n240), .o1(new_n255));
  nona22aa1n03x5               g160(.a(new_n255), .b(new_n253), .c(new_n252), .out0(new_n256));
  nanp02aa1n03x5               g161(.a(new_n254), .b(new_n256), .o1(\s[24] ));
  norb02aa1n03x5               g162(.a(new_n248), .b(new_n253), .out0(new_n258));
  inv040aa1n02x5               g163(.a(new_n258), .o1(new_n259));
  nano32aa1n03x7               g164(.a(new_n259), .b(new_n200), .c(new_n239), .d(new_n238), .out0(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  aoai13aa1n06x5               g166(.a(new_n239), .b(new_n223), .c(new_n238), .d(new_n210), .o1(new_n262));
  aoi112aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n263));
  oab012aa1n02x4               g168(.a(new_n263), .b(\a[24] ), .c(\b[23] ), .out0(new_n264));
  aoai13aa1n09x5               g169(.a(new_n264), .b(new_n259), .c(new_n262), .d(new_n244), .o1(new_n265));
  inv000aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  tech160nm_fioai012aa1n05x5   g171(.a(new_n266), .b(new_n188), .c(new_n261), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  tech160nm_fixorc02aa1n05x5   g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xnrc02aa1n12x5               g175(.a(\b[25] ), .b(\a[26] ), .out0(new_n271));
  aoai13aa1n02x7               g176(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n270), .o1(new_n272));
  aoai13aa1n04x5               g177(.a(new_n270), .b(new_n265), .c(new_n209), .d(new_n260), .o1(new_n273));
  nona22aa1n03x5               g178(.a(new_n273), .b(new_n271), .c(new_n269), .out0(new_n274));
  nanp02aa1n03x5               g179(.a(new_n272), .b(new_n274), .o1(\s[26] ));
  norb02aa1n06x5               g180(.a(new_n270), .b(new_n271), .out0(new_n276));
  nano23aa1n06x5               g181(.a(new_n221), .b(new_n259), .c(new_n276), .d(new_n239), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n192), .c(new_n126), .d(new_n182), .o1(new_n278));
  inv020aa1n02x5               g183(.a(new_n277), .o1(new_n279));
  inv000aa1d42x5               g184(.a(\a[26] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(\b[25] ), .o1(new_n281));
  tech160nm_fioaoi03aa1n03p5x5 g186(.a(new_n280), .b(new_n281), .c(new_n269), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  aoi012aa1n09x5               g188(.a(new_n283), .b(new_n265), .c(new_n276), .o1(new_n284));
  tech160nm_fioai012aa1n05x5   g189(.a(new_n284), .b(new_n188), .c(new_n279), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  aoi112aa1n02x5               g191(.a(new_n286), .b(new_n283), .c(new_n265), .d(new_n276), .o1(new_n287));
  aoi022aa1n03x5               g192(.a(new_n285), .b(new_n286), .c(new_n278), .d(new_n287), .o1(\s[27] ));
  norp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  nor002aa1n03x5               g194(.a(\b[27] ), .b(\a[28] ), .o1(new_n290));
  nand02aa1n06x5               g195(.a(\b[27] ), .b(\a[28] ), .o1(new_n291));
  nanb02aa1n06x5               g196(.a(new_n290), .b(new_n291), .out0(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n289), .c(new_n285), .d(new_n286), .o1(new_n293));
  aoai13aa1n09x5               g198(.a(new_n258), .b(new_n245), .c(new_n224), .d(new_n239), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n276), .o1(new_n295));
  aoai13aa1n04x5               g200(.a(new_n282), .b(new_n295), .c(new_n294), .d(new_n264), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n286), .b(new_n296), .c(new_n209), .d(new_n277), .o1(new_n297));
  nona22aa1n02x4               g202(.a(new_n297), .b(new_n292), .c(new_n289), .out0(new_n298));
  nanp02aa1n03x5               g203(.a(new_n293), .b(new_n298), .o1(\s[28] ));
  norb02aa1n03x5               g204(.a(new_n286), .b(new_n292), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n209), .d(new_n277), .o1(new_n301));
  norp02aa1n02x5               g206(.a(\b[28] ), .b(\a[29] ), .o1(new_n302));
  nand42aa1n03x5               g207(.a(\b[28] ), .b(\a[29] ), .o1(new_n303));
  norb02aa1n02x5               g208(.a(new_n303), .b(new_n302), .out0(new_n304));
  oai022aa1n02x5               g209(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n305));
  aboi22aa1n03x5               g210(.a(new_n302), .b(new_n303), .c(new_n305), .d(new_n291), .out0(new_n306));
  inv000aa1d42x5               g211(.a(new_n300), .o1(new_n307));
  oai012aa1n02x5               g212(.a(new_n291), .b(new_n290), .c(new_n289), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n307), .c(new_n278), .d(new_n284), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n309), .b(new_n304), .c(new_n301), .d(new_n306), .o1(\s[29] ));
  xnrb03aa1n02x5               g215(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g216(.a(new_n292), .b(new_n286), .c(new_n304), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n296), .c(new_n209), .d(new_n277), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .out0(new_n314));
  aoi113aa1n02x5               g219(.a(new_n314), .b(new_n302), .c(new_n303), .d(new_n305), .e(new_n291), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n312), .o1(new_n316));
  aoi013aa1n02x4               g221(.a(new_n302), .b(new_n305), .c(new_n303), .d(new_n291), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n316), .c(new_n278), .d(new_n284), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n313), .d(new_n315), .o1(\s[30] ));
  nand03aa1n02x5               g224(.a(new_n300), .b(new_n304), .c(new_n314), .o1(new_n320));
  nanb02aa1n03x5               g225(.a(new_n320), .b(new_n285), .out0(new_n321));
  xorc02aa1n02x5               g226(.a(\a[31] ), .b(\b[30] ), .out0(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n323));
  norb02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(new_n324));
  aoai13aa1n02x7               g229(.a(new_n323), .b(new_n320), .c(new_n278), .d(new_n284), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n325), .b(new_n322), .c(new_n321), .d(new_n324), .o1(\s[31] ));
  xorb03aa1n02x5               g231(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g232(.a(new_n111), .b(new_n112), .o1(new_n328));
  aoi112aa1n02x5               g233(.a(new_n108), .b(new_n107), .c(new_n104), .d(new_n109), .o1(new_n329));
  oaoi13aa1n02x5               g234(.a(new_n329), .b(new_n328), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g235(.a(new_n119), .b(new_n111), .c(new_n112), .out0(\s[5] ));
  nanp02aa1n02x5               g236(.a(new_n328), .b(new_n119), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n118), .b(new_n332), .c(new_n122), .out0(\s[6] ));
  nanb02aa1n02x5               g238(.a(new_n115), .b(new_n116), .out0(new_n334));
  nanp02aa1n02x5               g239(.a(\b[5] ), .b(\a[6] ), .o1(new_n335));
  nanp03aa1n02x5               g240(.a(new_n332), .b(new_n118), .c(new_n122), .o1(new_n336));
  xnbna2aa1n03x5               g241(.a(new_n334), .b(new_n336), .c(new_n335), .out0(\s[7] ));
  aoi013aa1n02x4               g242(.a(new_n115), .b(new_n336), .c(new_n335), .d(new_n116), .o1(new_n338));
  xnrb03aa1n02x5               g243(.a(new_n338), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  nanb02aa1n02x5               g244(.a(new_n120), .b(new_n328), .out0(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n128), .b(new_n340), .c(new_n125), .out0(\s[9] ));
endmodule


