// Benchmark "adder" written by ABC on Thu Jul 18 10:21:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n318, new_n320, new_n321, new_n324, new_n325, new_n327,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand22aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  norp02aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[1] ), .o1(new_n102));
  nand42aa1n03x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  oao003aa1n02x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .carry(new_n104));
  xorc02aa1n02x5               g009(.a(\a[4] ), .b(\b[3] ), .out0(new_n105));
  xorc02aa1n02x5               g010(.a(\a[3] ), .b(\b[2] ), .out0(new_n106));
  nanp03aa1n02x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  orn002aa1n02x5               g012(.a(\a[4] ), .b(\b[3] ), .o(new_n108));
  aoi112aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n109));
  norb02aa1n06x4               g014(.a(new_n108), .b(new_n109), .out0(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .out0(new_n111));
  tech160nm_fixorc02aa1n03p5x5 g016(.a(\a[5] ), .b(\b[4] ), .out0(new_n112));
  xorc02aa1n12x5               g017(.a(\a[8] ), .b(\b[7] ), .out0(new_n113));
  nor002aa1d32x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanb02aa1n06x5               g020(.a(new_n114), .b(new_n115), .out0(new_n116));
  nona23aa1n09x5               g021(.a(new_n112), .b(new_n113), .c(new_n111), .d(new_n116), .out0(new_n117));
  nanp02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nano22aa1n09x5               g023(.a(new_n114), .b(new_n118), .c(new_n115), .out0(new_n119));
  oai022aa1n06x5               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n114), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[8] ), .b(\b[7] ), .c(new_n121), .o1(new_n122));
  aoi013aa1n09x5               g027(.a(new_n122), .b(new_n119), .c(new_n113), .d(new_n120), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n123), .b(new_n117), .c(new_n107), .d(new_n110), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n99), .b(new_n100), .c(new_n124), .d(new_n125), .o1(new_n126));
  oaoi03aa1n02x5               g031(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n127));
  xnrc02aa1n02x5               g032(.a(\b[3] ), .b(\a[4] ), .out0(new_n128));
  xnrc02aa1n02x5               g033(.a(\b[2] ), .b(\a[3] ), .out0(new_n129));
  oai013aa1n02x4               g034(.a(new_n110), .b(new_n127), .c(new_n128), .d(new_n129), .o1(new_n130));
  xorc02aa1n02x5               g035(.a(\a[6] ), .b(\b[5] ), .out0(new_n131));
  nano32aa1n02x5               g036(.a(new_n116), .b(new_n113), .c(new_n112), .d(new_n131), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n123), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n125), .b(new_n133), .c(new_n132), .d(new_n130), .o1(new_n134));
  norb03aa1n02x5               g039(.a(new_n98), .b(new_n97), .c(new_n100), .out0(new_n135));
  nand42aa1n03x5               g040(.a(new_n134), .b(new_n135), .o1(new_n136));
  nanp02aa1n02x5               g041(.a(new_n126), .b(new_n136), .o1(\s[10] ));
  nanp02aa1n02x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  inv000aa1d42x5               g043(.a(\a[11] ), .o1(new_n139));
  inv000aa1d42x5               g044(.a(\b[10] ), .o1(new_n140));
  nand42aa1n03x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  nanp03aa1n02x5               g046(.a(new_n141), .b(new_n98), .c(new_n138), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n142), .b(new_n136), .out0(new_n143));
  aoi022aa1n02x5               g048(.a(new_n136), .b(new_n98), .c(new_n141), .d(new_n138), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(\s[11] ));
  tech160nm_fixorc02aa1n03p5x5 g050(.a(\a[12] ), .b(\b[11] ), .out0(new_n146));
  orn002aa1n02x5               g051(.a(\a[12] ), .b(\b[11] ), .o(new_n147));
  and002aa1n02x5               g052(.a(\b[11] ), .b(\a[12] ), .o(new_n148));
  aboi22aa1n03x5               g053(.a(new_n148), .b(new_n147), .c(new_n140), .d(new_n139), .out0(new_n149));
  aoai13aa1n02x5               g054(.a(new_n141), .b(new_n142), .c(new_n134), .d(new_n135), .o1(new_n150));
  aoi022aa1n02x5               g055(.a(new_n143), .b(new_n149), .c(new_n150), .d(new_n146), .o1(\s[12] ));
  nanp02aa1n03x5               g056(.a(new_n141), .b(new_n138), .o1(new_n152));
  nona23aa1d18x5               g057(.a(new_n146), .b(new_n125), .c(new_n99), .d(new_n152), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n133), .c(new_n132), .d(new_n130), .o1(new_n155));
  aoai13aa1n02x5               g060(.a(new_n138), .b(new_n97), .c(new_n100), .d(new_n98), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n147), .b(new_n148), .c(new_n156), .d(new_n141), .o1(new_n157));
  nanb02aa1n02x5               g062(.a(new_n157), .b(new_n155), .out0(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g064(.a(\a[13] ), .o1(new_n160));
  nanb02aa1d24x5               g065(.a(\b[12] ), .b(new_n160), .out0(new_n161));
  xorc02aa1n02x5               g066(.a(\a[13] ), .b(\b[12] ), .out0(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n157), .c(new_n124), .d(new_n154), .o1(new_n163));
  xorc02aa1n02x5               g068(.a(\a[14] ), .b(\b[13] ), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n163), .c(new_n161), .out0(\s[14] ));
  inv000aa1d42x5               g070(.a(\a[14] ), .o1(new_n166));
  xroi22aa1d04x5               g071(.a(new_n160), .b(\b[12] ), .c(new_n166), .d(\b[13] ), .out0(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n157), .c(new_n124), .d(new_n154), .o1(new_n168));
  oaoi03aa1n09x5               g073(.a(\a[14] ), .b(\b[13] ), .c(new_n161), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  xorc02aa1n12x5               g075(.a(\a[15] ), .b(\b[14] ), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n168), .c(new_n170), .out0(\s[15] ));
  aoai13aa1n02x5               g077(.a(new_n171), .b(new_n169), .c(new_n158), .d(new_n167), .o1(new_n173));
  tech160nm_fixorc02aa1n04x5   g078(.a(\a[16] ), .b(\b[15] ), .out0(new_n174));
  nor042aa1n03x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  norp02aa1n02x5               g080(.a(new_n174), .b(new_n175), .o1(new_n176));
  inv000aa1d42x5               g081(.a(new_n175), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n171), .o1(new_n178));
  aoai13aa1n02x5               g083(.a(new_n177), .b(new_n178), .c(new_n168), .d(new_n170), .o1(new_n179));
  aoi022aa1n02x5               g084(.a(new_n179), .b(new_n174), .c(new_n173), .d(new_n176), .o1(\s[16] ));
  nanp02aa1n02x5               g085(.a(new_n164), .b(new_n162), .o1(new_n181));
  nanp02aa1n06x5               g086(.a(new_n174), .b(new_n171), .o1(new_n182));
  nor043aa1n06x5               g087(.a(new_n153), .b(new_n181), .c(new_n182), .o1(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n133), .c(new_n132), .d(new_n130), .o1(new_n184));
  nano22aa1n02x4               g089(.a(new_n182), .b(new_n162), .c(new_n164), .out0(new_n185));
  nanp02aa1n03x5               g090(.a(new_n185), .b(new_n157), .o1(new_n186));
  oaoi03aa1n02x5               g091(.a(\a[16] ), .b(\b[15] ), .c(new_n177), .o1(new_n187));
  aoi013aa1n06x4               g092(.a(new_n187), .b(new_n169), .c(new_n171), .d(new_n174), .o1(new_n188));
  nanp02aa1n09x5               g093(.a(new_n186), .b(new_n188), .o1(new_n189));
  nanb02aa1n06x5               g094(.a(new_n189), .b(new_n184), .out0(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(\b[16] ), .b(new_n192), .out0(new_n193));
  xorc02aa1n02x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n194), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n195));
  xorc02aa1n02x5               g100(.a(\a[18] ), .b(\b[17] ), .out0(new_n196));
  xnbna2aa1n03x5               g101(.a(new_n196), .b(new_n195), .c(new_n193), .out0(\s[18] ));
  inv000aa1d42x5               g102(.a(\a[18] ), .o1(new_n198));
  xroi22aa1d04x5               g103(.a(new_n192), .b(\b[16] ), .c(new_n198), .d(\b[17] ), .out0(new_n199));
  aoai13aa1n02x5               g104(.a(new_n199), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n200));
  oai022aa1n02x5               g105(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n201));
  oaib12aa1n06x5               g106(.a(new_n201), .b(new_n198), .c(\b[17] ), .out0(new_n202));
  nor042aa1n06x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand42aa1n02x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n200), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n209));
  aoai13aa1n02x5               g114(.a(new_n206), .b(new_n209), .c(new_n190), .d(new_n199), .o1(new_n210));
  nor042aa1n02x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nand02aa1n03x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  aoib12aa1n02x5               g118(.a(new_n203), .b(new_n212), .c(new_n211), .out0(new_n214));
  inv000aa1n02x5               g119(.a(new_n203), .o1(new_n215));
  aoai13aa1n02x5               g120(.a(new_n215), .b(new_n205), .c(new_n200), .d(new_n202), .o1(new_n216));
  aoi022aa1n02x5               g121(.a(new_n216), .b(new_n213), .c(new_n210), .d(new_n214), .o1(\s[20] ));
  nano23aa1n06x5               g122(.a(new_n203), .b(new_n211), .c(new_n212), .d(new_n204), .out0(new_n218));
  nand23aa1n06x5               g123(.a(new_n218), .b(new_n194), .c(new_n196), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n02x5               g125(.a(new_n220), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n221));
  nona23aa1n09x5               g126(.a(new_n212), .b(new_n204), .c(new_n203), .d(new_n211), .out0(new_n222));
  oaoi03aa1n02x5               g127(.a(\a[20] ), .b(\b[19] ), .c(new_n215), .o1(new_n223));
  oabi12aa1n18x5               g128(.a(new_n223), .b(new_n222), .c(new_n202), .out0(new_n224));
  inv000aa1d42x5               g129(.a(new_n224), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  xnbna2aa1n03x5               g132(.a(new_n227), .b(new_n221), .c(new_n225), .out0(\s[21] ));
  aoai13aa1n02x5               g133(.a(new_n227), .b(new_n224), .c(new_n190), .d(new_n220), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[21] ), .b(\a[22] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  nor042aa1n06x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n230), .b(new_n232), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n232), .o1(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n226), .c(new_n221), .d(new_n225), .o1(new_n235));
  aoi022aa1n02x5               g140(.a(new_n235), .b(new_n231), .c(new_n229), .d(new_n233), .o1(\s[22] ));
  nor042aa1n06x5               g141(.a(new_n230), .b(new_n226), .o1(new_n237));
  norb02aa1n02x7               g142(.a(new_n237), .b(new_n219), .out0(new_n238));
  aoai13aa1n04x5               g143(.a(new_n238), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n239));
  oao003aa1n12x5               g144(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .carry(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoi012aa1n02x5               g146(.a(new_n241), .b(new_n224), .c(new_n237), .o1(new_n242));
  xorc02aa1n12x5               g147(.a(\a[23] ), .b(\b[22] ), .out0(new_n243));
  aob012aa1n06x5               g148(.a(new_n243), .b(new_n239), .c(new_n242), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n237), .b(new_n223), .c(new_n218), .d(new_n209), .o1(new_n245));
  nano32aa1n02x4               g150(.a(new_n243), .b(new_n239), .c(new_n245), .d(new_n240), .out0(new_n246));
  norb02aa1n02x5               g151(.a(new_n244), .b(new_n246), .out0(\s[23] ));
  xorc02aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .out0(new_n248));
  nor042aa1n03x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  norp02aa1n02x5               g154(.a(new_n248), .b(new_n249), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n249), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n243), .o1(new_n252));
  aoai13aa1n02x5               g157(.a(new_n251), .b(new_n252), .c(new_n239), .d(new_n242), .o1(new_n253));
  aoi022aa1n02x5               g158(.a(new_n253), .b(new_n248), .c(new_n244), .d(new_n250), .o1(\s[24] ));
  nano32aa1n06x5               g159(.a(new_n219), .b(new_n248), .c(new_n237), .d(new_n243), .out0(new_n255));
  aoai13aa1n02x5               g160(.a(new_n255), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n256));
  and002aa1n06x5               g161(.a(new_n248), .b(new_n243), .o(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  oao003aa1n02x5               g163(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .carry(new_n259));
  aoai13aa1n12x5               g164(.a(new_n259), .b(new_n258), .c(new_n245), .d(new_n240), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  xorc02aa1n12x5               g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xnbna2aa1n03x5               g167(.a(new_n262), .b(new_n256), .c(new_n261), .out0(\s[25] ));
  aoai13aa1n02x5               g168(.a(new_n262), .b(new_n260), .c(new_n190), .d(new_n255), .o1(new_n264));
  xorc02aa1n02x5               g169(.a(\a[26] ), .b(\b[25] ), .out0(new_n265));
  nor042aa1n03x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  norp02aa1n02x5               g171(.a(new_n265), .b(new_n266), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n266), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n262), .o1(new_n269));
  aoai13aa1n02x5               g174(.a(new_n268), .b(new_n269), .c(new_n256), .d(new_n261), .o1(new_n270));
  aoi022aa1n03x5               g175(.a(new_n270), .b(new_n265), .c(new_n264), .d(new_n267), .o1(\s[26] ));
  and002aa1n02x5               g176(.a(new_n265), .b(new_n262), .o(new_n272));
  inv000aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  nano23aa1n06x5               g178(.a(new_n273), .b(new_n219), .c(new_n257), .d(new_n237), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n189), .c(new_n124), .d(new_n183), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[26] ), .b(\b[25] ), .c(new_n268), .carry(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoi012aa1n12x5               g182(.a(new_n277), .b(new_n260), .c(new_n272), .o1(new_n278));
  xorc02aa1n12x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  xnbna2aa1n03x5               g184(.a(new_n279), .b(new_n278), .c(new_n275), .out0(\s[27] ));
  aoai13aa1n04x5               g185(.a(new_n257), .b(new_n241), .c(new_n224), .d(new_n237), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n276), .b(new_n273), .c(new_n281), .d(new_n259), .o1(new_n282));
  aoai13aa1n02x5               g187(.a(new_n279), .b(new_n282), .c(new_n190), .d(new_n274), .o1(new_n283));
  xorc02aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .out0(new_n284));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  norp02aa1n02x5               g190(.a(new_n284), .b(new_n285), .o1(new_n286));
  inv000aa1n03x5               g191(.a(new_n285), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n279), .o1(new_n288));
  aoai13aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n278), .d(new_n275), .o1(new_n289));
  aoi022aa1n03x5               g194(.a(new_n289), .b(new_n284), .c(new_n283), .d(new_n286), .o1(\s[28] ));
  and002aa1n02x5               g195(.a(new_n284), .b(new_n279), .o(new_n291));
  aoai13aa1n02x5               g196(.a(new_n291), .b(new_n282), .c(new_n190), .d(new_n274), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n291), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .carry(new_n294));
  aoai13aa1n02x5               g199(.a(new_n294), .b(new_n293), .c(new_n278), .d(new_n275), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[29] ), .b(\b[28] ), .out0(new_n296));
  norb02aa1n02x5               g201(.a(new_n294), .b(new_n296), .out0(new_n297));
  aoi022aa1n03x5               g202(.a(new_n295), .b(new_n296), .c(new_n292), .d(new_n297), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g204(.a(new_n288), .b(new_n284), .c(new_n296), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n282), .c(new_n190), .d(new_n274), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n300), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n302), .c(new_n278), .d(new_n275), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n303), .b(new_n305), .out0(new_n306));
  aoi022aa1n02x5               g211(.a(new_n304), .b(new_n305), .c(new_n301), .d(new_n306), .o1(\s[30] ));
  nano32aa1n03x7               g212(.a(new_n288), .b(new_n305), .c(new_n284), .d(new_n296), .out0(new_n308));
  aoai13aa1n02x5               g213(.a(new_n308), .b(new_n282), .c(new_n190), .d(new_n274), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[31] ), .b(\b[30] ), .out0(new_n310));
  and002aa1n02x5               g215(.a(\b[29] ), .b(\a[30] ), .o(new_n311));
  oabi12aa1n02x5               g216(.a(new_n310), .b(\a[30] ), .c(\b[29] ), .out0(new_n312));
  oab012aa1n02x4               g217(.a(new_n312), .b(new_n303), .c(new_n311), .out0(new_n313));
  inv000aa1d42x5               g218(.a(new_n308), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n303), .carry(new_n315));
  aoai13aa1n02x5               g220(.a(new_n315), .b(new_n314), .c(new_n278), .d(new_n275), .o1(new_n316));
  aoi022aa1n03x5               g221(.a(new_n316), .b(new_n310), .c(new_n309), .d(new_n313), .o1(\s[31] ));
  inv000aa1d42x5               g222(.a(\a[3] ), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n127), .b(\b[2] ), .c(new_n318), .out0(\s[3] ));
  nanp02aa1n02x5               g224(.a(new_n104), .b(new_n106), .o1(new_n320));
  aoib12aa1n02x5               g225(.a(new_n105), .b(new_n318), .c(\b[2] ), .out0(new_n321));
  aoi022aa1n02x5               g226(.a(new_n130), .b(new_n108), .c(new_n321), .d(new_n320), .o1(\s[4] ));
  xnbna2aa1n03x5               g227(.a(new_n112), .b(new_n107), .c(new_n110), .out0(\s[5] ));
  norp02aa1n02x5               g228(.a(\b[4] ), .b(\a[5] ), .o1(new_n324));
  aoi012aa1n02x5               g229(.a(new_n324), .b(new_n130), .c(new_n112), .o1(new_n325));
  xnrc02aa1n02x5               g230(.a(new_n325), .b(new_n131), .out0(\s[6] ));
  nanp02aa1n02x5               g231(.a(new_n325), .b(new_n131), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n116), .b(new_n327), .c(new_n118), .out0(\s[7] ));
  nanp02aa1n02x5               g233(.a(new_n327), .b(new_n119), .o1(new_n329));
  xnbna2aa1n03x5               g234(.a(new_n113), .b(new_n329), .c(new_n121), .out0(\s[8] ));
  xorb03aa1n02x5               g235(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


