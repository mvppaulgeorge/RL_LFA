// Benchmark "adder" written by ABC on Thu Jul 18 11:17:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n351, new_n352,
    new_n354, new_n356, new_n357, new_n358, new_n360, new_n361, new_n362,
    new_n364, new_n365, new_n366, new_n368, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  nand02aa1d24x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  inv040aa1n06x5               g004(.a(new_n99), .o1(new_n100));
  oaoi03aa1n09x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand42aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n06x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nor042aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n09x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n06x4               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  nand23aa1n06x5               g012(.a(new_n101), .b(new_n104), .c(new_n107), .o1(new_n108));
  tech160nm_fiaoi012aa1n05x5   g013(.a(new_n102), .b(new_n105), .c(new_n103), .o1(new_n109));
  nor042aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nor002aa1d24x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nano23aa1n06x5               g018(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n114));
  nanp02aa1n04x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor002aa1d32x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  norb02aa1n03x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  nor002aa1n03x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand02aa1d06x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  norb02aa1n03x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  nand23aa1n06x5               g025(.a(new_n114), .b(new_n117), .c(new_n120), .o1(new_n121));
  nano22aa1n12x5               g026(.a(new_n110), .b(new_n111), .c(new_n119), .out0(new_n122));
  oai012aa1n02x5               g027(.a(new_n115), .b(\b[7] ), .c(\a[8] ), .o1(new_n123));
  oab012aa1n03x5               g028(.a(new_n123), .b(new_n112), .c(new_n116), .out0(new_n124));
  tech160nm_fiaoi012aa1n05x5   g029(.a(new_n118), .b(new_n110), .c(new_n119), .o1(new_n125));
  inv000aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  aoi012aa1n06x5               g031(.a(new_n126), .b(new_n124), .c(new_n122), .o1(new_n127));
  aoai13aa1n12x5               g032(.a(new_n127), .b(new_n121), .c(new_n108), .d(new_n109), .o1(new_n128));
  tech160nm_fixorc02aa1n03p5x5 g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  nanp02aa1n02x5               g034(.a(new_n128), .b(new_n129), .o1(new_n130));
  tech160nm_fixorc02aa1n03p5x5 g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  oa0022aa1n03x5               g037(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n133));
  nanp02aa1n02x5               g038(.a(new_n130), .b(new_n133), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nand42aa1n03x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nor042aa1n06x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanb03aa1n02x5               g042(.a(new_n137), .b(new_n135), .c(new_n136), .out0(new_n138));
  nanb02aa1n02x5               g043(.a(new_n138), .b(new_n134), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n137), .o1(new_n140));
  aoi022aa1n02x5               g045(.a(new_n134), .b(new_n135), .c(new_n140), .d(new_n136), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n139), .b(new_n141), .out0(\s[11] ));
  nor042aa1n03x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  aoib12aa1n02x5               g050(.a(new_n137), .b(new_n144), .c(new_n143), .out0(new_n146));
  aoai13aa1n02x5               g051(.a(new_n140), .b(new_n138), .c(new_n130), .d(new_n133), .o1(new_n147));
  aoi022aa1n02x5               g052(.a(new_n139), .b(new_n146), .c(new_n147), .d(new_n145), .o1(\s[12] ));
  nano23aa1n03x7               g053(.a(new_n143), .b(new_n137), .c(new_n144), .d(new_n136), .out0(new_n149));
  and003aa1n02x5               g054(.a(new_n149), .b(new_n131), .c(new_n129), .o(new_n150));
  nanp02aa1n02x5               g055(.a(new_n128), .b(new_n150), .o1(new_n151));
  nano22aa1n03x5               g056(.a(new_n143), .b(new_n136), .c(new_n144), .out0(new_n152));
  nona23aa1n06x5               g057(.a(new_n152), .b(new_n135), .c(new_n133), .d(new_n137), .out0(new_n153));
  aoi012aa1n03x5               g058(.a(new_n143), .b(new_n137), .c(new_n144), .o1(new_n154));
  nand42aa1n04x5               g059(.a(new_n153), .b(new_n154), .o1(new_n155));
  nanb02aa1n02x5               g060(.a(new_n155), .b(new_n151), .out0(new_n156));
  xorc02aa1n12x5               g061(.a(\a[13] ), .b(\b[12] ), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  and003aa1n02x5               g063(.a(new_n153), .b(new_n158), .c(new_n154), .o(new_n159));
  aoi022aa1n02x5               g064(.a(new_n156), .b(new_n157), .c(new_n151), .d(new_n159), .o1(\s[13] ));
  orn002aa1n02x5               g065(.a(\a[13] ), .b(\b[12] ), .o(new_n161));
  aoai13aa1n02x5               g066(.a(new_n157), .b(new_n155), .c(new_n128), .d(new_n150), .o1(new_n162));
  xorc02aa1n06x5               g067(.a(\a[14] ), .b(\b[13] ), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n162), .c(new_n161), .out0(\s[14] ));
  and002aa1n02x5               g069(.a(new_n163), .b(new_n157), .o(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n155), .c(new_n128), .d(new_n150), .o1(new_n166));
  oaoi03aa1n02x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n161), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  nor042aa1n09x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand42aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  norb02aa1n06x4               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n166), .c(new_n168), .out0(\s[15] ));
  aob012aa1n03x5               g077(.a(new_n171), .b(new_n166), .c(new_n168), .out0(new_n173));
  nor002aa1n04x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  norp02aa1n02x5               g081(.a(new_n176), .b(new_n169), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n169), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n171), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n178), .b(new_n179), .c(new_n166), .d(new_n168), .o1(new_n180));
  aoi022aa1n03x5               g085(.a(new_n180), .b(new_n176), .c(new_n173), .d(new_n177), .o1(\s[16] ));
  nano23aa1n06x5               g086(.a(new_n169), .b(new_n174), .c(new_n175), .d(new_n170), .out0(new_n182));
  nand23aa1n06x5               g087(.a(new_n182), .b(new_n157), .c(new_n163), .o1(new_n183));
  nano32aa1n09x5               g088(.a(new_n183), .b(new_n149), .c(new_n131), .d(new_n129), .out0(new_n184));
  nanp02aa1n09x5               g089(.a(new_n128), .b(new_n184), .o1(new_n185));
  inv000aa1n02x5               g090(.a(new_n183), .o1(new_n186));
  nanb03aa1n02x5               g091(.a(new_n174), .b(new_n175), .c(new_n170), .out0(new_n187));
  inv000aa1d42x5               g092(.a(\a[14] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[13] ), .o1(new_n189));
  oaih22aa1n04x5               g094(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n190));
  oai122aa1n02x7               g095(.a(new_n190), .b(\a[15] ), .c(\b[14] ), .d(new_n188), .e(new_n189), .o1(new_n191));
  aoi012aa1n02x5               g096(.a(new_n174), .b(new_n169), .c(new_n175), .o1(new_n192));
  oa0012aa1n06x5               g097(.a(new_n192), .b(new_n191), .c(new_n187), .o(new_n193));
  aobi12aa1n12x5               g098(.a(new_n193), .b(new_n155), .c(new_n186), .out0(new_n194));
  nand22aa1n12x5               g099(.a(new_n185), .b(new_n194), .o1(new_n195));
  xorc02aa1n12x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  norb02aa1n02x5               g101(.a(new_n192), .b(new_n196), .out0(new_n197));
  oai012aa1n02x5               g102(.a(new_n197), .b(new_n191), .c(new_n187), .o1(new_n198));
  aoi012aa1n02x5               g103(.a(new_n198), .b(new_n155), .c(new_n186), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n195), .b(new_n196), .c(new_n185), .d(new_n199), .o1(\s[17] ));
  nor002aa1d32x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n193), .b(new_n183), .c(new_n153), .d(new_n154), .o1(new_n203));
  aoai13aa1n02x5               g108(.a(new_n196), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n204));
  nor002aa1n12x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nand22aa1n09x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  norb02aa1n09x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n204), .c(new_n202), .out0(\s[18] ));
  and002aa1n02x5               g113(.a(new_n196), .b(new_n207), .o(new_n209));
  aoai13aa1n03x5               g114(.a(new_n209), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n210));
  oaoi03aa1n02x5               g115(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor042aa1d18x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand02aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n03x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n210), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n06x5               g122(.a(new_n215), .b(new_n211), .c(new_n195), .d(new_n209), .o1(new_n218));
  nor042aa1n12x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand02aa1d24x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  norb02aa1n06x4               g125(.a(new_n220), .b(new_n219), .out0(new_n221));
  inv000aa1d42x5               g126(.a(\a[19] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(\b[18] ), .o1(new_n223));
  aboi22aa1n03x5               g128(.a(new_n219), .b(new_n220), .c(new_n222), .d(new_n223), .out0(new_n224));
  inv040aa1n02x5               g129(.a(new_n213), .o1(new_n225));
  inv000aa1n02x5               g130(.a(new_n215), .o1(new_n226));
  aoai13aa1n02x5               g131(.a(new_n225), .b(new_n226), .c(new_n210), .d(new_n212), .o1(new_n227));
  aoi022aa1n03x5               g132(.a(new_n227), .b(new_n221), .c(new_n218), .d(new_n224), .o1(\s[20] ));
  nano32aa1n03x7               g133(.a(new_n226), .b(new_n196), .c(new_n221), .d(new_n207), .out0(new_n229));
  aoai13aa1n02x5               g134(.a(new_n229), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n230));
  nanb03aa1n12x5               g135(.a(new_n219), .b(new_n220), .c(new_n214), .out0(new_n231));
  oai112aa1n06x5               g136(.a(new_n225), .b(new_n206), .c(new_n205), .d(new_n201), .o1(new_n232));
  aoi012aa1n12x5               g137(.a(new_n219), .b(new_n213), .c(new_n220), .o1(new_n233));
  oaih12aa1n12x5               g138(.a(new_n233), .b(new_n232), .c(new_n231), .o1(new_n234));
  nor042aa1d18x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nand42aa1d28x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n12x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n234), .c(new_n195), .d(new_n229), .o1(new_n238));
  nano22aa1n03x5               g143(.a(new_n219), .b(new_n214), .c(new_n220), .out0(new_n239));
  oaih12aa1n02x5               g144(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .o1(new_n240));
  oab012aa1n03x5               g145(.a(new_n240), .b(new_n201), .c(new_n205), .out0(new_n241));
  inv020aa1n03x5               g146(.a(new_n233), .o1(new_n242));
  aoi112aa1n02x5               g147(.a(new_n242), .b(new_n237), .c(new_n241), .d(new_n239), .o1(new_n243));
  aobi12aa1n03x7               g148(.a(new_n238), .b(new_n243), .c(new_n230), .out0(\s[21] ));
  nor042aa1n06x5               g149(.a(\b[21] ), .b(\a[22] ), .o1(new_n245));
  nand02aa1d24x5               g150(.a(\b[21] ), .b(\a[22] ), .o1(new_n246));
  norb02aa1n02x7               g151(.a(new_n246), .b(new_n245), .out0(new_n247));
  aoib12aa1n02x5               g152(.a(new_n235), .b(new_n246), .c(new_n245), .out0(new_n248));
  inv000aa1d42x5               g153(.a(new_n234), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n235), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n237), .o1(new_n251));
  aoai13aa1n03x5               g156(.a(new_n250), .b(new_n251), .c(new_n230), .d(new_n249), .o1(new_n252));
  aoi022aa1n03x5               g157(.a(new_n252), .b(new_n247), .c(new_n238), .d(new_n248), .o1(\s[22] ));
  nano23aa1d15x5               g158(.a(new_n235), .b(new_n245), .c(new_n246), .d(new_n236), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  nano32aa1n02x5               g160(.a(new_n255), .b(new_n209), .c(new_n215), .d(new_n221), .out0(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n257));
  aoi012aa1n12x5               g162(.a(new_n245), .b(new_n235), .c(new_n246), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n258), .o1(new_n259));
  aoi012aa1n02x5               g164(.a(new_n259), .b(new_n234), .c(new_n254), .o1(new_n260));
  inv040aa1n03x5               g165(.a(new_n260), .o1(new_n261));
  xorc02aa1n12x5               g166(.a(\a[23] ), .b(\b[22] ), .out0(new_n262));
  aoai13aa1n06x5               g167(.a(new_n262), .b(new_n261), .c(new_n195), .d(new_n256), .o1(new_n263));
  aoi112aa1n02x5               g168(.a(new_n262), .b(new_n259), .c(new_n234), .d(new_n254), .o1(new_n264));
  aobi12aa1n02x7               g169(.a(new_n263), .b(new_n264), .c(new_n257), .out0(\s[23] ));
  xorc02aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .out0(new_n266));
  nor042aa1n06x5               g171(.a(\b[22] ), .b(\a[23] ), .o1(new_n267));
  norp02aa1n02x5               g172(.a(new_n266), .b(new_n267), .o1(new_n268));
  inv000aa1d42x5               g173(.a(new_n267), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n262), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n269), .b(new_n270), .c(new_n257), .d(new_n260), .o1(new_n271));
  aoi022aa1n02x7               g176(.a(new_n271), .b(new_n266), .c(new_n263), .d(new_n268), .o1(\s[24] ));
  nano32aa1n03x7               g177(.a(new_n270), .b(new_n266), .c(new_n237), .d(new_n247), .out0(new_n273));
  and002aa1n02x5               g178(.a(new_n273), .b(new_n229), .o(new_n274));
  aoai13aa1n02x5               g179(.a(new_n274), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n275));
  aoai13aa1n06x5               g180(.a(new_n254), .b(new_n242), .c(new_n241), .d(new_n239), .o1(new_n276));
  and002aa1n03x5               g181(.a(new_n266), .b(new_n262), .o(new_n277));
  inv000aa1n06x5               g182(.a(new_n277), .o1(new_n278));
  oao003aa1n02x5               g183(.a(\a[24] ), .b(\b[23] ), .c(new_n269), .carry(new_n279));
  aoai13aa1n12x5               g184(.a(new_n279), .b(new_n278), .c(new_n276), .d(new_n258), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[25] ), .b(\b[24] ), .out0(new_n281));
  aoai13aa1n06x5               g186(.a(new_n281), .b(new_n280), .c(new_n195), .d(new_n274), .o1(new_n282));
  aoai13aa1n06x5               g187(.a(new_n277), .b(new_n259), .c(new_n234), .d(new_n254), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n281), .o1(new_n284));
  and003aa1n02x5               g189(.a(new_n283), .b(new_n284), .c(new_n279), .o(new_n285));
  aobi12aa1n03x7               g190(.a(new_n282), .b(new_n285), .c(new_n275), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g191(.a(\a[26] ), .b(\b[25] ), .out0(new_n287));
  nor042aa1n03x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  norp02aa1n02x5               g193(.a(new_n287), .b(new_n288), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n280), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n288), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n284), .c(new_n275), .d(new_n290), .o1(new_n292));
  aoi022aa1n03x5               g197(.a(new_n292), .b(new_n287), .c(new_n282), .d(new_n289), .o1(\s[26] ));
  and002aa1n12x5               g198(.a(new_n287), .b(new_n281), .o(new_n294));
  and003aa1n18x5               g199(.a(new_n273), .b(new_n229), .c(new_n294), .o(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n203), .c(new_n128), .d(new_n184), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n294), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[26] ), .b(\b[25] ), .c(new_n291), .carry(new_n298));
  aoai13aa1n04x5               g203(.a(new_n298), .b(new_n297), .c(new_n283), .d(new_n279), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  aoai13aa1n06x5               g205(.a(new_n300), .b(new_n299), .c(new_n195), .d(new_n295), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n298), .o1(new_n302));
  aoi112aa1n02x5               g207(.a(new_n300), .b(new_n302), .c(new_n280), .d(new_n294), .o1(new_n303));
  aobi12aa1n02x7               g208(.a(new_n301), .b(new_n303), .c(new_n296), .out0(\s[27] ));
  tech160nm_fixorc02aa1n04x5   g209(.a(\a[28] ), .b(\b[27] ), .out0(new_n305));
  norp02aa1n02x5               g210(.a(\b[26] ), .b(\a[27] ), .o1(new_n306));
  norp02aa1n02x5               g211(.a(new_n305), .b(new_n306), .o1(new_n307));
  tech160nm_fiaoi012aa1n05x5   g212(.a(new_n302), .b(new_n280), .c(new_n294), .o1(new_n308));
  inv000aa1n03x5               g213(.a(new_n306), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n300), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n309), .b(new_n310), .c(new_n308), .d(new_n296), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n311), .b(new_n305), .c(new_n301), .d(new_n307), .o1(\s[28] ));
  and002aa1n02x5               g217(.a(new_n305), .b(new_n300), .o(new_n313));
  aoai13aa1n03x5               g218(.a(new_n313), .b(new_n299), .c(new_n195), .d(new_n295), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[29] ), .b(\b[28] ), .out0(new_n315));
  oao003aa1n02x5               g220(.a(\a[28] ), .b(\b[27] ), .c(new_n309), .carry(new_n316));
  norb02aa1n02x5               g221(.a(new_n316), .b(new_n315), .out0(new_n317));
  inv000aa1d42x5               g222(.a(new_n313), .o1(new_n318));
  aoai13aa1n02x7               g223(.a(new_n316), .b(new_n318), .c(new_n308), .d(new_n296), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n319), .b(new_n315), .c(new_n314), .d(new_n317), .o1(\s[29] ));
  xorb03aa1n02x5               g225(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g226(.a(new_n310), .b(new_n305), .c(new_n315), .out0(new_n322));
  aoai13aa1n06x5               g227(.a(new_n322), .b(new_n299), .c(new_n195), .d(new_n295), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .out0(new_n324));
  inv000aa1d42x5               g229(.a(\a[29] ), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[28] ), .o1(new_n326));
  oaib12aa1n02x5               g231(.a(new_n316), .b(\b[28] ), .c(new_n325), .out0(new_n327));
  oaoi13aa1n02x5               g232(.a(new_n324), .b(new_n327), .c(new_n325), .d(new_n326), .o1(new_n328));
  inv000aa1n02x5               g233(.a(new_n322), .o1(new_n329));
  oaib12aa1n02x5               g234(.a(new_n327), .b(new_n326), .c(\a[29] ), .out0(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n329), .c(new_n308), .d(new_n296), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n331), .b(new_n324), .c(new_n323), .d(new_n328), .o1(\s[30] ));
  nano32aa1n02x4               g237(.a(new_n310), .b(new_n324), .c(new_n305), .d(new_n315), .out0(new_n333));
  aoai13aa1n03x5               g238(.a(new_n333), .b(new_n299), .c(new_n195), .d(new_n295), .o1(new_n334));
  aoi022aa1n02x5               g239(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n335));
  norb02aa1n02x5               g240(.a(\b[30] ), .b(\a[31] ), .out0(new_n336));
  obai22aa1n02x7               g241(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n337));
  aoi112aa1n02x5               g242(.a(new_n337), .b(new_n336), .c(new_n327), .d(new_n335), .o1(new_n338));
  inv000aa1n02x5               g243(.a(new_n333), .o1(new_n339));
  norp02aa1n02x5               g244(.a(\b[29] ), .b(\a[30] ), .o1(new_n340));
  aoi012aa1n02x5               g245(.a(new_n340), .b(new_n327), .c(new_n335), .o1(new_n341));
  aoai13aa1n02x7               g246(.a(new_n341), .b(new_n339), .c(new_n308), .d(new_n296), .o1(new_n342));
  xorc02aa1n02x5               g247(.a(\a[31] ), .b(\b[30] ), .out0(new_n343));
  aoi022aa1n02x7               g248(.a(new_n342), .b(new_n343), .c(new_n338), .d(new_n334), .o1(\s[31] ));
  inv000aa1d42x5               g249(.a(\b[1] ), .o1(new_n345));
  inv000aa1d42x5               g250(.a(\a[2] ), .o1(new_n346));
  aoi022aa1n02x5               g251(.a(new_n345), .b(new_n346), .c(\a[1] ), .d(\b[0] ), .o1(new_n347));
  oaib12aa1n02x5               g252(.a(new_n347), .b(new_n345), .c(\a[2] ), .out0(new_n348));
  aboi22aa1n03x5               g253(.a(new_n105), .b(new_n106), .c(new_n346), .d(new_n345), .out0(new_n349));
  aoi022aa1n02x5               g254(.a(new_n348), .b(new_n349), .c(new_n101), .d(new_n107), .o1(\s[3] ));
  aoai13aa1n02x5               g255(.a(new_n104), .b(new_n105), .c(new_n101), .d(new_n106), .o1(new_n351));
  aoi112aa1n02x5               g256(.a(new_n105), .b(new_n104), .c(new_n101), .d(new_n106), .o1(new_n352));
  norb02aa1n02x5               g257(.a(new_n351), .b(new_n352), .out0(\s[4] ));
  norb02aa1n02x5               g258(.a(new_n113), .b(new_n112), .out0(new_n354));
  xnbna2aa1n03x5               g259(.a(new_n354), .b(new_n108), .c(new_n109), .out0(\s[5] ));
  inv000aa1d42x5               g260(.a(new_n112), .o1(new_n356));
  nanp02aa1n02x5               g261(.a(new_n108), .b(new_n109), .o1(new_n357));
  nanp02aa1n02x5               g262(.a(new_n357), .b(new_n354), .o1(new_n358));
  xnbna2aa1n03x5               g263(.a(new_n117), .b(new_n358), .c(new_n356), .out0(\s[6] ));
  norb02aa1n02x5               g264(.a(new_n111), .b(new_n110), .out0(new_n360));
  inv000aa1d42x5               g265(.a(new_n116), .o1(new_n361));
  aoai13aa1n02x5               g266(.a(new_n117), .b(new_n112), .c(new_n357), .d(new_n113), .o1(new_n362));
  xnbna2aa1n03x5               g267(.a(new_n360), .b(new_n362), .c(new_n361), .out0(\s[7] ));
  aob012aa1n02x5               g268(.a(new_n360), .b(new_n362), .c(new_n361), .out0(new_n364));
  oai012aa1n02x5               g269(.a(new_n364), .b(\b[6] ), .c(\a[7] ), .o1(new_n365));
  aoib12aa1n02x5               g270(.a(new_n110), .b(new_n119), .c(new_n118), .out0(new_n366));
  aoi022aa1n02x5               g271(.a(new_n365), .b(new_n120), .c(new_n364), .d(new_n366), .o1(\s[8] ));
  aoi012aa1n02x5               g272(.a(new_n121), .b(new_n108), .c(new_n109), .o1(new_n368));
  aoi112aa1n02x5               g273(.a(new_n126), .b(new_n129), .c(new_n124), .d(new_n122), .o1(new_n369));
  aboi22aa1n03x5               g274(.a(new_n368), .b(new_n369), .c(new_n128), .d(new_n129), .out0(\s[9] ));
endmodule


