// Benchmark "adder" written by ABC on Thu Jul 18 11:53:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n342, new_n343, new_n344, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n352, new_n353, new_n354,
    new_n356, new_n358, new_n359, new_n360;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  oai022aa1n02x5               g002(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n98));
  xorc02aa1n03x5               g003(.a(\a[3] ), .b(\b[2] ), .out0(new_n99));
  and002aa1n12x5               g004(.a(\b[1] ), .b(\a[2] ), .o(new_n100));
  nand22aa1n06x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor022aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oab012aa1n09x5               g007(.a(new_n100), .b(new_n102), .c(new_n101), .out0(new_n103));
  aoi012aa1n12x5               g008(.a(new_n98), .b(new_n103), .c(new_n99), .o1(new_n104));
  nand42aa1n10x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  aob012aa1d18x5               g010(.a(new_n105), .b(\b[7] ), .c(\a[8] ), .out0(new_n106));
  nor002aa1d32x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nor042aa1d18x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand02aa1n06x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  norb03aa1d15x5               g014(.a(new_n109), .b(new_n107), .c(new_n108), .out0(new_n110));
  inv000aa1d42x5               g015(.a(\a[8] ), .o1(new_n111));
  inv000aa1d42x5               g016(.a(\b[7] ), .o1(new_n112));
  aoi022aa1n12x5               g017(.a(new_n112), .b(new_n111), .c(\a[5] ), .d(\b[4] ), .o1(new_n113));
  nand02aa1d16x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  oai012aa1n12x5               g019(.a(new_n114), .b(\b[4] ), .c(\a[5] ), .o1(new_n115));
  nona23aa1d24x5               g020(.a(new_n110), .b(new_n113), .c(new_n106), .d(new_n115), .out0(new_n116));
  inv000aa1d42x5               g021(.a(new_n108), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\a[5] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[4] ), .o1(new_n119));
  aoai13aa1n12x5               g024(.a(new_n114), .b(new_n107), .c(new_n118), .d(new_n119), .o1(new_n120));
  nand02aa1n02x5               g025(.a(new_n120), .b(new_n117), .o1(new_n121));
  aoi022aa1n12x5               g026(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n122));
  aoi022aa1n12x5               g027(.a(new_n121), .b(new_n122), .c(new_n112), .d(new_n111), .o1(new_n123));
  oai012aa1d24x5               g028(.a(new_n123), .b(new_n104), .c(new_n116), .o1(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  nor042aa1n03x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand42aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1n06x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n97), .c(new_n124), .d(new_n125), .o1(new_n129));
  aoi112aa1n02x5               g034(.a(new_n128), .b(new_n97), .c(new_n124), .d(new_n125), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(\s[10] ));
  oai012aa1n02x5               g036(.a(new_n127), .b(new_n126), .c(new_n97), .o1(new_n132));
  nor042aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n129), .c(new_n132), .out0(\s[11] ));
  nand02aa1n03x5               g041(.a(new_n129), .b(new_n132), .o1(new_n137));
  nor042aa1n03x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1n06x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n133), .c(new_n137), .d(new_n134), .o1(new_n142));
  aoi112aa1n02x5               g047(.a(new_n133), .b(new_n141), .c(new_n137), .d(new_n134), .o1(new_n143));
  nanb02aa1n03x5               g048(.a(new_n143), .b(new_n142), .out0(\s[12] ));
  xnrc02aa1n02x5               g049(.a(\b[2] ), .b(\a[3] ), .out0(new_n145));
  oabi12aa1n02x5               g050(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n146));
  oabi12aa1n02x5               g051(.a(new_n98), .b(new_n146), .c(new_n145), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n116), .o1(new_n148));
  nanp02aa1n02x5               g053(.a(new_n112), .b(new_n111), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n122), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n149), .b(new_n150), .c(new_n120), .d(new_n117), .o1(new_n151));
  nano23aa1n09x5               g056(.a(new_n133), .b(new_n138), .c(new_n139), .d(new_n134), .out0(new_n152));
  nand23aa1d12x5               g057(.a(new_n152), .b(new_n125), .c(new_n128), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n02x5               g059(.a(new_n154), .b(new_n151), .c(new_n148), .d(new_n147), .o1(new_n155));
  nano22aa1n03x7               g060(.a(new_n138), .b(new_n134), .c(new_n139), .out0(new_n156));
  oai012aa1n02x5               g061(.a(new_n127), .b(\b[10] ), .c(\a[11] ), .o1(new_n157));
  oab012aa1n04x5               g062(.a(new_n157), .b(new_n97), .c(new_n126), .out0(new_n158));
  nanp02aa1n02x5               g063(.a(new_n158), .b(new_n156), .o1(new_n159));
  aoi012aa1n09x5               g064(.a(new_n138), .b(new_n133), .c(new_n139), .o1(new_n160));
  nand02aa1d04x5               g065(.a(new_n159), .b(new_n160), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nor042aa1n09x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nand42aa1n03x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  xobna2aa1n03x5               g070(.a(new_n165), .b(new_n155), .c(new_n162), .out0(\s[13] ));
  inv000aa1d42x5               g071(.a(new_n163), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n167), .b(new_n165), .c(new_n155), .d(new_n162), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n02x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nanp02aa1n04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nano23aa1d12x5               g076(.a(new_n163), .b(new_n170), .c(new_n171), .d(new_n164), .out0(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n161), .c(new_n124), .d(new_n154), .o1(new_n173));
  aoi012aa1n09x5               g078(.a(new_n170), .b(new_n163), .c(new_n171), .o1(new_n174));
  xorc02aa1n12x5               g079(.a(\a[15] ), .b(\b[14] ), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n173), .c(new_n174), .out0(\s[15] ));
  nanp02aa1n06x5               g081(.a(new_n173), .b(new_n174), .o1(new_n177));
  nor002aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  xorc02aa1n12x5               g083(.a(\a[16] ), .b(\b[15] ), .out0(new_n179));
  inv000aa1d42x5               g084(.a(new_n179), .o1(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n178), .c(new_n177), .d(new_n175), .o1(new_n181));
  aoi112aa1n03x4               g086(.a(new_n178), .b(new_n180), .c(new_n177), .d(new_n175), .o1(new_n182));
  nanb02aa1n03x5               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  nano32aa1d12x5               g088(.a(new_n153), .b(new_n179), .c(new_n172), .d(new_n175), .out0(new_n184));
  nand22aa1n06x5               g089(.a(new_n124), .b(new_n184), .o1(new_n185));
  and002aa1n06x5               g090(.a(new_n179), .b(new_n175), .o(new_n186));
  inv030aa1n03x5               g091(.a(new_n160), .o1(new_n187));
  aoai13aa1n06x5               g092(.a(new_n172), .b(new_n187), .c(new_n158), .d(new_n156), .o1(new_n188));
  nand42aa1n02x5               g093(.a(new_n188), .b(new_n174), .o1(new_n189));
  nanp02aa1n06x5               g094(.a(new_n189), .b(new_n186), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\a[16] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[15] ), .o1(new_n192));
  oao003aa1n02x5               g097(.a(new_n191), .b(new_n192), .c(new_n178), .carry(new_n193));
  inv000aa1n02x5               g098(.a(new_n193), .o1(new_n194));
  nand23aa1n09x5               g099(.a(new_n185), .b(new_n190), .c(new_n194), .o1(new_n195));
  nor042aa1d18x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nand02aa1n06x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  aoi112aa1n02x5               g103(.a(new_n193), .b(new_n198), .c(new_n189), .d(new_n186), .o1(new_n199));
  aoi022aa1n02x5               g104(.a(new_n195), .b(new_n198), .c(new_n199), .d(new_n185), .o1(\s[17] ));
  inv000aa1n04x5               g105(.a(new_n186), .o1(new_n201));
  tech160nm_fiaoi012aa1n04x5   g106(.a(new_n201), .b(new_n188), .c(new_n174), .o1(new_n202));
  aoi112aa1n09x5               g107(.a(new_n202), .b(new_n193), .c(new_n124), .d(new_n184), .o1(new_n203));
  oaoi03aa1n03x5               g108(.a(\a[17] ), .b(\b[16] ), .c(new_n203), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor002aa1n20x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand42aa1n16x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nano23aa1n06x5               g112(.a(new_n196), .b(new_n206), .c(new_n207), .d(new_n197), .out0(new_n208));
  inv000aa1n04x5               g113(.a(new_n208), .o1(new_n209));
  oa0012aa1n02x5               g114(.a(new_n207), .b(new_n206), .c(new_n196), .o(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  oaih12aa1n04x5               g116(.a(new_n211), .b(new_n203), .c(new_n209), .o1(new_n212));
  nor042aa1d18x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand02aa1d10x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n06x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  aoi112aa1n03x4               g120(.a(new_n215), .b(new_n210), .c(new_n195), .d(new_n208), .o1(new_n216));
  aoi012aa1n02x5               g121(.a(new_n216), .b(new_n212), .c(new_n215), .o1(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand02aa1d28x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nanb02aa1n02x5               g125(.a(new_n219), .b(new_n220), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n213), .c(new_n212), .d(new_n214), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n215), .b(new_n210), .c(new_n195), .d(new_n208), .o1(new_n223));
  nona22aa1n06x5               g128(.a(new_n223), .b(new_n221), .c(new_n213), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n222), .b(new_n224), .o1(\s[20] ));
  inv000aa1d42x5               g130(.a(new_n219), .o1(new_n226));
  nano32aa1n03x7               g131(.a(new_n209), .b(new_n220), .c(new_n215), .d(new_n226), .out0(new_n227));
  inv000aa1n03x5               g132(.a(new_n227), .o1(new_n228));
  nanb03aa1n12x5               g133(.a(new_n219), .b(new_n220), .c(new_n214), .out0(new_n229));
  orn002aa1n03x5               g134(.a(\a[19] ), .b(\b[18] ), .o(new_n230));
  oai112aa1n06x5               g135(.a(new_n230), .b(new_n207), .c(new_n206), .d(new_n196), .o1(new_n231));
  aoi012aa1d24x5               g136(.a(new_n219), .b(new_n213), .c(new_n220), .o1(new_n232));
  oai012aa1d24x5               g137(.a(new_n232), .b(new_n231), .c(new_n229), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  oai012aa1n06x5               g139(.a(new_n234), .b(new_n203), .c(new_n228), .o1(new_n235));
  nor002aa1d32x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nand42aa1d28x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  aoi112aa1n02x5               g143(.a(new_n238), .b(new_n233), .c(new_n195), .d(new_n227), .o1(new_n239));
  aoi012aa1n02x5               g144(.a(new_n239), .b(new_n235), .c(new_n238), .o1(\s[21] ));
  nor002aa1n20x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  nand42aa1n20x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  nanb02aa1n02x5               g147(.a(new_n241), .b(new_n242), .out0(new_n243));
  aoai13aa1n03x5               g148(.a(new_n243), .b(new_n236), .c(new_n235), .d(new_n238), .o1(new_n244));
  aoai13aa1n03x5               g149(.a(new_n238), .b(new_n233), .c(new_n195), .d(new_n227), .o1(new_n245));
  nona22aa1n03x5               g150(.a(new_n245), .b(new_n243), .c(new_n236), .out0(new_n246));
  nanp02aa1n03x5               g151(.a(new_n244), .b(new_n246), .o1(\s[22] ));
  aoai13aa1n03x5               g152(.a(new_n194), .b(new_n201), .c(new_n188), .d(new_n174), .o1(new_n248));
  nano23aa1d15x5               g153(.a(new_n236), .b(new_n241), .c(new_n242), .d(new_n237), .out0(new_n249));
  nano32aa1n03x7               g154(.a(new_n221), .b(new_n249), .c(new_n208), .d(new_n215), .out0(new_n250));
  aoai13aa1n02x5               g155(.a(new_n250), .b(new_n248), .c(new_n124), .d(new_n184), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n250), .o1(new_n252));
  oa0012aa1n06x5               g157(.a(new_n242), .b(new_n241), .c(new_n236), .o(new_n253));
  aoi012aa1d24x5               g158(.a(new_n253), .b(new_n233), .c(new_n249), .o1(new_n254));
  oai012aa1n06x5               g159(.a(new_n254), .b(new_n203), .c(new_n252), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  aoi112aa1n02x5               g161(.a(new_n256), .b(new_n253), .c(new_n233), .d(new_n249), .o1(new_n257));
  aoi022aa1n02x5               g162(.a(new_n255), .b(new_n256), .c(new_n251), .d(new_n257), .o1(\s[23] ));
  norp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[23] ), .b(\a[24] ), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n259), .c(new_n255), .d(new_n256), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n254), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n256), .b(new_n262), .c(new_n195), .d(new_n250), .o1(new_n263));
  nona22aa1n03x5               g168(.a(new_n263), .b(new_n260), .c(new_n259), .out0(new_n264));
  nanp02aa1n03x5               g169(.a(new_n261), .b(new_n264), .o1(\s[24] ));
  norb02aa1n06x4               g170(.a(new_n256), .b(new_n260), .out0(new_n266));
  nano22aa1n03x7               g171(.a(new_n228), .b(new_n249), .c(new_n266), .out0(new_n267));
  aoai13aa1n02x5               g172(.a(new_n267), .b(new_n248), .c(new_n124), .d(new_n184), .o1(new_n268));
  inv000aa1n02x5               g173(.a(new_n267), .o1(new_n269));
  nano22aa1n02x5               g174(.a(new_n219), .b(new_n214), .c(new_n220), .out0(new_n270));
  tech160nm_fioai012aa1n03p5x5 g175(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .o1(new_n271));
  oab012aa1n02x5               g176(.a(new_n271), .b(new_n196), .c(new_n206), .out0(new_n272));
  inv020aa1n03x5               g177(.a(new_n232), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n249), .b(new_n273), .c(new_n272), .d(new_n270), .o1(new_n274));
  inv040aa1n03x5               g179(.a(new_n253), .o1(new_n275));
  inv040aa1n02x5               g180(.a(new_n266), .o1(new_n276));
  oai022aa1n02x5               g181(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n277));
  aob012aa1n02x5               g182(.a(new_n277), .b(\b[23] ), .c(\a[24] ), .out0(new_n278));
  aoai13aa1n12x5               g183(.a(new_n278), .b(new_n276), .c(new_n274), .d(new_n275), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  oai012aa1n04x7               g185(.a(new_n280), .b(new_n203), .c(new_n269), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n266), .b(new_n253), .c(new_n233), .d(new_n249), .o1(new_n283));
  nano22aa1n02x4               g188(.a(new_n282), .b(new_n283), .c(new_n278), .out0(new_n284));
  aoi022aa1n02x5               g189(.a(new_n281), .b(new_n282), .c(new_n268), .d(new_n284), .o1(\s[25] ));
  nor002aa1n02x5               g190(.a(\b[24] ), .b(\a[25] ), .o1(new_n286));
  xnrc02aa1n12x5               g191(.a(\b[25] ), .b(\a[26] ), .out0(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n286), .c(new_n281), .d(new_n282), .o1(new_n288));
  aoai13aa1n02x7               g193(.a(new_n282), .b(new_n279), .c(new_n195), .d(new_n267), .o1(new_n289));
  nona22aa1n03x5               g194(.a(new_n289), .b(new_n287), .c(new_n286), .out0(new_n290));
  nanp02aa1n03x5               g195(.a(new_n288), .b(new_n290), .o1(\s[26] ));
  norb02aa1n15x5               g196(.a(new_n282), .b(new_n287), .out0(new_n292));
  nano32aa1n03x7               g197(.a(new_n228), .b(new_n292), .c(new_n249), .d(new_n266), .out0(new_n293));
  aoai13aa1n06x5               g198(.a(new_n293), .b(new_n248), .c(new_n124), .d(new_n184), .o1(new_n294));
  inv000aa1n02x5               g199(.a(new_n293), .o1(new_n295));
  inv000aa1d42x5               g200(.a(\a[26] ), .o1(new_n296));
  inv000aa1d42x5               g201(.a(\b[25] ), .o1(new_n297));
  oao003aa1n02x5               g202(.a(new_n296), .b(new_n297), .c(new_n286), .carry(new_n298));
  aoi012aa1n09x5               g203(.a(new_n298), .b(new_n279), .c(new_n292), .o1(new_n299));
  oai012aa1n06x5               g204(.a(new_n299), .b(new_n203), .c(new_n295), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  aoi112aa1n02x5               g206(.a(new_n301), .b(new_n298), .c(new_n279), .d(new_n292), .o1(new_n302));
  aoi022aa1n02x5               g207(.a(new_n300), .b(new_n301), .c(new_n294), .d(new_n302), .o1(\s[27] ));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  norp02aa1n04x5               g209(.a(\b[27] ), .b(\a[28] ), .o1(new_n305));
  nand42aa1n03x5               g210(.a(\b[27] ), .b(\a[28] ), .o1(new_n306));
  nanb02aa1n06x5               g211(.a(new_n305), .b(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n304), .c(new_n300), .d(new_n301), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n292), .o1(new_n309));
  inv000aa1n02x5               g214(.a(new_n298), .o1(new_n310));
  aoai13aa1n04x5               g215(.a(new_n310), .b(new_n309), .c(new_n283), .d(new_n278), .o1(new_n311));
  aoai13aa1n02x5               g216(.a(new_n301), .b(new_n311), .c(new_n195), .d(new_n293), .o1(new_n312));
  nona22aa1n02x4               g217(.a(new_n312), .b(new_n307), .c(new_n304), .out0(new_n313));
  nanp02aa1n03x5               g218(.a(new_n308), .b(new_n313), .o1(\s[28] ));
  norb02aa1n03x5               g219(.a(new_n301), .b(new_n307), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n195), .d(new_n293), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n315), .o1(new_n317));
  aoi012aa1n02x5               g222(.a(new_n305), .b(new_n304), .c(new_n306), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n317), .c(new_n294), .d(new_n299), .o1(new_n319));
  xorc02aa1n12x5               g224(.a(\a[29] ), .b(\b[28] ), .out0(new_n320));
  norb02aa1n02x5               g225(.a(new_n318), .b(new_n320), .out0(new_n321));
  aoi022aa1n03x5               g226(.a(new_n319), .b(new_n320), .c(new_n316), .d(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g228(.a(new_n307), .b(new_n301), .c(new_n320), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n311), .c(new_n195), .d(new_n293), .o1(new_n325));
  inv000aa1d42x5               g230(.a(new_n324), .o1(new_n326));
  oao003aa1n02x5               g231(.a(\a[29] ), .b(\b[28] ), .c(new_n318), .carry(new_n327));
  aoai13aa1n02x7               g232(.a(new_n327), .b(new_n326), .c(new_n294), .d(new_n299), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[30] ), .b(\b[29] ), .out0(new_n329));
  norb02aa1n02x5               g234(.a(new_n327), .b(new_n329), .out0(new_n330));
  aoi022aa1n03x5               g235(.a(new_n328), .b(new_n329), .c(new_n325), .d(new_n330), .o1(\s[30] ));
  nand03aa1n02x5               g236(.a(new_n315), .b(new_n320), .c(new_n329), .o1(new_n332));
  nanb02aa1n03x5               g237(.a(new_n332), .b(new_n300), .out0(new_n333));
  oao003aa1n02x5               g238(.a(\a[30] ), .b(\b[29] ), .c(new_n327), .carry(new_n334));
  aoai13aa1n02x7               g239(.a(new_n334), .b(new_n332), .c(new_n294), .d(new_n299), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  and002aa1n02x5               g241(.a(\b[29] ), .b(\a[30] ), .o(new_n337));
  oabi12aa1n02x5               g242(.a(new_n336), .b(\a[30] ), .c(\b[29] ), .out0(new_n338));
  oab012aa1n02x4               g243(.a(new_n338), .b(new_n327), .c(new_n337), .out0(new_n339));
  aoi022aa1n03x5               g244(.a(new_n335), .b(new_n336), .c(new_n333), .d(new_n339), .o1(\s[31] ));
  xorb03aa1n02x5               g245(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g246(.a(new_n103), .b(new_n99), .o1(new_n342));
  xorc02aa1n02x5               g247(.a(\a[4] ), .b(\b[3] ), .out0(new_n343));
  oab012aa1n02x4               g248(.a(new_n343), .b(\a[3] ), .c(\b[2] ), .out0(new_n344));
  aoi022aa1n02x5               g249(.a(new_n147), .b(new_n343), .c(new_n344), .d(new_n342), .o1(\s[4] ));
  nanp02aa1n02x5               g250(.a(\b[4] ), .b(\a[5] ), .o1(new_n346));
  nanp02aa1n02x5               g251(.a(new_n119), .b(new_n118), .o1(new_n347));
  aoi022aa1n02x5               g252(.a(new_n147), .b(new_n105), .c(new_n347), .d(new_n346), .o1(new_n348));
  aoi022aa1n02x5               g253(.a(new_n119), .b(new_n118), .c(\a[4] ), .d(\b[3] ), .o1(new_n349));
  nano22aa1n03x7               g254(.a(new_n104), .b(new_n346), .c(new_n349), .out0(new_n350));
  norp02aa1n02x5               g255(.a(new_n348), .b(new_n350), .o1(\s[5] ));
  norb02aa1n02x5               g256(.a(new_n114), .b(new_n107), .out0(new_n352));
  aoai13aa1n06x5               g257(.a(new_n352), .b(new_n350), .c(new_n118), .d(new_n119), .o1(new_n353));
  aoi112aa1n02x5               g258(.a(new_n350), .b(new_n352), .c(new_n118), .d(new_n119), .o1(new_n354));
  norb02aa1n02x5               g259(.a(new_n353), .b(new_n354), .out0(\s[6] ));
  norb02aa1n02x5               g260(.a(new_n109), .b(new_n108), .out0(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n356), .b(new_n353), .c(new_n120), .out0(\s[7] ));
  nanp02aa1n02x5               g262(.a(new_n353), .b(new_n120), .o1(new_n358));
  nanp02aa1n02x5               g263(.a(new_n358), .b(new_n356), .o1(new_n359));
  xorc02aa1n02x5               g264(.a(\a[8] ), .b(\b[7] ), .out0(new_n360));
  xnbna2aa1n03x5               g265(.a(new_n360), .b(new_n359), .c(new_n117), .out0(\s[8] ));
  xorb03aa1n02x5               g266(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


