// Benchmark "adder" written by ABC on Thu Jul 18 05:33:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n322, new_n325, new_n327,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n09x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n16x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n06x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nand42aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor042aa1d18x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  orn002aa1n03x5               g006(.a(\a[2] ), .b(\b[1] ), .o(new_n102));
  nand02aa1d08x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  nand02aa1d16x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  aob012aa1n06x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .out0(new_n105));
  nor042aa1n04x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nand02aa1d08x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  norb02aa1n03x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nor042aa1n06x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nand02aa1d04x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  norb02aa1n03x5               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  nand23aa1n06x5               g016(.a(new_n105), .b(new_n108), .c(new_n111), .o1(new_n112));
  tech160nm_fiaoi012aa1n04x5   g017(.a(new_n106), .b(new_n109), .c(new_n107), .o1(new_n113));
  nor042aa1n03x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand42aa1d28x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nor002aa1n06x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n16x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nano23aa1n09x5               g022(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n118));
  nor022aa1n16x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nand02aa1n04x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nor022aa1n16x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nand02aa1n06x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  nano23aa1n03x7               g027(.a(new_n119), .b(new_n121), .c(new_n122), .d(new_n120), .out0(new_n123));
  nand02aa1n02x5               g028(.a(new_n123), .b(new_n118), .o1(new_n124));
  and002aa1n12x5               g029(.a(\b[5] ), .b(\a[6] ), .o(new_n125));
  oab012aa1n09x5               g030(.a(new_n125), .b(new_n119), .c(new_n121), .out0(new_n126));
  oai022aa1n09x5               g031(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n127));
  aoi022aa1n12x5               g032(.a(new_n118), .b(new_n126), .c(new_n115), .d(new_n127), .o1(new_n128));
  aoai13aa1n12x5               g033(.a(new_n128), .b(new_n124), .c(new_n112), .d(new_n113), .o1(new_n129));
  nor042aa1n03x5               g034(.a(new_n129), .b(new_n101), .o1(new_n130));
  nano22aa1n03x7               g035(.a(new_n130), .b(new_n99), .c(new_n100), .out0(new_n131));
  oaoi13aa1n02x5               g036(.a(new_n99), .b(new_n100), .c(new_n129), .d(new_n101), .o1(new_n132));
  norp02aa1n02x5               g037(.a(new_n132), .b(new_n131), .o1(\s[10] ));
  oai112aa1n04x5               g038(.a(new_n100), .b(new_n99), .c(new_n129), .d(new_n101), .o1(new_n134));
  aoi012aa1d18x5               g039(.a(new_n97), .b(new_n101), .c(new_n98), .o1(new_n135));
  nor002aa1d32x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand42aa1n16x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanb02aa1d36x5               g042(.a(new_n136), .b(new_n137), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n134), .c(new_n135), .out0(\s[11] ));
  inv000aa1d42x5               g045(.a(new_n136), .o1(new_n141));
  inv000aa1d42x5               g046(.a(new_n135), .o1(new_n142));
  tech160nm_fioai012aa1n03p5x5 g047(.a(new_n139), .b(new_n131), .c(new_n142), .o1(new_n143));
  nor002aa1n03x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand02aa1n06x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nanb02aa1n12x5               g050(.a(new_n144), .b(new_n145), .out0(new_n146));
  aoi012aa1n02x5               g051(.a(new_n146), .b(new_n143), .c(new_n141), .o1(new_n147));
  aoi012aa1n02x5               g052(.a(new_n138), .b(new_n134), .c(new_n135), .o1(new_n148));
  nano22aa1n03x5               g053(.a(new_n148), .b(new_n141), .c(new_n146), .out0(new_n149));
  norp02aa1n02x5               g054(.a(new_n147), .b(new_n149), .o1(\s[12] ));
  norb02aa1n06x5               g055(.a(new_n100), .b(new_n101), .out0(new_n151));
  nona23aa1d24x5               g056(.a(new_n99), .b(new_n151), .c(new_n146), .d(new_n138), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n06x5               g058(.a(new_n137), .b(new_n97), .c(new_n101), .d(new_n98), .o1(new_n154));
  nor002aa1n02x5               g059(.a(new_n144), .b(new_n136), .o1(new_n155));
  aob012aa1d15x5               g060(.a(new_n145), .b(new_n154), .c(new_n155), .out0(new_n156));
  aob012aa1n02x5               g061(.a(new_n156), .b(new_n129), .c(new_n153), .out0(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n08x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norp02aa1n12x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand42aa1n08x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  aoi112aa1n02x5               g068(.a(new_n159), .b(new_n163), .c(new_n157), .d(new_n160), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n156), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n159), .b(new_n161), .c(new_n162), .d(new_n160), .out0(new_n166));
  aoai13aa1n06x5               g071(.a(new_n166), .b(new_n165), .c(new_n129), .d(new_n153), .o1(new_n167));
  oa0012aa1n12x5               g072(.a(new_n162), .b(new_n161), .c(new_n159), .o(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  aoi012aa1n02x5               g074(.a(new_n161), .b(new_n167), .c(new_n169), .o1(new_n170));
  norp02aa1n02x5               g075(.a(new_n164), .b(new_n170), .o1(\s[14] ));
  xnrc02aa1n12x5               g076(.a(\b[14] ), .b(\a[15] ), .out0(new_n172));
  xobna2aa1n03x5               g077(.a(new_n172), .b(new_n167), .c(new_n169), .out0(\s[15] ));
  norp02aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  aoai13aa1n04x5               g080(.a(new_n175), .b(new_n172), .c(new_n167), .d(new_n169), .o1(new_n176));
  xnrc02aa1n03x5               g081(.a(\b[15] ), .b(\a[16] ), .out0(new_n177));
  nanp02aa1n02x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  oai022aa1n02x5               g083(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n02x5               g085(.a(new_n180), .b(new_n172), .c(new_n167), .d(new_n169), .o1(new_n181));
  aob012aa1n03x5               g086(.a(new_n181), .b(new_n176), .c(new_n177), .out0(\s[16] ));
  nona22aa1n09x5               g087(.a(new_n166), .b(new_n172), .c(new_n177), .out0(new_n183));
  nor042aa1d18x5               g088(.a(new_n152), .b(new_n183), .o1(new_n184));
  tech160nm_finand02aa1n05x5   g089(.a(new_n129), .b(new_n184), .o1(new_n185));
  nor022aa1n04x5               g090(.a(new_n177), .b(new_n172), .o1(new_n186));
  aoi022aa1n06x5               g091(.a(new_n186), .b(new_n168), .c(new_n178), .d(new_n179), .o1(new_n187));
  oaih12aa1n12x5               g092(.a(new_n187), .b(new_n156), .c(new_n183), .o1(new_n188));
  nanb02aa1n09x5               g093(.a(new_n188), .b(new_n185), .out0(new_n189));
  xorc02aa1n12x5               g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  aob012aa1n02x5               g095(.a(new_n186), .b(new_n167), .c(new_n169), .out0(new_n191));
  aoi012aa1n02x5               g096(.a(new_n190), .b(new_n178), .c(new_n179), .o1(new_n192));
  aoi022aa1n02x5               g097(.a(new_n191), .b(new_n192), .c(new_n190), .d(new_n189), .o1(\s[17] ));
  nor042aa1n03x5               g098(.a(\b[17] ), .b(\a[18] ), .o1(new_n194));
  inv040aa1d32x5               g099(.a(\a[17] ), .o1(new_n195));
  inv040aa1n20x5               g100(.a(\b[16] ), .o1(new_n196));
  nanp02aa1n12x5               g101(.a(new_n196), .b(new_n195), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  oaib12aa1n02x5               g103(.a(new_n197), .b(new_n194), .c(new_n198), .out0(new_n199));
  aoi012aa1n02x5               g104(.a(new_n199), .b(new_n189), .c(new_n190), .o1(new_n200));
  nano22aa1n12x5               g105(.a(new_n194), .b(new_n190), .c(new_n198), .out0(new_n201));
  oaoi03aa1n12x5               g106(.a(\a[18] ), .b(\b[17] ), .c(new_n197), .o1(new_n202));
  aoi012aa1n06x5               g107(.a(new_n202), .b(new_n189), .c(new_n201), .o1(new_n203));
  oab012aa1n03x5               g108(.a(new_n200), .b(new_n203), .c(new_n194), .out0(\s[18] ));
  nor002aa1d32x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  inv040aa1n02x5               g110(.a(new_n205), .o1(new_n206));
  nand42aa1d28x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n203), .b(new_n207), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g114(.a(new_n205), .b(new_n207), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n04x5               g116(.a(new_n211), .b(new_n202), .c(new_n189), .d(new_n201), .o1(new_n212));
  nor042aa1n06x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand42aa1d28x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  norb03aa1n02x5               g120(.a(new_n214), .b(new_n205), .c(new_n213), .out0(new_n216));
  nanp02aa1n03x5               g121(.a(new_n212), .b(new_n216), .o1(new_n217));
  aoai13aa1n03x5               g122(.a(new_n217), .b(new_n215), .c(new_n206), .d(new_n212), .o1(\s[20] ));
  nano23aa1n09x5               g123(.a(new_n205), .b(new_n213), .c(new_n214), .d(new_n207), .out0(new_n219));
  nand02aa1d04x5               g124(.a(new_n201), .b(new_n219), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n188), .c(new_n129), .d(new_n184), .o1(new_n222));
  oaoi03aa1n03x5               g127(.a(\a[20] ), .b(\b[19] ), .c(new_n206), .o1(new_n223));
  aoi012aa1n02x5               g128(.a(new_n223), .b(new_n219), .c(new_n202), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xnbna2aa1n03x5               g130(.a(new_n225), .b(new_n222), .c(new_n224), .out0(\s[21] ));
  nor042aa1n12x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aob012aa1n03x5               g133(.a(new_n225), .b(new_n222), .c(new_n224), .out0(new_n229));
  xorc02aa1n02x5               g134(.a(\a[22] ), .b(\b[21] ), .out0(new_n230));
  nand02aa1d06x5               g135(.a(\b[21] ), .b(\a[22] ), .o1(new_n231));
  oai022aa1n02x5               g136(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n231), .b(new_n232), .out0(new_n233));
  nand02aa1n04x5               g138(.a(new_n229), .b(new_n233), .o1(new_n234));
  aoai13aa1n03x5               g139(.a(new_n234), .b(new_n230), .c(new_n228), .d(new_n229), .o1(\s[22] ));
  nanp02aa1n02x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nor042aa1n02x5               g141(.a(\b[21] ), .b(\a[22] ), .o1(new_n237));
  nano23aa1n06x5               g142(.a(new_n227), .b(new_n237), .c(new_n231), .d(new_n236), .out0(new_n238));
  and003aa1n02x5               g143(.a(new_n201), .b(new_n238), .c(new_n219), .o(new_n239));
  aoai13aa1n06x5               g144(.a(new_n238), .b(new_n223), .c(new_n219), .d(new_n202), .o1(new_n240));
  oaih12aa1n06x5               g145(.a(new_n231), .b(new_n237), .c(new_n227), .o1(new_n241));
  nanp02aa1n02x5               g146(.a(new_n240), .b(new_n241), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[22] ), .b(\a[23] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n242), .c(new_n189), .d(new_n239), .o1(new_n245));
  aoi112aa1n02x7               g150(.a(new_n244), .b(new_n242), .c(new_n189), .d(new_n239), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n245), .b(new_n246), .out0(\s[23] ));
  norp02aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[24] ), .b(\b[23] ), .out0(new_n250));
  nanp02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  oai022aa1n02x5               g156(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(new_n253));
  nand02aa1n02x5               g158(.a(new_n245), .b(new_n253), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n250), .c(new_n249), .d(new_n245), .o1(\s[24] ));
  norb02aa1n09x5               g160(.a(new_n250), .b(new_n243), .out0(new_n256));
  nano22aa1n02x5               g161(.a(new_n220), .b(new_n256), .c(new_n238), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n188), .c(new_n129), .d(new_n184), .o1(new_n258));
  inv040aa1n04x5               g163(.a(new_n256), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(new_n252), .b(new_n251), .o1(new_n260));
  aoai13aa1n12x5               g165(.a(new_n260), .b(new_n259), .c(new_n240), .d(new_n241), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  tech160nm_fixorc02aa1n03p5x5 g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  xnbna2aa1n03x5               g168(.a(new_n263), .b(new_n258), .c(new_n262), .out0(\s[25] ));
  norp02aa1n02x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  aob012aa1n03x5               g171(.a(new_n263), .b(new_n258), .c(new_n262), .out0(new_n267));
  tech160nm_fixorc02aa1n03p5x5 g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  nanp02aa1n02x5               g173(.a(\b[25] ), .b(\a[26] ), .o1(new_n269));
  oai022aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n269), .b(new_n270), .out0(new_n271));
  nand02aa1n03x5               g176(.a(new_n267), .b(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n268), .c(new_n266), .d(new_n267), .o1(\s[26] ));
  and002aa1n02x5               g178(.a(new_n268), .b(new_n263), .o(new_n274));
  nano32aa1n03x7               g179(.a(new_n220), .b(new_n274), .c(new_n238), .d(new_n256), .out0(new_n275));
  aoai13aa1n12x5               g180(.a(new_n275), .b(new_n188), .c(new_n129), .d(new_n184), .o1(new_n276));
  aoi022aa1n09x5               g181(.a(new_n261), .b(new_n274), .c(new_n269), .d(new_n270), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n277), .c(new_n276), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  nand02aa1n04x5               g186(.a(new_n261), .b(new_n274), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(new_n270), .b(new_n269), .o1(new_n283));
  nanp03aa1d12x5               g188(.a(new_n282), .b(new_n276), .c(new_n283), .o1(new_n284));
  nanp02aa1n03x5               g189(.a(new_n284), .b(new_n278), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .out0(new_n286));
  inv000aa1d42x5               g191(.a(new_n278), .o1(new_n287));
  oai022aa1n02x5               g192(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n288));
  aoi012aa1n02x5               g193(.a(new_n288), .b(\a[28] ), .c(\b[27] ), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n287), .c(new_n277), .d(new_n276), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n286), .c(new_n285), .d(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g196(.a(new_n286), .b(new_n278), .o(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  oaib12aa1n09x5               g199(.a(new_n288), .b(new_n294), .c(\a[28] ), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  tech160nm_fixorc02aa1n03p5x5 g201(.a(\a[29] ), .b(\b[28] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n297), .b(new_n296), .out0(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n293), .c(new_n277), .d(new_n276), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n297), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n284), .d(new_n292), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n301), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g208(.a(new_n300), .b(new_n278), .c(new_n286), .out0(new_n304));
  oaoi03aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .o1(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n305), .c(new_n284), .d(new_n304), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n304), .o1(new_n308));
  norp02aa1n02x5               g213(.a(new_n305), .b(new_n306), .o1(new_n309));
  aoai13aa1n02x5               g214(.a(new_n309), .b(new_n308), .c(new_n277), .d(new_n276), .o1(new_n310));
  nanp02aa1n03x5               g215(.a(new_n307), .b(new_n310), .o1(\s[30] ));
  nano32aa1n03x7               g216(.a(new_n306), .b(new_n297), .c(new_n286), .d(new_n278), .out0(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  aoi012aa1n02x5               g218(.a(new_n309), .b(\a[30] ), .c(\b[29] ), .o1(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  norp02aa1n02x5               g220(.a(new_n314), .b(new_n315), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n313), .c(new_n277), .d(new_n276), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n315), .b(new_n314), .c(new_n284), .d(new_n312), .o1(new_n318));
  nanp02aa1n03x5               g223(.a(new_n318), .b(new_n317), .o1(\s[31] ));
  xorb03aa1n02x5               g224(.a(new_n105), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g225(.a(new_n112), .b(new_n113), .o1(new_n321));
  oaoi13aa1n02x5               g226(.a(new_n108), .b(new_n110), .c(new_n105), .d(new_n109), .o1(new_n322));
  aoib12aa1n02x5               g227(.a(new_n322), .b(new_n321), .c(new_n106), .out0(\s[4] ));
  xorb03aa1n02x5               g228(.a(new_n321), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g229(.a(new_n121), .b(new_n321), .c(new_n122), .o1(new_n325));
  xnrb03aa1n02x5               g230(.a(new_n325), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g231(.a(new_n126), .b(new_n321), .c(new_n123), .o(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g233(.a(new_n116), .b(new_n327), .c(new_n117), .o1(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g235(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


