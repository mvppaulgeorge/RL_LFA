// Benchmark "adder" written by ABC on Wed Jul 17 23:22:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n313, new_n315, new_n318, new_n319,
    new_n321, new_n322, new_n323, new_n325;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(new_n98), .o1(new_n99));
  norp02aa1n04x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor022aa1n12x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  inv000aa1n06x5               g006(.a(new_n101), .o1(new_n102));
  oaoi03aa1n06x5               g007(.a(\a[8] ), .b(\b[7] ), .c(new_n102), .o1(new_n103));
  inv000aa1n02x5               g008(.a(new_n103), .o1(new_n104));
  norp02aa1n12x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  oab012aa1n12x5               g010(.a(new_n105), .b(\a[5] ), .c(\b[4] ), .out0(new_n106));
  and002aa1n06x5               g011(.a(\b[5] ), .b(\a[6] ), .o(new_n107));
  nanp02aa1n04x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor022aa1n08x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nanp02aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nona23aa1n09x5               g015(.a(new_n108), .b(new_n110), .c(new_n101), .d(new_n109), .out0(new_n111));
  oai013aa1n03x5               g016(.a(new_n104), .b(new_n111), .c(new_n106), .d(new_n107), .o1(new_n112));
  nor042aa1d18x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  inv040aa1n02x5               g018(.a(new_n113), .o1(new_n114));
  oao003aa1n09x5               g019(.a(\a[4] ), .b(\b[3] ), .c(new_n114), .carry(new_n115));
  tech160nm_fixnrc02aa1n04x5   g020(.a(\b[3] ), .b(\a[4] ), .out0(new_n116));
  nand02aa1d28x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  nand42aa1d28x5               g022(.a(\b[2] ), .b(\a[3] ), .o1(new_n118));
  nanb03aa1d18x5               g023(.a(new_n113), .b(new_n118), .c(new_n117), .out0(new_n119));
  nand22aa1n06x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  nor002aa1n04x5               g025(.a(\b[1] ), .b(\a[2] ), .o1(new_n121));
  norb03aa1n09x5               g026(.a(new_n117), .b(new_n121), .c(new_n120), .out0(new_n122));
  oai013aa1d12x5               g027(.a(new_n115), .b(new_n122), .c(new_n119), .d(new_n116), .o1(new_n123));
  xnrc02aa1n02x5               g028(.a(\b[5] ), .b(\a[6] ), .out0(new_n124));
  xnrc02aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .out0(new_n125));
  nor043aa1n03x5               g030(.a(new_n111), .b(new_n124), .c(new_n125), .o1(new_n126));
  nand02aa1d06x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n100), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n112), .c(new_n123), .d(new_n126), .o1(new_n129));
  obai22aa1n02x7               g034(.a(new_n129), .b(new_n100), .c(new_n97), .d(new_n99), .out0(new_n130));
  nona32aa1n02x4               g035(.a(new_n129), .b(new_n100), .c(new_n99), .d(new_n97), .out0(new_n131));
  nanp02aa1n02x5               g036(.a(new_n130), .b(new_n131), .o1(\s[10] ));
  xnrc02aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n133), .b(new_n131), .c(new_n98), .out0(\s[11] ));
  inv000aa1d42x5               g039(.a(\a[11] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(\b[10] ), .o1(new_n136));
  nand02aa1d08x5               g041(.a(new_n136), .b(new_n135), .o1(new_n137));
  nona22aa1n02x4               g042(.a(new_n131), .b(new_n133), .c(new_n99), .out0(new_n138));
  norp02aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  and002aa1n03x5               g044(.a(\b[11] ), .b(\a[12] ), .o(new_n140));
  norp02aa1n02x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n138), .c(new_n137), .out0(\s[12] ));
  inv000aa1d42x5               g047(.a(new_n106), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n107), .o1(new_n144));
  nano23aa1n03x7               g049(.a(new_n101), .b(new_n109), .c(new_n110), .d(new_n108), .out0(new_n145));
  aoi013aa1n06x4               g050(.a(new_n103), .b(new_n145), .c(new_n144), .d(new_n143), .o1(new_n146));
  nanp02aa1n02x5               g051(.a(new_n123), .b(new_n126), .o1(new_n147));
  nano23aa1n06x5               g052(.a(new_n97), .b(new_n100), .c(new_n127), .d(new_n98), .out0(new_n148));
  aoi112aa1n06x5               g053(.a(new_n140), .b(new_n139), .c(\a[11] ), .d(\b[10] ), .o1(new_n149));
  nand23aa1n03x5               g054(.a(new_n148), .b(new_n137), .c(new_n149), .o1(new_n150));
  oai022aa1n02x5               g055(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n151));
  aoi022aa1n02x5               g056(.a(new_n135), .b(new_n136), .c(\a[10] ), .d(\b[9] ), .o1(new_n152));
  oaoi03aa1n09x5               g057(.a(\a[12] ), .b(\b[11] ), .c(new_n137), .o1(new_n153));
  aoi013aa1n03x5               g058(.a(new_n153), .b(new_n149), .c(new_n151), .d(new_n152), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n150), .c(new_n147), .d(new_n146), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nanp02aa1n24x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  aoi012aa1n02x5               g063(.a(new_n157), .b(new_n155), .c(new_n158), .o1(new_n159));
  xnrb03aa1n03x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand42aa1n08x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nano23aa1d15x5               g067(.a(new_n157), .b(new_n161), .c(new_n162), .d(new_n158), .out0(new_n163));
  oa0012aa1n06x5               g068(.a(new_n162), .b(new_n161), .c(new_n157), .o(new_n164));
  xorc02aa1n12x5               g069(.a(\a[15] ), .b(\b[14] ), .out0(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n164), .c(new_n155), .d(new_n163), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n165), .b(new_n164), .c(new_n155), .d(new_n163), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(\s[15] ));
  orn002aa1n02x5               g073(.a(\a[15] ), .b(\b[14] ), .o(new_n169));
  xorc02aa1n12x5               g074(.a(\a[16] ), .b(\b[15] ), .out0(new_n170));
  aobi12aa1n02x5               g075(.a(new_n170), .b(new_n166), .c(new_n169), .out0(new_n171));
  norp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nona22aa1n02x4               g077(.a(new_n166), .b(new_n170), .c(new_n172), .out0(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n171), .out0(\s[16] ));
  nand23aa1n04x5               g079(.a(new_n163), .b(new_n165), .c(new_n170), .o1(new_n175));
  nor042aa1n03x5               g080(.a(new_n175), .b(new_n150), .o1(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n112), .c(new_n123), .d(new_n126), .o1(new_n177));
  nand43aa1n02x5               g082(.a(new_n164), .b(new_n165), .c(new_n170), .o1(new_n178));
  nanp03aa1n02x5               g083(.a(new_n149), .b(new_n151), .c(new_n152), .o1(new_n179));
  inv000aa1n02x5               g084(.a(new_n153), .o1(new_n180));
  aoi012aa1n02x7               g085(.a(new_n175), .b(new_n179), .c(new_n180), .o1(new_n181));
  oao003aa1n02x5               g086(.a(\a[16] ), .b(\b[15] ), .c(new_n169), .carry(new_n182));
  nano22aa1n03x7               g087(.a(new_n181), .b(new_n178), .c(new_n182), .out0(new_n183));
  nand02aa1d06x5               g088(.a(new_n177), .b(new_n183), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g090(.a(\a[18] ), .o1(new_n186));
  inv040aa1d32x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  oaoi03aa1n03x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n186), .out0(\s[18] ));
  xroi22aa1d04x5               g095(.a(new_n187), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(new_n188), .b(new_n187), .o1(new_n192));
  oaoi03aa1n12x5               g097(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n193));
  nor042aa1n09x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand02aa1n06x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  aoai13aa1n06x5               g101(.a(new_n196), .b(new_n193), .c(new_n184), .d(new_n191), .o1(new_n197));
  aoi112aa1n02x5               g102(.a(new_n196), .b(new_n193), .c(new_n184), .d(new_n191), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n197), .b(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n12x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand42aa1n06x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  oaoi13aa1n06x5               g109(.a(new_n204), .b(new_n197), .c(\a[19] ), .d(\b[18] ), .o1(new_n205));
  nona22aa1n02x5               g110(.a(new_n197), .b(new_n203), .c(new_n194), .out0(new_n206));
  norb02aa1n03x4               g111(.a(new_n206), .b(new_n205), .out0(\s[20] ));
  nano23aa1n09x5               g112(.a(new_n194), .b(new_n201), .c(new_n202), .d(new_n195), .out0(new_n208));
  nanp02aa1n02x5               g113(.a(new_n191), .b(new_n208), .o1(new_n209));
  oai022aa1n04x7               g114(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n210));
  oaib12aa1n06x5               g115(.a(new_n210), .b(new_n186), .c(\b[17] ), .out0(new_n211));
  nona23aa1d18x5               g116(.a(new_n202), .b(new_n195), .c(new_n194), .d(new_n201), .out0(new_n212));
  oai012aa1n12x5               g117(.a(new_n202), .b(new_n201), .c(new_n194), .o1(new_n213));
  oai012aa1d24x5               g118(.a(new_n213), .b(new_n212), .c(new_n211), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n215), .b(new_n209), .c(new_n177), .d(new_n183), .o1(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  xorc02aa1n02x5               g123(.a(\a[21] ), .b(\b[20] ), .out0(new_n219));
  xorc02aa1n02x5               g124(.a(\a[22] ), .b(\b[21] ), .out0(new_n220));
  aoai13aa1n03x5               g125(.a(new_n220), .b(new_n218), .c(new_n216), .d(new_n219), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(new_n218), .b(new_n220), .c(new_n216), .d(new_n219), .o1(new_n222));
  norb02aa1n02x7               g127(.a(new_n221), .b(new_n222), .out0(\s[22] ));
  inv000aa1d42x5               g128(.a(\a[21] ), .o1(new_n224));
  inv040aa1d32x5               g129(.a(\a[22] ), .o1(new_n225));
  xroi22aa1d06x4               g130(.a(new_n224), .b(\b[20] ), .c(new_n225), .d(\b[21] ), .out0(new_n226));
  and003aa1n02x5               g131(.a(new_n191), .b(new_n226), .c(new_n208), .o(new_n227));
  inv040aa1n03x5               g132(.a(new_n213), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n226), .b(new_n228), .c(new_n208), .d(new_n193), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\b[21] ), .o1(new_n230));
  oao003aa1n02x5               g135(.a(new_n225), .b(new_n230), .c(new_n218), .carry(new_n231));
  inv000aa1n02x5               g136(.a(new_n231), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(new_n229), .b(new_n232), .o1(new_n233));
  xorc02aa1n02x5               g138(.a(\a[23] ), .b(\b[22] ), .out0(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n233), .c(new_n184), .d(new_n227), .o1(new_n235));
  aoi112aa1n02x5               g140(.a(new_n234), .b(new_n233), .c(new_n184), .d(new_n227), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n235), .b(new_n236), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  xorc02aa1n02x5               g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  aobi12aa1n06x5               g145(.a(new_n240), .b(new_n235), .c(new_n239), .out0(new_n241));
  nona22aa1n02x5               g146(.a(new_n235), .b(new_n240), .c(new_n238), .out0(new_n242));
  norb02aa1n03x4               g147(.a(new_n242), .b(new_n241), .out0(\s[24] ));
  inv000aa1d42x5               g148(.a(\a[23] ), .o1(new_n244));
  inv020aa1n04x5               g149(.a(\a[24] ), .o1(new_n245));
  xroi22aa1d06x4               g150(.a(new_n244), .b(\b[22] ), .c(new_n245), .d(\b[23] ), .out0(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  oao003aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .c(new_n239), .carry(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n247), .c(new_n229), .d(new_n232), .o1(new_n249));
  nano22aa1n02x4               g154(.a(new_n209), .b(new_n226), .c(new_n246), .out0(new_n250));
  xorc02aa1n02x5               g155(.a(\a[25] ), .b(\b[24] ), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n249), .c(new_n184), .d(new_n250), .o1(new_n252));
  aoi112aa1n02x5               g157(.a(new_n249), .b(new_n251), .c(new_n184), .d(new_n250), .o1(new_n253));
  norb02aa1n02x5               g158(.a(new_n252), .b(new_n253), .out0(\s[25] ));
  nor042aa1n03x5               g159(.a(\b[24] ), .b(\a[25] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  xorc02aa1n02x5               g161(.a(\a[26] ), .b(\b[25] ), .out0(new_n257));
  aobi12aa1n06x5               g162(.a(new_n257), .b(new_n252), .c(new_n256), .out0(new_n258));
  nona22aa1n03x5               g163(.a(new_n252), .b(new_n257), .c(new_n255), .out0(new_n259));
  norb02aa1n03x4               g164(.a(new_n259), .b(new_n258), .out0(\s[26] ));
  xorc02aa1n02x5               g165(.a(\a[4] ), .b(\b[3] ), .out0(new_n261));
  nona22aa1n03x5               g166(.a(new_n117), .b(new_n121), .c(new_n120), .out0(new_n262));
  nanb03aa1n06x5               g167(.a(new_n119), .b(new_n262), .c(new_n261), .out0(new_n263));
  nona22aa1n02x4               g168(.a(new_n145), .b(new_n125), .c(new_n124), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n146), .b(new_n264), .c(new_n263), .d(new_n115), .o1(new_n265));
  oai112aa1n02x5               g170(.a(new_n178), .b(new_n182), .c(new_n154), .d(new_n175), .o1(new_n266));
  inv000aa1d42x5               g171(.a(\a[25] ), .o1(new_n267));
  inv020aa1n04x5               g172(.a(\a[26] ), .o1(new_n268));
  xroi22aa1d06x4               g173(.a(new_n267), .b(\b[24] ), .c(new_n268), .d(\b[25] ), .out0(new_n269));
  nano32aa1n03x7               g174(.a(new_n209), .b(new_n269), .c(new_n226), .d(new_n246), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n266), .c(new_n265), .d(new_n176), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[26] ), .b(\b[25] ), .c(new_n256), .carry(new_n272));
  aobi12aa1n06x5               g177(.a(new_n272), .b(new_n249), .c(new_n269), .out0(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n271), .out0(\s[27] ));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  inv040aa1n03x5               g181(.a(new_n276), .o1(new_n277));
  aobi12aa1n06x5               g182(.a(new_n270), .b(new_n177), .c(new_n183), .out0(new_n278));
  aoai13aa1n04x5               g183(.a(new_n246), .b(new_n231), .c(new_n214), .d(new_n226), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n269), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n272), .b(new_n280), .c(new_n279), .d(new_n248), .o1(new_n281));
  oaih12aa1n02x5               g186(.a(new_n274), .b(new_n281), .c(new_n278), .o1(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n283), .b(new_n282), .c(new_n277), .o1(new_n284));
  aobi12aa1n02x7               g189(.a(new_n274), .b(new_n273), .c(new_n271), .out0(new_n285));
  nano22aa1n03x5               g190(.a(new_n285), .b(new_n277), .c(new_n283), .out0(new_n286));
  norp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n274), .b(new_n283), .out0(new_n288));
  oaih12aa1n02x5               g193(.a(new_n288), .b(new_n281), .c(new_n278), .o1(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n277), .carry(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n291), .b(new_n289), .c(new_n290), .o1(new_n292));
  aobi12aa1n02x7               g197(.a(new_n288), .b(new_n273), .c(new_n271), .out0(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n291), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g201(.a(new_n274), .b(new_n291), .c(new_n283), .out0(new_n297));
  oaih12aa1n02x5               g202(.a(new_n297), .b(new_n281), .c(new_n278), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[29] ), .b(\a[30] ), .out0(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n300), .b(new_n298), .c(new_n299), .o1(new_n301));
  aobi12aa1n02x7               g206(.a(new_n297), .b(new_n273), .c(new_n271), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n299), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[30] ));
  norb02aa1n02x5               g209(.a(new_n297), .b(new_n300), .out0(new_n305));
  aobi12aa1n02x7               g210(.a(new_n305), .b(new_n273), .c(new_n271), .out0(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  nano22aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n308), .out0(new_n309));
  oaih12aa1n02x5               g214(.a(new_n305), .b(new_n281), .c(new_n278), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n308), .b(new_n310), .c(new_n307), .o1(new_n311));
  norp02aa1n03x5               g216(.a(new_n311), .b(new_n309), .o1(\s[31] ));
  aoi022aa1n02x5               g217(.a(new_n262), .b(new_n117), .c(new_n114), .d(new_n118), .o1(new_n313));
  aoib12aa1n02x5               g218(.a(new_n313), .b(new_n262), .c(new_n119), .out0(\s[3] ));
  oai012aa1n02x5               g219(.a(new_n114), .b(new_n122), .c(new_n119), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g221(.a(new_n123), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  orn002aa1n02x5               g222(.a(\a[5] ), .b(\b[4] ), .o(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n125), .c(new_n263), .d(new_n115), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g225(.a(new_n110), .b(new_n101), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n105), .c(new_n319), .d(new_n144), .o1(new_n322));
  aoi112aa1n02x5               g227(.a(new_n321), .b(new_n105), .c(new_n319), .d(new_n144), .o1(new_n323));
  norb02aa1n02x5               g228(.a(new_n322), .b(new_n323), .out0(\s[7] ));
  norb02aa1n02x5               g229(.a(new_n108), .b(new_n109), .out0(new_n325));
  xnbna2aa1n03x5               g230(.a(new_n325), .b(new_n322), .c(new_n102), .out0(\s[8] ));
  xorb03aa1n02x5               g231(.a(new_n265), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


