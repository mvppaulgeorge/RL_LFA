// Benchmark "adder" written by ABC on Thu Jul 18 02:09:55 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n330,
    new_n332, new_n335, new_n337, new_n339, new_n340, new_n341, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand22aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nanp02aa1n06x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nor042aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  oai112aa1n06x5               g007(.a(new_n102), .b(new_n100), .c(new_n101), .d(new_n99), .o1(new_n103));
  oa0022aa1n06x5               g008(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n104));
  aoi022aa1d18x5               g009(.a(new_n103), .b(new_n104), .c(\b[3] ), .d(\a[4] ), .o1(new_n105));
  nor022aa1n08x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand02aa1n06x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand02aa1n04x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nona23aa1d18x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .out0(new_n111));
  tech160nm_fixnrc02aa1n04x5   g016(.a(\b[4] ), .b(\a[5] ), .out0(new_n112));
  nor043aa1n06x5               g017(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n113));
  inv000aa1d42x5               g018(.a(\a[6] ), .o1(new_n114));
  inv000aa1d42x5               g019(.a(\b[5] ), .o1(new_n115));
  nor042aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  tech160nm_fioaoi03aa1n03p5x5 g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  inv040aa1d30x5               g022(.a(new_n108), .o1(new_n118));
  oaoi03aa1n09x5               g023(.a(\a[8] ), .b(\b[7] ), .c(new_n118), .o1(new_n119));
  oabi12aa1n06x5               g024(.a(new_n119), .b(new_n110), .c(new_n117), .out0(new_n120));
  nand02aa1n12x5               g025(.a(\b[8] ), .b(\a[9] ), .o1(new_n121));
  norb02aa1n02x5               g026(.a(new_n121), .b(new_n97), .out0(new_n122));
  aoai13aa1n06x5               g027(.a(new_n122), .b(new_n120), .c(new_n113), .d(new_n105), .o1(new_n123));
  nor002aa1d24x5               g028(.a(\b[9] ), .b(\a[10] ), .o1(new_n124));
  nand02aa1d28x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n126), .b(new_n123), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(new_n124), .o1(new_n128));
  inv000aa1n02x5               g033(.a(new_n126), .o1(new_n129));
  aoai13aa1n06x5               g034(.a(new_n128), .b(new_n129), .c(new_n123), .d(new_n98), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1d18x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1d28x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  nor042aa1d18x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nand42aa1d28x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  aoai13aa1n03x5               g043(.a(new_n138), .b(new_n132), .c(new_n130), .d(new_n134), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n130), .b(new_n134), .o1(new_n140));
  nona22aa1n02x4               g045(.a(new_n140), .b(new_n138), .c(new_n132), .out0(new_n141));
  nanp02aa1n02x5               g046(.a(new_n141), .b(new_n139), .o1(\s[12] ));
  nano23aa1n09x5               g047(.a(new_n132), .b(new_n135), .c(new_n136), .d(new_n133), .out0(new_n143));
  nano23aa1n09x5               g048(.a(new_n97), .b(new_n124), .c(new_n125), .d(new_n121), .out0(new_n144));
  nand22aa1n09x5               g049(.a(new_n144), .b(new_n143), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  aoai13aa1n06x5               g051(.a(new_n146), .b(new_n120), .c(new_n113), .d(new_n105), .o1(new_n147));
  aoi012aa1n06x5               g052(.a(new_n124), .b(new_n97), .c(new_n125), .o1(new_n148));
  inv020aa1n04x5               g053(.a(new_n148), .o1(new_n149));
  tech160nm_fioai012aa1n03p5x5 g054(.a(new_n136), .b(new_n135), .c(new_n132), .o1(new_n150));
  aobi12aa1n06x5               g055(.a(new_n150), .b(new_n143), .c(new_n149), .out0(new_n151));
  nor002aa1d32x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1n08x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  norb02aa1n03x5               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  xnbna2aa1n03x5               g059(.a(new_n154), .b(new_n147), .c(new_n151), .out0(\s[13] ));
  orn002aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .o(new_n156));
  nanp02aa1n02x5               g061(.a(\b[3] ), .b(\a[4] ), .o1(new_n157));
  nanp02aa1n03x5               g062(.a(new_n103), .b(new_n104), .o1(new_n158));
  nanp02aa1n03x5               g063(.a(new_n158), .b(new_n157), .o1(new_n159));
  nano23aa1n02x5               g064(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n160));
  xorc02aa1n02x5               g065(.a(\a[6] ), .b(\b[5] ), .out0(new_n161));
  xorc02aa1n02x5               g066(.a(\a[5] ), .b(\b[4] ), .out0(new_n162));
  nand03aa1n02x5               g067(.a(new_n160), .b(new_n161), .c(new_n162), .o1(new_n163));
  oab012aa1n06x5               g068(.a(new_n119), .b(new_n110), .c(new_n117), .out0(new_n164));
  tech160nm_fioai012aa1n03p5x5 g069(.a(new_n164), .b(new_n159), .c(new_n163), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n136), .b(new_n133), .c(new_n132), .d(new_n135), .out0(new_n166));
  oai012aa1n06x5               g071(.a(new_n150), .b(new_n166), .c(new_n148), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n154), .b(new_n167), .c(new_n165), .d(new_n146), .o1(new_n168));
  nor002aa1d32x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1d28x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n03x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n168), .c(new_n156), .out0(\s[14] ));
  nona23aa1n09x5               g077(.a(new_n170), .b(new_n153), .c(new_n152), .d(new_n169), .out0(new_n173));
  aoi012aa1n02x5               g078(.a(new_n169), .b(new_n152), .c(new_n170), .o1(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n173), .c(new_n147), .d(new_n151), .o1(new_n175));
  xorb03aa1n02x5               g080(.a(new_n175), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n16x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand22aa1n09x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nor022aa1n08x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand02aa1n12x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  aoai13aa1n03x5               g086(.a(new_n181), .b(new_n177), .c(new_n175), .d(new_n178), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n178), .b(new_n177), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n175), .b(new_n183), .o1(new_n184));
  nona22aa1n02x4               g089(.a(new_n184), .b(new_n181), .c(new_n177), .out0(new_n185));
  nanp02aa1n03x5               g090(.a(new_n185), .b(new_n182), .o1(\s[16] ));
  nano23aa1n06x5               g091(.a(new_n177), .b(new_n179), .c(new_n180), .d(new_n178), .out0(new_n187));
  nano32aa1d12x5               g092(.a(new_n145), .b(new_n187), .c(new_n154), .d(new_n171), .out0(new_n188));
  aoai13aa1n12x5               g093(.a(new_n188), .b(new_n120), .c(new_n105), .d(new_n113), .o1(new_n189));
  nona23aa1n03x5               g094(.a(new_n180), .b(new_n178), .c(new_n177), .d(new_n179), .out0(new_n190));
  nor002aa1n04x5               g095(.a(new_n190), .b(new_n173), .o1(new_n191));
  aoai13aa1n04x5               g096(.a(new_n178), .b(new_n169), .c(new_n152), .d(new_n170), .o1(new_n192));
  nona22aa1n03x5               g097(.a(new_n192), .b(new_n179), .c(new_n177), .out0(new_n193));
  aoi022aa1d18x5               g098(.a(new_n167), .b(new_n191), .c(new_n180), .d(new_n193), .o1(new_n194));
  xnrc02aa1n02x5               g099(.a(\b[16] ), .b(\a[17] ), .out0(new_n195));
  xobna2aa1n03x5               g100(.a(new_n195), .b(new_n189), .c(new_n194), .out0(\s[17] ));
  nanp02aa1n03x5               g101(.a(new_n113), .b(new_n105), .o1(new_n197));
  nona23aa1n03x5               g102(.a(new_n187), .b(new_n144), .c(new_n166), .d(new_n173), .out0(new_n198));
  aoai13aa1n12x5               g103(.a(new_n194), .b(new_n198), .c(new_n197), .d(new_n164), .o1(new_n199));
  nor042aa1d18x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  nand42aa1d28x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  nor002aa1n20x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand42aa1d28x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  aoai13aa1n03x5               g109(.a(new_n204), .b(new_n200), .c(new_n199), .d(new_n201), .o1(new_n205));
  aoi112aa1n02x7               g110(.a(new_n200), .b(new_n204), .c(new_n199), .d(new_n201), .o1(new_n206));
  norb02aa1n03x4               g111(.a(new_n205), .b(new_n206), .out0(\s[18] ));
  nano23aa1d15x5               g112(.a(new_n200), .b(new_n202), .c(new_n203), .d(new_n201), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoi012aa1d18x5               g114(.a(new_n202), .b(new_n200), .c(new_n203), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n209), .c(new_n189), .d(new_n194), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1d18x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nand42aa1n16x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  xnrc02aa1n12x5               g120(.a(\b[19] ), .b(\a[20] ), .out0(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n214), .c(new_n211), .d(new_n215), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n210), .o1(new_n218));
  nanb02aa1n18x5               g123(.a(new_n214), .b(new_n215), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n220), .b(new_n218), .c(new_n199), .d(new_n208), .o1(new_n221));
  nona22aa1n03x5               g126(.a(new_n221), .b(new_n216), .c(new_n214), .out0(new_n222));
  nanp02aa1n03x5               g127(.a(new_n217), .b(new_n222), .o1(\s[20] ));
  nona22aa1d36x5               g128(.a(new_n208), .b(new_n216), .c(new_n219), .out0(new_n224));
  inv000aa1d42x5               g129(.a(\b[19] ), .o1(new_n225));
  norp02aa1n02x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n215), .b(new_n202), .c(new_n200), .d(new_n203), .o1(new_n227));
  nona22aa1n06x5               g132(.a(new_n227), .b(new_n226), .c(new_n214), .out0(new_n228));
  oaib12aa1n18x5               g133(.a(new_n228), .b(new_n225), .c(\a[20] ), .out0(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n224), .c(new_n189), .d(new_n194), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[20] ), .b(\a[21] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  nor022aa1n06x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  nanp02aa1n06x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  nanb02aa1n09x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n232), .c(new_n230), .d(new_n234), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n224), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n229), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n234), .b(new_n240), .c(new_n199), .d(new_n239), .o1(new_n241));
  nona22aa1n03x5               g146(.a(new_n241), .b(new_n237), .c(new_n232), .out0(new_n242));
  nanp02aa1n03x5               g147(.a(new_n238), .b(new_n242), .o1(\s[22] ));
  nor042aa1n12x5               g148(.a(new_n233), .b(new_n237), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  nor042aa1n04x5               g150(.a(new_n224), .b(new_n245), .o1(new_n246));
  inv020aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  aoi012aa1n02x7               g152(.a(new_n235), .b(new_n232), .c(new_n236), .o1(new_n248));
  oa0012aa1n06x5               g153(.a(new_n248), .b(new_n229), .c(new_n245), .o(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n247), .c(new_n189), .d(new_n194), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  xnrc02aa1n12x5               g157(.a(\b[22] ), .b(\a[23] ), .out0(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[23] ), .b(\a[24] ), .out0(new_n255));
  aoai13aa1n03x5               g160(.a(new_n255), .b(new_n252), .c(new_n250), .d(new_n254), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n249), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n254), .b(new_n257), .c(new_n199), .d(new_n246), .o1(new_n258));
  nona22aa1n03x5               g163(.a(new_n258), .b(new_n255), .c(new_n252), .out0(new_n259));
  nanp02aa1n03x5               g164(.a(new_n256), .b(new_n259), .o1(\s[24] ));
  nor042aa1n03x5               g165(.a(new_n255), .b(new_n253), .o1(new_n261));
  nano22aa1n03x7               g166(.a(new_n224), .b(new_n261), .c(new_n244), .out0(new_n262));
  inv020aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  nand02aa1d06x5               g168(.a(new_n261), .b(new_n244), .o1(new_n264));
  orn002aa1n02x5               g169(.a(\a[24] ), .b(\b[23] ), .o(new_n265));
  aob012aa1n02x5               g170(.a(new_n252), .b(\b[23] ), .c(\a[24] ), .out0(new_n266));
  nor003aa1n02x5               g171(.a(new_n255), .b(new_n253), .c(new_n248), .o1(new_n267));
  nano22aa1n03x7               g172(.a(new_n267), .b(new_n265), .c(new_n266), .out0(new_n268));
  oai012aa1n18x5               g173(.a(new_n268), .b(new_n229), .c(new_n264), .o1(new_n269));
  inv040aa1n04x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n263), .c(new_n189), .d(new_n194), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  tech160nm_fixorc02aa1n04x5   g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  xnrc02aa1n12x5               g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  aoai13aa1n03x5               g180(.a(new_n275), .b(new_n273), .c(new_n271), .d(new_n274), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n274), .b(new_n269), .c(new_n199), .d(new_n262), .o1(new_n277));
  nona22aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .out0(new_n278));
  nanp02aa1n03x5               g183(.a(new_n276), .b(new_n278), .o1(\s[26] ));
  nanp02aa1n02x5               g184(.a(new_n193), .b(new_n180), .o1(new_n280));
  oaib12aa1n02x5               g185(.a(new_n280), .b(new_n151), .c(new_n191), .out0(new_n281));
  norb02aa1n06x5               g186(.a(new_n274), .b(new_n275), .out0(new_n282));
  nano32aa1d12x5               g187(.a(new_n224), .b(new_n282), .c(new_n244), .d(new_n261), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n281), .c(new_n165), .d(new_n188), .o1(new_n284));
  nanp02aa1n02x5               g189(.a(\b[25] ), .b(\a[26] ), .o1(new_n285));
  oai022aa1n02x5               g190(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n286));
  aoi022aa1n12x5               g191(.a(new_n269), .b(new_n282), .c(new_n285), .d(new_n286), .o1(new_n287));
  xnrc02aa1n12x5               g192(.a(\b[26] ), .b(\a[27] ), .out0(new_n288));
  xobna2aa1n03x5               g193(.a(new_n288), .b(new_n284), .c(new_n287), .out0(\s[27] ));
  aobi12aa1n02x7               g194(.a(new_n283), .b(new_n189), .c(new_n194), .out0(new_n290));
  nanp02aa1n06x5               g195(.a(new_n269), .b(new_n282), .o1(new_n291));
  nanp02aa1n02x5               g196(.a(new_n286), .b(new_n285), .o1(new_n292));
  tech160nm_finand02aa1n05x5   g197(.a(new_n291), .b(new_n292), .o1(new_n293));
  and002aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o(new_n294));
  oabi12aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(new_n290), .out0(new_n295));
  nor042aa1n03x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  inv000aa1n03x5               g201(.a(new_n296), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n294), .c(new_n284), .d(new_n287), .o1(new_n298));
  tech160nm_fixorc02aa1n02p5x5 g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  norp02aa1n02x5               g204(.a(new_n299), .b(new_n296), .o1(new_n300));
  aoi022aa1n03x5               g205(.a(new_n298), .b(new_n299), .c(new_n295), .d(new_n300), .o1(\s[28] ));
  norb02aa1n06x4               g206(.a(new_n299), .b(new_n288), .out0(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n293), .c(new_n199), .d(new_n283), .o1(new_n303));
  inv000aa1n02x5               g208(.a(new_n302), .o1(new_n304));
  oao003aa1n03x5               g209(.a(\a[28] ), .b(\b[27] ), .c(new_n297), .carry(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n304), .c(new_n284), .d(new_n287), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g215(.a(new_n288), .b(new_n299), .c(new_n307), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n293), .c(new_n199), .d(new_n283), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  oaoi03aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .o1(new_n314));
  inv000aa1n03x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n284), .d(new_n287), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .out0(new_n317));
  and002aa1n02x5               g222(.a(\b[28] ), .b(\a[29] ), .o(new_n318));
  oabi12aa1n02x5               g223(.a(new_n317), .b(\a[29] ), .c(\b[28] ), .out0(new_n319));
  oab012aa1n02x4               g224(.a(new_n319), .b(new_n305), .c(new_n318), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n316), .b(new_n317), .c(new_n312), .d(new_n320), .o1(\s[30] ));
  nano32aa1d12x5               g226(.a(new_n288), .b(new_n317), .c(new_n299), .d(new_n307), .out0(new_n322));
  aoai13aa1n03x5               g227(.a(new_n322), .b(new_n293), .c(new_n199), .d(new_n283), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[31] ), .b(\b[30] ), .out0(new_n324));
  oao003aa1n02x5               g229(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n325));
  norb02aa1n02x5               g230(.a(new_n325), .b(new_n324), .out0(new_n326));
  inv000aa1n02x5               g231(.a(new_n322), .o1(new_n327));
  aoai13aa1n03x5               g232(.a(new_n325), .b(new_n327), .c(new_n284), .d(new_n287), .o1(new_n328));
  aoi022aa1n03x5               g233(.a(new_n328), .b(new_n324), .c(new_n323), .d(new_n326), .o1(\s[31] ));
  oai012aa1n02x5               g234(.a(new_n100), .b(new_n101), .c(new_n99), .o1(new_n330));
  xnrb03aa1n02x5               g235(.a(new_n330), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g236(.a(\a[3] ), .b(\b[2] ), .c(new_n330), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g238(.a(new_n105), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g239(.a(\a[5] ), .b(\b[4] ), .c(new_n159), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fioaoi03aa1n03p5x5 g241(.a(new_n114), .b(new_n115), .c(new_n335), .o1(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n337), .b(new_n118), .c(new_n109), .out0(\s[7] ));
  norb02aa1n02x5               g243(.a(new_n107), .b(new_n106), .out0(new_n339));
  nano22aa1n03x7               g244(.a(new_n337), .b(new_n118), .c(new_n109), .out0(new_n340));
  oabi12aa1n03x5               g245(.a(new_n339), .b(new_n340), .c(new_n108), .out0(new_n341));
  nano22aa1n02x4               g246(.a(new_n340), .b(new_n339), .c(new_n118), .out0(new_n342));
  nanb02aa1n03x5               g247(.a(new_n342), .b(new_n341), .out0(\s[8] ));
  xnbna2aa1n03x5               g248(.a(new_n122), .b(new_n197), .c(new_n164), .out0(\s[9] ));
endmodule


