// Benchmark "adder" written by ABC on Thu Jul 11 11:46:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n325, new_n327,
    new_n329, new_n330;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  xorc02aa1n02x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  and002aa1n02x5               g003(.a(\b[3] ), .b(\a[4] ), .o(new_n99));
  160nm_ficinv00aa1n08x5       g004(.clk(\a[3] ), .clkout(new_n100));
  160nm_ficinv00aa1n08x5       g005(.clk(\b[2] ), .clkout(new_n101));
  nanp02aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(new_n102), .b(new_n103), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  norp02aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  oai012aa1n02x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .o1(new_n108));
  160nm_ficinv00aa1n08x5       g013(.clk(\b[3] ), .clkout(new_n109));
  aboi22aa1n03x5               g014(.a(\a[4] ), .b(new_n109), .c(new_n100), .d(new_n101), .out0(new_n110));
  oaoi13aa1n02x5               g015(.a(new_n99), .b(new_n110), .c(new_n108), .d(new_n104), .o1(new_n111));
  norp02aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanb02aa1n02x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .out0(new_n115));
  norp02aa1n02x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  norp02aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nona23aa1n02x4               g024(.a(new_n119), .b(new_n117), .c(new_n116), .d(new_n118), .out0(new_n120));
  norp03aa1n02x5               g025(.a(new_n120), .b(new_n115), .c(new_n114), .o1(new_n121));
  aoi112aa1n02x5               g026(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n122));
  norb02aa1n02x5               g027(.a(new_n113), .b(new_n112), .out0(new_n123));
  xorc02aa1n02x5               g028(.a(\a[7] ), .b(\b[6] ), .out0(new_n124));
  aoi112aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  oai112aa1n02x5               g030(.a(new_n124), .b(new_n123), .c(new_n116), .d(new_n125), .o1(new_n126));
  nona22aa1n02x4               g031(.a(new_n126), .b(new_n122), .c(new_n112), .out0(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n111), .d(new_n121), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n97), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  norp02aa1n02x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  oai012aa1n02x5               g038(.a(new_n110), .b(new_n108), .c(new_n104), .o1(new_n134));
  oaib12aa1n02x5               g039(.a(new_n134), .b(new_n109), .c(\a[4] ), .out0(new_n135));
  norp02aa1n02x5               g040(.a(new_n115), .b(new_n114), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n120), .b(new_n136), .out0(new_n137));
  aoi012aa1n02x5               g042(.a(new_n116), .b(new_n118), .c(new_n117), .o1(new_n138));
  norp03aa1n02x5               g043(.a(new_n115), .b(new_n138), .c(new_n114), .o1(new_n139));
  norp03aa1n02x5               g044(.a(new_n139), .b(new_n122), .c(new_n112), .o1(new_n140));
  oai012aa1n02x5               g045(.a(new_n140), .b(new_n135), .c(new_n137), .o1(new_n141));
  and002aa1n02x5               g046(.a(new_n128), .b(new_n97), .o(new_n142));
  norp02aa1n02x5               g047(.a(\b[9] ), .b(\a[10] ), .o1(new_n143));
  aoi112aa1n02x5               g048(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n144));
  norp02aa1n02x5               g049(.a(new_n144), .b(new_n143), .o1(new_n145));
  aobi12aa1n02x5               g050(.a(new_n145), .b(new_n141), .c(new_n142), .out0(new_n146));
  xnrc02aa1n02x5               g051(.a(new_n146), .b(new_n133), .out0(\s[11] ));
  oaoi03aa1n02x5               g052(.a(\a[11] ), .b(\b[10] ), .c(new_n146), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norp02aa1n02x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nano23aa1n02x4               g056(.a(new_n131), .b(new_n150), .c(new_n151), .d(new_n132), .out0(new_n152));
  and003aa1n02x5               g057(.a(new_n152), .b(new_n128), .c(new_n97), .o(new_n153));
  aoai13aa1n02x5               g058(.a(new_n153), .b(new_n127), .c(new_n111), .d(new_n121), .o1(new_n154));
  aoi112aa1n02x5               g059(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n151), .b(new_n150), .out0(new_n156));
  oai112aa1n02x5               g061(.a(new_n156), .b(new_n133), .c(new_n144), .d(new_n143), .o1(new_n157));
  nona22aa1n02x4               g062(.a(new_n157), .b(new_n155), .c(new_n150), .out0(new_n158));
  160nm_ficinv00aa1n08x5       g063(.clk(new_n158), .clkout(new_n159));
  nanp02aa1n02x5               g064(.a(new_n154), .b(new_n159), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n162), .b(new_n160), .c(new_n163), .o1(new_n164));
  xnrb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n02x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nona23aa1n02x4               g072(.a(new_n167), .b(new_n163), .c(new_n162), .d(new_n166), .out0(new_n168));
  aoi012aa1n02x5               g073(.a(new_n166), .b(new_n162), .c(new_n167), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n168), .c(new_n154), .d(new_n159), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  160nm_ficinv00aa1n08x5       g079(.clk(new_n174), .clkout(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  aoi122aa1n02x5               g081(.a(new_n172), .b(new_n176), .c(new_n175), .d(new_n170), .e(new_n173), .o1(new_n177));
  aoi012aa1n02x5               g082(.a(new_n172), .b(new_n170), .c(new_n173), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n174), .b(new_n176), .out0(new_n179));
  norp02aa1n02x5               g084(.a(new_n178), .b(new_n179), .o1(new_n180));
  norp02aa1n02x5               g085(.a(new_n180), .b(new_n177), .o1(\s[16] ));
  nano23aa1n02x4               g086(.a(new_n162), .b(new_n166), .c(new_n167), .d(new_n163), .out0(new_n182));
  nano23aa1n02x4               g087(.a(new_n172), .b(new_n174), .c(new_n176), .d(new_n173), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n183), .b(new_n182), .o1(new_n184));
  nano32aa1n02x4               g089(.a(new_n184), .b(new_n152), .c(new_n128), .d(new_n97), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n127), .c(new_n111), .d(new_n121), .o1(new_n186));
  nanb02aa1n02x5               g091(.a(new_n172), .b(new_n173), .out0(new_n187));
  norp03aa1n02x5               g092(.a(new_n168), .b(new_n179), .c(new_n187), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n189));
  oai013aa1n02x4               g094(.a(new_n175), .b(new_n169), .c(new_n187), .d(new_n179), .o1(new_n190));
  aoi112aa1n02x5               g095(.a(new_n190), .b(new_n189), .c(new_n158), .d(new_n188), .o1(new_n191));
  norp02aa1n02x5               g096(.a(\b[16] ), .b(\a[17] ), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  norb02aa1n02x5               g098(.a(new_n193), .b(new_n192), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n191), .c(new_n186), .out0(\s[17] ));
  nanp03aa1n02x5               g100(.a(new_n191), .b(new_n186), .c(new_n194), .o1(new_n196));
  xnrc02aa1n02x5               g101(.a(\b[17] ), .b(\a[18] ), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n196), .c(new_n193), .out0(\s[18] ));
  norb02aa1n02x5               g103(.a(new_n194), .b(new_n197), .out0(new_n199));
  160nm_ficinv00aa1n08x5       g104(.clk(new_n199), .clkout(new_n200));
  160nm_ficinv00aa1n08x5       g105(.clk(\a[18] ), .clkout(new_n201));
  160nm_ficinv00aa1n08x5       g106(.clk(\b[17] ), .clkout(new_n202));
  oao003aa1n02x5               g107(.a(new_n201), .b(new_n202), .c(new_n192), .carry(new_n203));
  160nm_ficinv00aa1n08x5       g108(.clk(new_n203), .clkout(new_n204));
  aoai13aa1n02x5               g109(.a(new_n204), .b(new_n200), .c(new_n191), .d(new_n186), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nanp02aa1n02x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  norp02aa1n02x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nanp02aa1n02x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  norb02aa1n02x5               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  aoi112aa1n02x5               g117(.a(new_n208), .b(new_n212), .c(new_n205), .d(new_n209), .o1(new_n213));
  aoai13aa1n02x5               g118(.a(new_n212), .b(new_n208), .c(new_n205), .d(new_n209), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(\s[20] ));
  nano23aa1n02x4               g120(.a(new_n208), .b(new_n210), .c(new_n211), .d(new_n209), .out0(new_n216));
  nanb03aa1n02x5               g121(.a(new_n197), .b(new_n216), .c(new_n194), .out0(new_n217));
  aoi112aa1n02x5               g122(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n218));
  aoi112aa1n02x5               g123(.a(new_n218), .b(new_n210), .c(new_n216), .d(new_n203), .o1(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n217), .c(new_n191), .d(new_n186), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  xnrc02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .out0(new_n223));
  160nm_ficinv00aa1n08x5       g128(.clk(new_n223), .clkout(new_n224));
  xnrc02aa1n02x5               g129(.a(\b[21] ), .b(\a[22] ), .out0(new_n225));
  160nm_ficinv00aa1n08x5       g130(.clk(new_n225), .clkout(new_n226));
  aoi112aa1n02x5               g131(.a(new_n222), .b(new_n226), .c(new_n220), .d(new_n224), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n226), .b(new_n222), .c(new_n220), .d(new_n224), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(\s[22] ));
  norp02aa1n02x5               g134(.a(new_n225), .b(new_n223), .o1(new_n230));
  nanp03aa1n02x5               g135(.a(new_n199), .b(new_n230), .c(new_n216), .o1(new_n231));
  norp02aa1n02x5               g136(.a(\b[17] ), .b(\a[18] ), .o1(new_n232));
  aoi112aa1n02x5               g137(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n209), .b(new_n208), .out0(new_n234));
  oai112aa1n02x5               g139(.a(new_n234), .b(new_n212), .c(new_n233), .d(new_n232), .o1(new_n235));
  nona22aa1n02x4               g140(.a(new_n235), .b(new_n218), .c(new_n210), .out0(new_n236));
  160nm_ficinv00aa1n08x5       g141(.clk(new_n222), .clkout(new_n237));
  oaoi03aa1n02x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(new_n236), .c(new_n230), .o1(new_n239));
  aoai13aa1n02x5               g144(.a(new_n239), .b(new_n231), .c(new_n191), .d(new_n186), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  nanp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  norp02aa1n02x5               g148(.a(\b[23] ), .b(\a[24] ), .o1(new_n244));
  nanp02aa1n02x5               g149(.a(\b[23] ), .b(\a[24] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  aoi112aa1n02x5               g151(.a(new_n242), .b(new_n246), .c(new_n240), .d(new_n243), .o1(new_n247));
  aoai13aa1n02x5               g152(.a(new_n246), .b(new_n242), .c(new_n240), .d(new_n243), .o1(new_n248));
  norb02aa1n02x5               g153(.a(new_n248), .b(new_n247), .out0(\s[24] ));
  nona23aa1n02x4               g154(.a(new_n245), .b(new_n243), .c(new_n242), .d(new_n244), .out0(new_n250));
  160nm_ficinv00aa1n08x5       g155(.clk(new_n250), .clkout(new_n251));
  nanb03aa1n02x5               g156(.a(new_n217), .b(new_n251), .c(new_n230), .out0(new_n252));
  nona32aa1n02x4               g157(.a(new_n236), .b(new_n250), .c(new_n225), .d(new_n223), .out0(new_n253));
  aoi112aa1n02x5               g158(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n254), .b(new_n244), .c(new_n251), .d(new_n238), .o1(new_n255));
  nanp02aa1n02x5               g160(.a(new_n253), .b(new_n255), .o1(new_n256));
  160nm_ficinv00aa1n08x5       g161(.clk(new_n256), .clkout(new_n257));
  aoai13aa1n02x5               g162(.a(new_n257), .b(new_n252), .c(new_n191), .d(new_n186), .o1(new_n258));
  xorb03aa1n02x5               g163(.a(new_n258), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g164(.a(\b[24] ), .b(\a[25] ), .o1(new_n260));
  xorc02aa1n02x5               g165(.a(\a[25] ), .b(\b[24] ), .out0(new_n261));
  xorc02aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .out0(new_n262));
  aoi112aa1n02x5               g167(.a(new_n260), .b(new_n262), .c(new_n258), .d(new_n261), .o1(new_n263));
  aoai13aa1n02x5               g168(.a(new_n262), .b(new_n260), .c(new_n258), .d(new_n261), .o1(new_n264));
  norb02aa1n02x5               g169(.a(new_n264), .b(new_n263), .out0(\s[26] ));
  nanp02aa1n02x5               g170(.a(new_n158), .b(new_n188), .o1(new_n266));
  nona22aa1n02x4               g171(.a(new_n266), .b(new_n190), .c(new_n189), .out0(new_n267));
  nano32aa1n02x4               g172(.a(new_n231), .b(new_n262), .c(new_n251), .d(new_n261), .out0(new_n268));
  aoai13aa1n02x5               g173(.a(new_n268), .b(new_n267), .c(new_n141), .d(new_n185), .o1(new_n269));
  nanp02aa1n02x5               g174(.a(\b[25] ), .b(\a[26] ), .o1(new_n270));
  and002aa1n02x5               g175(.a(new_n262), .b(new_n261), .o(new_n271));
  oai022aa1n02x5               g176(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n272));
  aoi022aa1n02x5               g177(.a(new_n256), .b(new_n271), .c(new_n270), .d(new_n272), .o1(new_n273));
  norp02aa1n02x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(\b[26] ), .b(\a[27] ), .o1(new_n275));
  norb02aa1n02x5               g180(.a(new_n275), .b(new_n274), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n269), .c(new_n273), .out0(\s[27] ));
  xorc02aa1n02x5               g182(.a(\a[28] ), .b(\b[27] ), .out0(new_n278));
  nanp02aa1n02x5               g183(.a(new_n191), .b(new_n186), .o1(new_n279));
  160nm_ficinv00aa1n08x5       g184(.clk(new_n271), .clkout(new_n280));
  nanp02aa1n02x5               g185(.a(new_n272), .b(new_n270), .o1(new_n281));
  aoai13aa1n02x5               g186(.a(new_n281), .b(new_n280), .c(new_n253), .d(new_n255), .o1(new_n282));
  aoi112aa1n02x5               g187(.a(new_n274), .b(new_n282), .c(new_n279), .d(new_n268), .o1(new_n283));
  nano22aa1n02x4               g188(.a(new_n283), .b(new_n275), .c(new_n278), .out0(new_n284));
  160nm_ficinv00aa1n08x5       g189(.clk(\a[28] ), .clkout(new_n285));
  160nm_ficinv00aa1n08x5       g190(.clk(\b[27] ), .clkout(new_n286));
  nanp02aa1n02x5               g191(.a(new_n286), .b(new_n285), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(\b[27] ), .b(\a[28] ), .o1(new_n288));
  160nm_ficinv00aa1n08x5       g193(.clk(new_n274), .clkout(new_n289));
  nanp03aa1n02x5               g194(.a(new_n269), .b(new_n273), .c(new_n289), .o1(new_n290));
  aoi022aa1n02x5               g195(.a(new_n290), .b(new_n275), .c(new_n287), .d(new_n288), .o1(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n284), .o1(\s[28] ));
  nano32aa1n02x4               g197(.a(new_n274), .b(new_n288), .c(new_n275), .d(new_n287), .out0(new_n293));
  aoai13aa1n02x5               g198(.a(new_n293), .b(new_n282), .c(new_n279), .d(new_n268), .o1(new_n294));
  oaoi03aa1n02x5               g199(.a(new_n285), .b(new_n286), .c(new_n274), .o1(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[28] ), .b(\a[29] ), .out0(new_n296));
  aoi012aa1n02x5               g201(.a(new_n296), .b(new_n294), .c(new_n295), .o1(new_n297));
  160nm_ficinv00aa1n08x5       g202(.clk(new_n293), .clkout(new_n298));
  aoi012aa1n02x5               g203(.a(new_n298), .b(new_n269), .c(new_n273), .o1(new_n299));
  nano22aa1n02x4               g204(.a(new_n299), .b(new_n295), .c(new_n296), .out0(new_n300));
  norp02aa1n02x5               g205(.a(new_n297), .b(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g206(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g207(.a(new_n296), .b(new_n276), .c(new_n287), .d(new_n288), .out0(new_n303));
  aoai13aa1n02x5               g208(.a(new_n303), .b(new_n282), .c(new_n279), .d(new_n268), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .carry(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .out0(new_n306));
  aoi012aa1n02x5               g211(.a(new_n306), .b(new_n304), .c(new_n305), .o1(new_n307));
  160nm_ficinv00aa1n08x5       g212(.clk(new_n303), .clkout(new_n308));
  aoi012aa1n02x5               g213(.a(new_n308), .b(new_n269), .c(new_n273), .o1(new_n309));
  nano22aa1n02x4               g214(.a(new_n309), .b(new_n305), .c(new_n306), .out0(new_n310));
  norp02aa1n02x5               g215(.a(new_n307), .b(new_n310), .o1(\s[30] ));
  nano23aa1n02x4               g216(.a(new_n306), .b(new_n296), .c(new_n278), .d(new_n276), .out0(new_n312));
  160nm_ficinv00aa1n08x5       g217(.clk(new_n312), .clkout(new_n313));
  aoi012aa1n02x5               g218(.a(new_n313), .b(new_n269), .c(new_n273), .o1(new_n314));
  oao003aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  nano22aa1n02x4               g221(.a(new_n314), .b(new_n315), .c(new_n316), .out0(new_n317));
  aoai13aa1n02x5               g222(.a(new_n312), .b(new_n282), .c(new_n279), .d(new_n268), .o1(new_n318));
  aoi012aa1n02x5               g223(.a(new_n316), .b(new_n318), .c(new_n315), .o1(new_n319));
  norp02aa1n02x5               g224(.a(new_n319), .b(new_n317), .o1(\s[31] ));
  xnbna2aa1n03x5               g225(.a(new_n108), .b(new_n102), .c(new_n103), .out0(\s[3] ));
  oaoi03aa1n02x5               g226(.a(\a[3] ), .b(\b[2] ), .c(new_n108), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g228(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g229(.a(new_n118), .b(new_n111), .c(new_n119), .o1(new_n325));
  xnrb03aa1n02x5               g230(.a(new_n325), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nona22aa1n02x4               g231(.a(new_n134), .b(new_n120), .c(new_n99), .out0(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n124), .b(new_n327), .c(new_n138), .out0(\s[7] ));
  orn002aa1n02x5               g233(.a(\a[7] ), .b(\b[6] ), .o(new_n329));
  aob012aa1n02x5               g234(.a(new_n124), .b(new_n327), .c(new_n138), .out0(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n123), .b(new_n330), .c(new_n329), .out0(\s[8] ));
  xorb03aa1n02x5               g236(.a(new_n141), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


