// Benchmark "adder" written by ABC on Wed Jul 17 12:52:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n325, new_n326,
    new_n328, new_n330;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  nor042aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  and002aa1n02x5               g003(.a(\b[8] ), .b(\a[9] ), .o(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  inv040aa1d32x5               g005(.a(\a[2] ), .o1(new_n101));
  inv040aa1d32x5               g006(.a(\b[1] ), .o1(new_n102));
  nand22aa1n06x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  oao003aa1n02x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .carry(new_n104));
  nor002aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nand42aa1d28x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nor022aa1n16x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1d28x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nano23aa1n02x5               g013(.a(new_n105), .b(new_n107), .c(new_n108), .d(new_n106), .out0(new_n109));
  oaih12aa1n02x5               g014(.a(new_n106), .b(new_n107), .c(new_n105), .o1(new_n110));
  aobi12aa1n06x5               g015(.a(new_n110), .b(new_n109), .c(new_n104), .out0(new_n111));
  xnrc02aa1n12x5               g016(.a(\b[5] ), .b(\a[6] ), .out0(new_n112));
  nor022aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand42aa1n06x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor002aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nano23aa1n03x7               g021(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n117));
  tech160nm_fixnrc02aa1n03p5x5 g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  nona22aa1n09x5               g023(.a(new_n117), .b(new_n118), .c(new_n112), .out0(new_n119));
  oaih12aa1n02x5               g024(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n120));
  orn002aa1n24x5               g025(.a(\a[5] ), .b(\b[4] ), .o(new_n121));
  oaoi03aa1n12x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n121), .o1(new_n122));
  aobi12aa1n06x5               g027(.a(new_n120), .b(new_n117), .c(new_n122), .out0(new_n123));
  oai012aa1n06x5               g028(.a(new_n123), .b(new_n111), .c(new_n119), .o1(new_n124));
  aoai13aa1n02x5               g029(.a(new_n97), .b(new_n98), .c(new_n124), .d(new_n100), .o1(new_n125));
  tech160nm_fioaoi03aa1n02p5x5 g030(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n126));
  nona23aa1n02x4               g031(.a(new_n108), .b(new_n106), .c(new_n105), .d(new_n107), .out0(new_n127));
  oaih12aa1n02x5               g032(.a(new_n110), .b(new_n127), .c(new_n126), .o1(new_n128));
  nona23aa1n03x5               g033(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n129));
  nor043aa1n02x5               g034(.a(new_n129), .b(new_n118), .c(new_n112), .o1(new_n130));
  oaib12aa1n03x5               g035(.a(new_n120), .b(new_n129), .c(new_n122), .out0(new_n131));
  aoai13aa1n03x5               g036(.a(new_n100), .b(new_n131), .c(new_n128), .d(new_n130), .o1(new_n132));
  nona22aa1n03x5               g037(.a(new_n132), .b(new_n98), .c(new_n97), .out0(new_n133));
  nanp02aa1n02x5               g038(.a(new_n125), .b(new_n133), .o1(\s[10] ));
  inv000aa1d42x5               g039(.a(\a[10] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(\b[9] ), .o1(new_n136));
  norp02aa1n12x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  tech160nm_finand02aa1n03p5x5 g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  oai112aa1n03x5               g044(.a(new_n133), .b(new_n139), .c(new_n136), .d(new_n135), .o1(new_n140));
  oaoi13aa1n02x5               g045(.a(new_n139), .b(new_n133), .c(new_n135), .d(new_n136), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(\s[11] ));
  inv000aa1n02x5               g047(.a(new_n137), .o1(new_n143));
  nor022aa1n16x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n03x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n140), .c(new_n143), .out0(\s[12] ));
  nona23aa1n09x5               g052(.a(new_n145), .b(new_n138), .c(new_n137), .d(new_n144), .out0(new_n148));
  oaoi03aa1n02x5               g053(.a(new_n135), .b(new_n136), .c(new_n98), .o1(new_n149));
  oaoi03aa1n03x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n143), .o1(new_n150));
  oabi12aa1n03x5               g055(.a(new_n150), .b(new_n148), .c(new_n149), .out0(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[8] ), .b(\a[9] ), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  norp02aa1n02x5               g058(.a(new_n148), .b(new_n97), .o1(new_n154));
  aoi013aa1n03x5               g059(.a(new_n151), .b(new_n124), .c(new_n153), .d(new_n154), .o1(new_n155));
  nor002aa1d32x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  nand22aa1n06x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n155), .b(new_n158), .c(new_n157), .out0(\s[13] ));
  oaoi03aa1n03x5               g064(.a(\a[13] ), .b(\b[12] ), .c(new_n155), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n16x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand02aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nona23aa1n09x5               g068(.a(new_n163), .b(new_n158), .c(new_n156), .d(new_n162), .out0(new_n164));
  nona23aa1n03x5               g069(.a(new_n124), .b(new_n154), .c(new_n164), .d(new_n152), .out0(new_n165));
  inv040aa1n02x5               g070(.a(new_n164), .o1(new_n166));
  aoi012aa1n12x5               g071(.a(new_n162), .b(new_n156), .c(new_n163), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n168), .b(new_n151), .c(new_n166), .o1(new_n169));
  nor002aa1d32x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand22aa1n12x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n165), .c(new_n169), .out0(\s[15] ));
  inv000aa1d42x5               g078(.a(new_n170), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n172), .o1(new_n175));
  aoai13aa1n03x5               g080(.a(new_n174), .b(new_n175), .c(new_n165), .d(new_n169), .o1(new_n176));
  xorb03aa1n02x5               g081(.a(new_n176), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  aoi012aa1n06x5               g082(.a(new_n131), .b(new_n128), .c(new_n130), .o1(new_n178));
  nor002aa1n06x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand02aa1n04x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nona23aa1n09x5               g085(.a(new_n180), .b(new_n171), .c(new_n170), .d(new_n179), .out0(new_n181));
  nor042aa1n02x5               g086(.a(new_n181), .b(new_n164), .o1(new_n182));
  nona32aa1n09x5               g087(.a(new_n182), .b(new_n148), .c(new_n152), .d(new_n97), .out0(new_n183));
  nano23aa1n02x4               g088(.a(new_n170), .b(new_n179), .c(new_n180), .d(new_n171), .out0(new_n184));
  aoai13aa1n04x5               g089(.a(new_n184), .b(new_n168), .c(new_n151), .d(new_n166), .o1(new_n185));
  aoi012aa1n02x7               g090(.a(new_n179), .b(new_n170), .c(new_n180), .o1(new_n186));
  oai112aa1n04x5               g091(.a(new_n185), .b(new_n186), .c(new_n178), .d(new_n183), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[16] ), .o1(new_n191));
  oaoi03aa1n03x5               g096(.a(new_n190), .b(new_n191), .c(new_n187), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(new_n189), .out0(\s[18] ));
  oaoi13aa1n12x5               g098(.a(new_n183), .b(new_n123), .c(new_n111), .d(new_n119), .o1(new_n194));
  nano23aa1n03x5               g099(.a(new_n137), .b(new_n144), .c(new_n145), .d(new_n138), .out0(new_n195));
  oao003aa1n03x5               g100(.a(new_n135), .b(new_n136), .c(new_n98), .carry(new_n196));
  aoai13aa1n04x5               g101(.a(new_n166), .b(new_n150), .c(new_n195), .d(new_n196), .o1(new_n197));
  aoai13aa1n09x5               g102(.a(new_n186), .b(new_n181), .c(new_n197), .d(new_n167), .o1(new_n198));
  xroi22aa1d06x4               g103(.a(new_n190), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n199));
  tech160nm_fioai012aa1n03p5x5 g104(.a(new_n199), .b(new_n198), .c(new_n194), .o1(new_n200));
  oaih22aa1n04x5               g105(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n201));
  oaib12aa1n09x5               g106(.a(new_n201), .b(new_n189), .c(\b[17] ), .out0(new_n202));
  nor042aa1n12x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand22aa1n12x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n203), .b(new_n204), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n200), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g113(.a(new_n203), .o1(new_n209));
  tech160nm_fiaoi012aa1n02p5x5 g114(.a(new_n205), .b(new_n200), .c(new_n202), .o1(new_n210));
  nor042aa1n04x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nand22aa1n12x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nanb02aa1n02x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  nano22aa1n03x5               g118(.a(new_n210), .b(new_n209), .c(new_n213), .out0(new_n214));
  nanp02aa1n02x5               g119(.a(new_n191), .b(new_n190), .o1(new_n215));
  oaoi03aa1n02x5               g120(.a(\a[18] ), .b(\b[17] ), .c(new_n215), .o1(new_n216));
  oaoi13aa1n03x5               g121(.a(new_n216), .b(new_n199), .c(new_n198), .d(new_n194), .o1(new_n217));
  oaoi13aa1n02x7               g122(.a(new_n213), .b(new_n209), .c(new_n217), .d(new_n205), .o1(new_n218));
  norp02aa1n03x5               g123(.a(new_n218), .b(new_n214), .o1(\s[20] ));
  nano23aa1n06x5               g124(.a(new_n203), .b(new_n211), .c(new_n212), .d(new_n204), .out0(new_n220));
  nand02aa1n03x5               g125(.a(new_n199), .b(new_n220), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  tech160nm_fioai012aa1n03p5x5 g127(.a(new_n222), .b(new_n198), .c(new_n194), .o1(new_n223));
  nona23aa1d18x5               g128(.a(new_n212), .b(new_n204), .c(new_n203), .d(new_n211), .out0(new_n224));
  aoi012aa1n09x5               g129(.a(new_n211), .b(new_n203), .c(new_n212), .o1(new_n225));
  oai012aa1d24x5               g130(.a(new_n225), .b(new_n224), .c(new_n202), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  nor042aa1n09x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  xnbna2aa1n03x5               g135(.a(new_n230), .b(new_n223), .c(new_n227), .out0(\s[21] ));
  inv000aa1d42x5               g136(.a(new_n228), .o1(new_n232));
  aobi12aa1n02x7               g137(.a(new_n230), .b(new_n223), .c(new_n227), .out0(new_n233));
  tech160nm_fixnrc02aa1n02p5x5 g138(.a(\b[21] ), .b(\a[22] ), .out0(new_n234));
  nano22aa1n03x5               g139(.a(new_n233), .b(new_n232), .c(new_n234), .out0(new_n235));
  aoai13aa1n03x5               g140(.a(new_n230), .b(new_n226), .c(new_n187), .d(new_n222), .o1(new_n236));
  tech160nm_fiaoi012aa1n02p5x5 g141(.a(new_n234), .b(new_n236), .c(new_n232), .o1(new_n237));
  norp02aa1n03x5               g142(.a(new_n237), .b(new_n235), .o1(\s[22] ));
  nano22aa1n03x7               g143(.a(new_n234), .b(new_n232), .c(new_n229), .out0(new_n239));
  and003aa1n02x5               g144(.a(new_n199), .b(new_n239), .c(new_n220), .o(new_n240));
  tech160nm_fioai012aa1n03p5x5 g145(.a(new_n240), .b(new_n198), .c(new_n194), .o1(new_n241));
  oao003aa1n12x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n232), .carry(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n243), .b(new_n226), .c(new_n239), .o1(new_n244));
  xnrc02aa1n12x5               g149(.a(\b[22] ), .b(\a[23] ), .out0(new_n245));
  inv000aa1d42x5               g150(.a(new_n245), .o1(new_n246));
  xnbna2aa1n03x5               g151(.a(new_n246), .b(new_n241), .c(new_n244), .out0(\s[23] ));
  nor042aa1n03x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  tech160nm_fiaoi012aa1n02p5x5 g154(.a(new_n245), .b(new_n241), .c(new_n244), .o1(new_n250));
  xnrc02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .out0(new_n251));
  nano22aa1n02x4               g156(.a(new_n250), .b(new_n249), .c(new_n251), .out0(new_n252));
  inv000aa1n03x5               g157(.a(new_n244), .o1(new_n253));
  oaoi13aa1n03x5               g158(.a(new_n253), .b(new_n240), .c(new_n198), .d(new_n194), .o1(new_n254));
  oaoi13aa1n02x7               g159(.a(new_n251), .b(new_n249), .c(new_n254), .d(new_n245), .o1(new_n255));
  norp02aa1n03x5               g160(.a(new_n255), .b(new_n252), .o1(\s[24] ));
  nor042aa1n02x5               g161(.a(new_n251), .b(new_n245), .o1(new_n257));
  nano22aa1n03x7               g162(.a(new_n221), .b(new_n239), .c(new_n257), .out0(new_n258));
  oaih12aa1n02x5               g163(.a(new_n258), .b(new_n198), .c(new_n194), .o1(new_n259));
  inv040aa1n03x5               g164(.a(new_n225), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n239), .b(new_n260), .c(new_n220), .d(new_n216), .o1(new_n261));
  inv000aa1n02x5               g166(.a(new_n257), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .carry(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n261), .d(new_n242), .o1(new_n264));
  xnrc02aa1n12x5               g169(.a(\b[24] ), .b(\a[25] ), .out0(new_n265));
  aoib12aa1n06x5               g170(.a(new_n265), .b(new_n259), .c(new_n264), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n265), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n267), .b(new_n264), .c(new_n187), .d(new_n258), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n266), .b(new_n268), .o1(\s[25] ));
  nor042aa1n03x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  tech160nm_fixnrc02aa1n04x5   g176(.a(\b[25] ), .b(\a[26] ), .out0(new_n272));
  nano22aa1n03x5               g177(.a(new_n266), .b(new_n271), .c(new_n272), .out0(new_n273));
  oaoi13aa1n03x5               g178(.a(new_n264), .b(new_n258), .c(new_n198), .d(new_n194), .o1(new_n274));
  oaoi13aa1n02x7               g179(.a(new_n272), .b(new_n271), .c(new_n274), .d(new_n265), .o1(new_n275));
  norp02aa1n03x5               g180(.a(new_n275), .b(new_n273), .o1(\s[26] ));
  nor042aa1n03x5               g181(.a(new_n272), .b(new_n265), .o1(new_n277));
  nano32aa1n03x7               g182(.a(new_n221), .b(new_n277), .c(new_n239), .d(new_n257), .out0(new_n278));
  oai012aa1n06x5               g183(.a(new_n278), .b(new_n198), .c(new_n194), .o1(new_n279));
  oao003aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .carry(new_n280));
  aobi12aa1n06x5               g185(.a(new_n280), .b(new_n264), .c(new_n277), .out0(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n279), .c(new_n281), .out0(\s[27] ));
  norp02aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  inv040aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  aobi12aa1n02x7               g190(.a(new_n282), .b(new_n279), .c(new_n281), .out0(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[27] ), .b(\a[28] ), .out0(new_n287));
  nano22aa1n03x5               g192(.a(new_n286), .b(new_n285), .c(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n257), .b(new_n243), .c(new_n226), .d(new_n239), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n277), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n280), .b(new_n290), .c(new_n289), .d(new_n263), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n282), .b(new_n291), .c(new_n187), .d(new_n278), .o1(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n287), .b(new_n292), .c(new_n285), .o1(new_n293));
  norp02aa1n03x5               g198(.a(new_n293), .b(new_n288), .o1(\s[28] ));
  norb02aa1n02x5               g199(.a(new_n282), .b(new_n287), .out0(new_n295));
  aobi12aa1n02x7               g200(.a(new_n295), .b(new_n279), .c(new_n281), .out0(new_n296));
  oao003aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[28] ), .b(\a[29] ), .out0(new_n298));
  nano22aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  aoai13aa1n02x5               g204(.a(new_n295), .b(new_n291), .c(new_n187), .d(new_n278), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  norp02aa1n03x5               g206(.a(new_n301), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g208(.a(new_n282), .b(new_n298), .c(new_n287), .out0(new_n304));
  aobi12aa1n02x7               g209(.a(new_n304), .b(new_n279), .c(new_n281), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[29] ), .b(\a[30] ), .out0(new_n307));
  nano22aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n307), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n304), .b(new_n291), .c(new_n187), .d(new_n278), .o1(new_n309));
  tech160nm_fiaoi012aa1n02p5x5 g214(.a(new_n307), .b(new_n309), .c(new_n306), .o1(new_n310));
  norp02aa1n03x5               g215(.a(new_n310), .b(new_n308), .o1(\s[30] ));
  norb02aa1n02x5               g216(.a(new_n304), .b(new_n307), .out0(new_n312));
  aobi12aa1n02x7               g217(.a(new_n312), .b(new_n279), .c(new_n281), .out0(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  nano22aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n315), .out0(new_n316));
  aoai13aa1n02x5               g221(.a(new_n312), .b(new_n291), .c(new_n187), .d(new_n278), .o1(new_n317));
  tech160nm_fiaoi012aa1n02p5x5 g222(.a(new_n315), .b(new_n317), .c(new_n314), .o1(new_n318));
  norp02aa1n03x5               g223(.a(new_n318), .b(new_n316), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n126), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n126), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n128), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g228(.a(new_n112), .o1(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n324), .b(new_n121), .c(new_n111), .d(new_n118), .o1(new_n325));
  oai112aa1n02x5               g230(.a(new_n121), .b(new_n324), .c(new_n111), .d(new_n118), .o1(new_n326));
  nanb02aa1n02x5               g231(.a(new_n325), .b(new_n326), .out0(\s[6] ));
  aob012aa1n02x5               g232(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g234(.a(\a[7] ), .b(\b[6] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrc02aa1n02x5               g236(.a(new_n178), .b(new_n153), .out0(\s[9] ));
endmodule


