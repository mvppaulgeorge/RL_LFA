// Benchmark "adder" written by ABC on Thu Jul 18 12:51:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n192, new_n193,
    new_n194, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n342, new_n343, new_n344,
    new_n345, new_n347, new_n349, new_n351, new_n352, new_n354, new_n355,
    new_n357, new_n358, new_n360;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n20x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv040aa1d32x5               g003(.a(\a[4] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[3] ), .o1(new_n100));
  nor042aa1n06x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  tech160nm_fioaoi03aa1n03p5x5 g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(new_n100), .b(new_n99), .o1(new_n103));
  nor042aa1n09x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand22aa1n12x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  oai112aa1n06x5               g011(.a(new_n103), .b(new_n105), .c(new_n104), .d(new_n106), .o1(new_n107));
  nanp02aa1n04x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand42aa1n04x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanb03aa1n09x5               g014(.a(new_n101), .b(new_n109), .c(new_n108), .out0(new_n110));
  oai012aa1n18x5               g015(.a(new_n102), .b(new_n107), .c(new_n110), .o1(new_n111));
  nor042aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand02aa1d10x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  norb02aa1n06x4               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  nor042aa1n06x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n06x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  norb02aa1n06x4               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nor042aa1n06x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nanp02aa1n06x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  nor002aa1d32x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nand02aa1n06x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nona23aa1n09x5               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  nano22aa1n12x5               g027(.a(new_n122), .b(new_n114), .c(new_n117), .out0(new_n123));
  nanb02aa1n12x5               g028(.a(new_n118), .b(new_n119), .out0(new_n124));
  nanb03aa1d24x5               g029(.a(new_n120), .b(new_n121), .c(new_n113), .out0(new_n125));
  nor042aa1n04x5               g030(.a(new_n115), .b(new_n112), .o1(new_n126));
  tech160nm_fioai012aa1n03p5x5 g031(.a(new_n119), .b(new_n120), .c(new_n118), .o1(new_n127));
  oai013aa1d12x5               g032(.a(new_n127), .b(new_n125), .c(new_n124), .d(new_n126), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  aoai13aa1n03x5               g034(.a(new_n129), .b(new_n128), .c(new_n111), .d(new_n123), .o1(new_n130));
  nor002aa1n20x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nand02aa1d28x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  norb02aa1d27x5               g037(.a(new_n132), .b(new_n131), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n133), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  aob012aa1n03x5               g039(.a(new_n133), .b(new_n130), .c(new_n98), .out0(new_n135));
  oai022aa1n09x5               g040(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n136));
  aob012aa1n02x5               g041(.a(new_n135), .b(new_n136), .c(new_n132), .out0(new_n137));
  nor022aa1n16x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nand02aa1n06x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aboi22aa1n03x5               g045(.a(new_n138), .b(new_n139), .c(new_n136), .d(new_n132), .out0(new_n141));
  aoi022aa1n02x5               g046(.a(new_n137), .b(new_n140), .c(new_n135), .d(new_n141), .o1(\s[11] ));
  nor002aa1n16x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand22aa1n09x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  aoai13aa1n02x5               g050(.a(new_n145), .b(new_n138), .c(new_n137), .d(new_n139), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n133), .o1(new_n147));
  aoi012aa1n02x5               g052(.a(new_n147), .b(new_n130), .c(new_n98), .o1(new_n148));
  aoai13aa1n02x5               g053(.a(new_n140), .b(new_n148), .c(new_n132), .d(new_n136), .o1(new_n149));
  nona22aa1n02x4               g054(.a(new_n149), .b(new_n145), .c(new_n138), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n146), .b(new_n150), .o1(\s[12] ));
  nand22aa1n06x5               g056(.a(new_n111), .b(new_n123), .o1(new_n152));
  norp03aa1n06x5               g057(.a(new_n125), .b(new_n124), .c(new_n126), .o1(new_n153));
  norb02aa1n09x5               g058(.a(new_n127), .b(new_n153), .out0(new_n154));
  nona23aa1d18x5               g059(.a(new_n144), .b(new_n139), .c(new_n138), .d(new_n143), .out0(new_n155));
  nano22aa1d15x5               g060(.a(new_n155), .b(new_n129), .c(new_n133), .out0(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n157), .b(new_n152), .c(new_n154), .o1(new_n158));
  aoi012aa1d24x5               g063(.a(new_n128), .b(new_n111), .c(new_n123), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nanb03aa1n02x5               g065(.a(new_n143), .b(new_n144), .c(new_n139), .out0(new_n161));
  oai112aa1n02x5               g066(.a(new_n136), .b(new_n132), .c(\b[10] ), .d(\a[11] ), .o1(new_n162));
  aoi012aa1n06x5               g067(.a(new_n143), .b(new_n138), .c(new_n144), .o1(new_n163));
  tech160nm_fioai012aa1n03p5x5 g068(.a(new_n163), .b(new_n162), .c(new_n161), .o1(new_n164));
  nor002aa1d32x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand02aa1n04x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n164), .c(new_n160), .d(new_n156), .o1(new_n169));
  oai112aa1n02x5               g074(.a(new_n163), .b(new_n167), .c(new_n162), .d(new_n161), .o1(new_n170));
  oa0012aa1n02x5               g075(.a(new_n169), .b(new_n170), .c(new_n158), .o(\s[13] ));
  oaoi13aa1n03x5               g076(.a(new_n165), .b(new_n166), .c(new_n158), .d(new_n164), .o1(new_n172));
  xnrb03aa1n02x5               g077(.a(new_n172), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nand02aa1n08x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nona23aa1d18x5               g080(.a(new_n175), .b(new_n166), .c(new_n165), .d(new_n174), .out0(new_n176));
  nona22aa1n02x4               g081(.a(new_n160), .b(new_n157), .c(new_n176), .out0(new_n177));
  inv040aa1n09x5               g082(.a(new_n176), .o1(new_n178));
  nona23aa1n02x4               g083(.a(new_n178), .b(new_n129), .c(new_n155), .d(new_n147), .out0(new_n179));
  nano22aa1n03x7               g084(.a(new_n143), .b(new_n139), .c(new_n144), .out0(new_n180));
  oai012aa1n02x5               g085(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .o1(new_n181));
  oab012aa1n04x5               g086(.a(new_n181), .b(new_n97), .c(new_n131), .out0(new_n182));
  inv000aa1n06x5               g087(.a(new_n163), .o1(new_n183));
  aoai13aa1n12x5               g088(.a(new_n178), .b(new_n183), .c(new_n182), .d(new_n180), .o1(new_n184));
  oai012aa1d24x5               g089(.a(new_n175), .b(new_n174), .c(new_n165), .o1(new_n185));
  oai112aa1n04x5               g090(.a(new_n184), .b(new_n185), .c(new_n159), .d(new_n179), .o1(new_n186));
  xnrc02aa1n12x5               g091(.a(\b[14] ), .b(\a[15] ), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(new_n185), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(new_n188), .b(new_n189), .c(new_n164), .d(new_n178), .o1(new_n190));
  aoi022aa1n02x5               g095(.a(new_n186), .b(new_n188), .c(new_n177), .d(new_n190), .o1(\s[15] ));
  inv000aa1d42x5               g096(.a(\a[16] ), .o1(new_n192));
  nor042aa1n04x5               g097(.a(\b[14] ), .b(\a[15] ), .o1(new_n193));
  tech160nm_fiaoi012aa1n05x5   g098(.a(new_n193), .b(new_n186), .c(new_n188), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[15] ), .c(new_n192), .out0(\s[16] ));
  tech160nm_fixnrc02aa1n04x5   g100(.a(\b[15] ), .b(\a[16] ), .out0(new_n196));
  nona32aa1d24x5               g101(.a(new_n156), .b(new_n196), .c(new_n187), .d(new_n176), .out0(new_n197));
  aoi012aa1d24x5               g102(.a(new_n197), .b(new_n152), .c(new_n154), .o1(new_n198));
  norp02aa1n04x5               g103(.a(new_n196), .b(new_n187), .o1(new_n199));
  aoai13aa1n04x5               g104(.a(new_n199), .b(new_n189), .c(new_n164), .d(new_n178), .o1(new_n200));
  inv000aa1d42x5               g105(.a(\b[15] ), .o1(new_n201));
  oao003aa1n02x5               g106(.a(new_n192), .b(new_n201), .c(new_n193), .carry(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  oai112aa1n06x5               g108(.a(new_n200), .b(new_n203), .c(new_n159), .d(new_n197), .o1(new_n204));
  xorc02aa1n12x5               g109(.a(\a[17] ), .b(\b[16] ), .out0(new_n205));
  nano22aa1n02x4               g110(.a(new_n205), .b(new_n200), .c(new_n203), .out0(new_n206));
  aboi22aa1n03x5               g111(.a(new_n198), .b(new_n206), .c(new_n204), .d(new_n205), .out0(\s[17] ));
  inv000aa1d42x5               g112(.a(\a[18] ), .o1(new_n208));
  inv000aa1n03x5               g113(.a(new_n199), .o1(new_n209));
  aoai13aa1n12x5               g114(.a(new_n203), .b(new_n209), .c(new_n184), .d(new_n185), .o1(new_n210));
  norp02aa1n24x5               g115(.a(\b[16] ), .b(\a[17] ), .o1(new_n211));
  oaoi13aa1n06x5               g116(.a(new_n211), .b(new_n205), .c(new_n210), .d(new_n198), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[17] ), .c(new_n208), .out0(\s[18] ));
  nor002aa1d32x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  nand02aa1d24x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  nano22aa1n12x5               g120(.a(new_n214), .b(new_n205), .c(new_n215), .out0(new_n216));
  oai012aa1n06x5               g121(.a(new_n216), .b(new_n210), .c(new_n198), .o1(new_n217));
  oa0012aa1n02x5               g122(.a(new_n215), .b(new_n214), .c(new_n211), .o(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  nor042aa1d18x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nand02aa1n06x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n06x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n217), .c(new_n219), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand02aa1d04x5               g129(.a(new_n217), .b(new_n219), .o1(new_n225));
  nor002aa1n16x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  nand02aa1d24x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nanb02aa1n02x5               g132(.a(new_n226), .b(new_n227), .out0(new_n228));
  aoai13aa1n03x5               g133(.a(new_n228), .b(new_n220), .c(new_n225), .d(new_n221), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n222), .b(new_n218), .c(new_n204), .d(new_n216), .o1(new_n230));
  nona22aa1n03x5               g135(.a(new_n230), .b(new_n228), .c(new_n220), .out0(new_n231));
  nanp02aa1n03x5               g136(.a(new_n229), .b(new_n231), .o1(\s[20] ));
  nanb03aa1d18x5               g137(.a(new_n228), .b(new_n216), .c(new_n222), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  oai012aa1n06x5               g139(.a(new_n234), .b(new_n210), .c(new_n198), .o1(new_n235));
  nanb03aa1n06x5               g140(.a(new_n226), .b(new_n227), .c(new_n221), .out0(new_n236));
  oai122aa1n06x5               g141(.a(new_n215), .b(new_n214), .c(new_n211), .d(\b[18] ), .e(\a[19] ), .o1(new_n237));
  aoi012aa1n12x5               g142(.a(new_n226), .b(new_n220), .c(new_n227), .o1(new_n238));
  oai012aa1n12x5               g143(.a(new_n238), .b(new_n237), .c(new_n236), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nanp02aa1n03x5               g145(.a(new_n235), .b(new_n240), .o1(new_n241));
  nor042aa1d18x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  nand42aa1n10x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n243), .b(new_n242), .out0(new_n244));
  nano22aa1n03x7               g149(.a(new_n226), .b(new_n221), .c(new_n227), .out0(new_n245));
  oai012aa1n04x7               g150(.a(new_n215), .b(\b[18] ), .c(\a[19] ), .o1(new_n246));
  oab012aa1n06x5               g151(.a(new_n246), .b(new_n211), .c(new_n214), .out0(new_n247));
  inv020aa1n03x5               g152(.a(new_n238), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n248), .b(new_n244), .c(new_n247), .d(new_n245), .o1(new_n249));
  aoi022aa1n02x5               g154(.a(new_n241), .b(new_n244), .c(new_n235), .d(new_n249), .o1(\s[21] ));
  nor042aa1d18x5               g155(.a(\b[21] ), .b(\a[22] ), .o1(new_n251));
  nand42aa1n10x5               g156(.a(\b[21] ), .b(\a[22] ), .o1(new_n252));
  nanb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n242), .c(new_n241), .d(new_n244), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n244), .b(new_n239), .c(new_n204), .d(new_n234), .o1(new_n255));
  nona22aa1n03x5               g160(.a(new_n255), .b(new_n253), .c(new_n242), .out0(new_n256));
  nanp02aa1n03x5               g161(.a(new_n254), .b(new_n256), .o1(\s[22] ));
  nano23aa1d15x5               g162(.a(new_n242), .b(new_n251), .c(new_n252), .d(new_n243), .out0(new_n258));
  nano32aa1n02x4               g163(.a(new_n228), .b(new_n216), .c(new_n258), .d(new_n222), .out0(new_n259));
  oai012aa1n06x5               g164(.a(new_n259), .b(new_n210), .c(new_n198), .o1(new_n260));
  oa0012aa1n06x5               g165(.a(new_n252), .b(new_n251), .c(new_n242), .o(new_n261));
  aoi012aa1n02x5               g166(.a(new_n261), .b(new_n239), .c(new_n258), .o1(new_n262));
  nanp02aa1n03x5               g167(.a(new_n260), .b(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  aoi112aa1n02x5               g169(.a(new_n264), .b(new_n261), .c(new_n239), .d(new_n258), .o1(new_n265));
  aoi022aa1n02x5               g170(.a(new_n263), .b(new_n264), .c(new_n260), .d(new_n265), .o1(\s[23] ));
  norp02aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .o1(new_n267));
  tech160nm_fixnrc02aa1n05x5   g172(.a(\b[23] ), .b(\a[24] ), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n263), .d(new_n264), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n262), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n264), .b(new_n270), .c(new_n204), .d(new_n259), .o1(new_n271));
  nona22aa1n02x4               g176(.a(new_n271), .b(new_n268), .c(new_n267), .out0(new_n272));
  nanp02aa1n03x5               g177(.a(new_n269), .b(new_n272), .o1(\s[24] ));
  norb02aa1n06x4               g178(.a(new_n264), .b(new_n268), .out0(new_n274));
  nano22aa1n03x7               g179(.a(new_n233), .b(new_n258), .c(new_n274), .out0(new_n275));
  oai012aa1n06x5               g180(.a(new_n275), .b(new_n210), .c(new_n198), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n258), .b(new_n248), .c(new_n247), .d(new_n245), .o1(new_n277));
  inv040aa1n02x5               g182(.a(new_n261), .o1(new_n278));
  inv040aa1n02x5               g183(.a(new_n274), .o1(new_n279));
  oai022aa1n02x5               g184(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n280));
  aob012aa1n02x5               g185(.a(new_n280), .b(\b[23] ), .c(\a[24] ), .out0(new_n281));
  aoai13aa1n12x5               g186(.a(new_n281), .b(new_n279), .c(new_n277), .d(new_n278), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n282), .o1(new_n283));
  nanp02aa1n06x5               g188(.a(new_n276), .b(new_n283), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  aoai13aa1n03x5               g190(.a(new_n274), .b(new_n261), .c(new_n239), .d(new_n258), .o1(new_n286));
  nano22aa1n02x4               g191(.a(new_n285), .b(new_n286), .c(new_n281), .out0(new_n287));
  aoi022aa1n02x5               g192(.a(new_n284), .b(new_n285), .c(new_n276), .d(new_n287), .o1(\s[25] ));
  norp02aa1n02x5               g193(.a(\b[24] ), .b(\a[25] ), .o1(new_n289));
  tech160nm_fixnrc02aa1n04x5   g194(.a(\b[25] ), .b(\a[26] ), .out0(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n289), .c(new_n284), .d(new_n285), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n285), .b(new_n282), .c(new_n204), .d(new_n275), .o1(new_n292));
  nona22aa1n03x5               g197(.a(new_n292), .b(new_n290), .c(new_n289), .out0(new_n293));
  nanp02aa1n03x5               g198(.a(new_n291), .b(new_n293), .o1(\s[26] ));
  norb02aa1n06x5               g199(.a(new_n285), .b(new_n290), .out0(new_n295));
  nano32aa1n03x7               g200(.a(new_n233), .b(new_n295), .c(new_n258), .d(new_n274), .out0(new_n296));
  oai012aa1n18x5               g201(.a(new_n296), .b(new_n210), .c(new_n198), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(\b[25] ), .b(\a[26] ), .o1(new_n298));
  oai022aa1n02x5               g203(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n299));
  aoi022aa1d18x5               g204(.a(new_n282), .b(new_n295), .c(new_n298), .d(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  xnbna2aa1n03x5               g206(.a(new_n301), .b(new_n297), .c(new_n300), .out0(\s[27] ));
  xnrc02aa1n02x5               g207(.a(\b[27] ), .b(\a[28] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  inv000aa1n03x5               g209(.a(new_n304), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n301), .o1(new_n306));
  aoai13aa1n06x5               g211(.a(new_n305), .b(new_n306), .c(new_n297), .d(new_n300), .o1(new_n307));
  nanp02aa1n03x5               g212(.a(new_n307), .b(new_n303), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n295), .o1(new_n309));
  nanp02aa1n02x5               g214(.a(new_n299), .b(new_n298), .o1(new_n310));
  aoai13aa1n02x7               g215(.a(new_n310), .b(new_n309), .c(new_n286), .d(new_n281), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n301), .b(new_n311), .c(new_n204), .d(new_n296), .o1(new_n312));
  nona22aa1n02x4               g217(.a(new_n312), .b(new_n303), .c(new_n304), .out0(new_n313));
  nanp02aa1n03x5               g218(.a(new_n308), .b(new_n313), .o1(\s[28] ));
  norb02aa1n02x5               g219(.a(new_n301), .b(new_n303), .out0(new_n315));
  aoai13aa1n02x5               g220(.a(new_n315), .b(new_n311), .c(new_n204), .d(new_n296), .o1(new_n316));
  tech160nm_fixorc02aa1n03p5x5 g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  oao003aa1n02x5               g222(.a(\a[28] ), .b(\b[27] ), .c(new_n305), .carry(new_n318));
  norb02aa1n02x5               g223(.a(new_n318), .b(new_n317), .out0(new_n319));
  inv000aa1n02x5               g224(.a(new_n315), .o1(new_n320));
  aoai13aa1n06x5               g225(.a(new_n318), .b(new_n320), .c(new_n297), .d(new_n300), .o1(new_n321));
  aoi022aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n316), .d(new_n319), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nand02aa1n03x5               g228(.a(new_n297), .b(new_n300), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n317), .o1(new_n325));
  nona32aa1n03x5               g230(.a(new_n324), .b(new_n325), .c(new_n303), .d(new_n306), .out0(new_n326));
  xorc02aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .out0(new_n327));
  oaoi03aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .c(new_n318), .o1(new_n328));
  norp02aa1n02x5               g233(.a(new_n328), .b(new_n327), .o1(new_n329));
  nanb03aa1n02x5               g234(.a(new_n303), .b(new_n317), .c(new_n301), .out0(new_n330));
  inv000aa1n03x5               g235(.a(new_n328), .o1(new_n331));
  aoai13aa1n06x5               g236(.a(new_n331), .b(new_n330), .c(new_n297), .d(new_n300), .o1(new_n332));
  aoi022aa1n02x7               g237(.a(new_n326), .b(new_n329), .c(new_n332), .d(new_n327), .o1(\s[30] ));
  inv000aa1n02x5               g238(.a(new_n327), .o1(new_n334));
  nona32aa1n03x5               g239(.a(new_n324), .b(new_n334), .c(new_n325), .d(new_n320), .out0(new_n335));
  xorc02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  oao003aa1n02x5               g241(.a(\a[30] ), .b(\b[29] ), .c(new_n331), .carry(new_n337));
  norb02aa1n02x5               g242(.a(new_n337), .b(new_n336), .out0(new_n338));
  nona22aa1n02x4               g243(.a(new_n315), .b(new_n325), .c(new_n334), .out0(new_n339));
  aoai13aa1n06x5               g244(.a(new_n337), .b(new_n339), .c(new_n297), .d(new_n300), .o1(new_n340));
  aoi022aa1n02x7               g245(.a(new_n335), .b(new_n338), .c(new_n340), .d(new_n336), .o1(\s[31] ));
  norb03aa1n02x5               g246(.a(new_n105), .b(new_n104), .c(new_n106), .out0(new_n342));
  oai012aa1n02x5               g247(.a(new_n105), .b(new_n104), .c(new_n106), .o1(new_n343));
  nanb03aa1n02x5               g248(.a(new_n101), .b(new_n343), .c(new_n109), .out0(new_n344));
  oaib12aa1n02x5               g249(.a(new_n105), .b(new_n101), .c(new_n109), .out0(new_n345));
  oai012aa1n02x5               g250(.a(new_n344), .b(new_n345), .c(new_n342), .o1(\s[3] ));
  nanp02aa1n02x5               g251(.a(new_n103), .b(new_n108), .o1(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n347), .b(new_n344), .c(new_n109), .out0(\s[4] ));
  orn002aa1n02x5               g253(.a(new_n107), .b(new_n110), .o(new_n349));
  xnbna2aa1n03x5               g254(.a(new_n117), .b(new_n349), .c(new_n102), .out0(\s[5] ));
  aoai13aa1n02x5               g255(.a(new_n114), .b(new_n115), .c(new_n111), .d(new_n116), .o1(new_n351));
  aoi112aa1n02x5               g256(.a(new_n115), .b(new_n114), .c(new_n111), .d(new_n117), .o1(new_n352));
  norb02aa1n02x5               g257(.a(new_n351), .b(new_n352), .out0(\s[6] ));
  nanb02aa1n02x5               g258(.a(new_n120), .b(new_n121), .out0(new_n354));
  oai012aa1n02x5               g259(.a(new_n113), .b(new_n115), .c(new_n112), .o1(new_n355));
  xobna2aa1n03x5               g260(.a(new_n354), .b(new_n351), .c(new_n355), .out0(\s[7] ));
  inv000aa1d42x5               g261(.a(new_n120), .o1(new_n357));
  aoai13aa1n02x5               g262(.a(new_n357), .b(new_n354), .c(new_n351), .d(new_n355), .o1(new_n358));
  xorb03aa1n02x5               g263(.a(new_n358), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  norb03aa1n02x5               g264(.a(new_n127), .b(new_n153), .c(new_n129), .out0(new_n360));
  aboi22aa1n03x5               g265(.a(new_n159), .b(new_n129), .c(new_n360), .d(new_n152), .out0(\s[9] ));
endmodule


