// Benchmark "adder" written by ABC on Wed Jul 17 21:41:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n310,
    new_n312, new_n314, new_n316, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n03x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n06x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  inv000aa1d42x5               g004(.a(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[8] ), .o1(new_n101));
  norp02aa1n06x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nand42aa1d28x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nor042aa1n09x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nanp02aa1n09x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nano23aa1n03x5               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  nanp02aa1n04x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor022aa1n16x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  oa0012aa1n03x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o(new_n110));
  oa0012aa1n02x5               g015(.a(new_n103), .b(new_n104), .c(new_n102), .o(new_n111));
  aoi012aa1n06x5               g016(.a(new_n111), .b(new_n106), .c(new_n110), .o1(new_n112));
  nor042aa1d18x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  inv030aa1n02x5               g018(.a(new_n113), .o1(new_n114));
  oao003aa1n06x5               g019(.a(\a[4] ), .b(\b[3] ), .c(new_n114), .carry(new_n115));
  tech160nm_fixorc02aa1n02p5x5 g020(.a(\a[4] ), .b(\b[3] ), .out0(new_n116));
  nand42aa1n16x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  norb02aa1n02x7               g022(.a(new_n117), .b(new_n113), .out0(new_n118));
  and002aa1n12x5               g023(.a(\b[1] ), .b(\a[2] ), .o(new_n119));
  nand22aa1n12x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  norp02aa1n06x5               g025(.a(\b[1] ), .b(\a[2] ), .o1(new_n121));
  oab012aa1n09x5               g026(.a(new_n119), .b(new_n121), .c(new_n120), .out0(new_n122));
  nand43aa1n06x5               g027(.a(new_n122), .b(new_n116), .c(new_n118), .o1(new_n123));
  nand02aa1n03x5               g028(.a(\b[4] ), .b(\a[5] ), .o1(new_n124));
  nano23aa1n02x5               g029(.a(new_n109), .b(new_n108), .c(new_n124), .d(new_n107), .out0(new_n125));
  nand02aa1n02x5               g030(.a(new_n125), .b(new_n106), .o1(new_n126));
  aoai13aa1n12x5               g031(.a(new_n112), .b(new_n126), .c(new_n123), .d(new_n115), .o1(new_n127));
  oaoi03aa1n09x5               g032(.a(new_n100), .b(new_n101), .c(new_n127), .o1(new_n128));
  xnrc02aa1n02x5               g033(.a(new_n128), .b(new_n99), .out0(\s[10] ));
  tech160nm_fioaoi03aa1n03p5x5 g034(.a(\a[10] ), .b(\b[9] ), .c(new_n128), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n20x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1n10x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  tech160nm_finand02aa1n05x5   g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  aoai13aa1n02x5               g041(.a(new_n136), .b(new_n132), .c(new_n130), .d(new_n133), .o1(new_n137));
  nanp02aa1n02x5               g042(.a(new_n128), .b(new_n99), .o1(new_n138));
  nanb02aa1n12x5               g043(.a(new_n132), .b(new_n133), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nand03aa1n02x5               g045(.a(new_n138), .b(new_n98), .c(new_n140), .o1(new_n141));
  nona22aa1n02x4               g046(.a(new_n141), .b(new_n136), .c(new_n132), .out0(new_n142));
  nanp02aa1n03x5               g047(.a(new_n137), .b(new_n142), .o1(\s[12] ));
  aoai13aa1n06x5               g048(.a(new_n98), .b(new_n97), .c(new_n100), .d(new_n101), .o1(new_n144));
  oa0012aa1n02x5               g049(.a(new_n135), .b(new_n134), .c(new_n132), .o(new_n145));
  inv000aa1n02x5               g050(.a(new_n145), .o1(new_n146));
  oai013aa1n03x5               g051(.a(new_n146), .b(new_n144), .c(new_n139), .d(new_n136), .o1(new_n147));
  nano23aa1n06x5               g052(.a(new_n132), .b(new_n134), .c(new_n135), .d(new_n133), .out0(new_n148));
  tech160nm_fixorc02aa1n03p5x5 g053(.a(\a[9] ), .b(\b[8] ), .out0(new_n149));
  nanp03aa1d12x5               g054(.a(new_n148), .b(new_n99), .c(new_n149), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[12] ), .b(\a[13] ), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n02x5               g058(.a(new_n153), .b(new_n147), .c(new_n127), .d(new_n151), .o1(new_n154));
  aoi112aa1n02x5               g059(.a(new_n147), .b(new_n153), .c(new_n127), .d(new_n151), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n154), .b(new_n155), .out0(\s[13] ));
  nor042aa1n03x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  inv000aa1n03x5               g062(.a(new_n157), .o1(new_n158));
  tech160nm_fixnrc02aa1n04x5   g063(.a(\b[13] ), .b(\a[14] ), .out0(new_n159));
  xobna2aa1n03x5               g064(.a(new_n159), .b(new_n154), .c(new_n158), .out0(\s[14] ));
  nor042aa1n09x5               g065(.a(new_n159), .b(new_n152), .o1(new_n161));
  oaoi03aa1n03x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n158), .o1(new_n162));
  aoi012aa1n06x5               g067(.a(new_n162), .b(new_n147), .c(new_n161), .o1(new_n163));
  nona32aa1n03x5               g068(.a(new_n127), .b(new_n159), .c(new_n152), .d(new_n150), .out0(new_n164));
  xnrc02aa1n12x5               g069(.a(\b[14] ), .b(\a[15] ), .out0(new_n165));
  xobna2aa1n03x5               g070(.a(new_n165), .b(new_n164), .c(new_n163), .out0(\s[15] ));
  nor042aa1n06x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n03x5               g073(.a(new_n168), .b(new_n165), .c(new_n164), .d(new_n163), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  inv040aa1d32x5               g075(.a(\a[17] ), .o1(new_n171));
  tech160nm_fixnrc02aa1n02p5x5 g076(.a(\b[15] ), .b(\a[16] ), .out0(new_n172));
  nor002aa1n03x5               g077(.a(new_n172), .b(new_n165), .o1(new_n173));
  nano22aa1n06x5               g078(.a(new_n150), .b(new_n161), .c(new_n173), .out0(new_n174));
  oaoi03aa1n12x5               g079(.a(\a[16] ), .b(\b[15] ), .c(new_n168), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n101), .b(new_n100), .o1(new_n176));
  oaoi03aa1n02x5               g081(.a(\a[10] ), .b(\b[9] ), .c(new_n176), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n161), .b(new_n145), .c(new_n148), .d(new_n177), .o1(new_n178));
  inv000aa1n02x5               g083(.a(new_n162), .o1(new_n179));
  inv000aa1n02x5               g084(.a(new_n173), .o1(new_n180));
  aoi012aa1n03x5               g085(.a(new_n180), .b(new_n178), .c(new_n179), .o1(new_n181));
  aoi112aa1n09x5               g086(.a(new_n181), .b(new_n175), .c(new_n127), .d(new_n174), .o1(new_n182));
  xorb03aa1n02x5               g087(.a(new_n182), .b(\b[16] ), .c(new_n171), .out0(\s[17] ));
  oaoi03aa1n03x5               g088(.a(\a[17] ), .b(\b[16] ), .c(new_n182), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g090(.a(\a[18] ), .o1(new_n186));
  xroi22aa1d06x4               g091(.a(new_n171), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n187));
  inv000aa1n02x5               g092(.a(new_n187), .o1(new_n188));
  oai022aa1n04x7               g093(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n189));
  oaib12aa1n06x5               g094(.a(new_n189), .b(new_n186), .c(\b[17] ), .out0(new_n190));
  tech160nm_fioai012aa1n05x5   g095(.a(new_n190), .b(new_n182), .c(new_n188), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g097(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand42aa1n04x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nanb02aa1n02x5               g100(.a(new_n194), .b(new_n195), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  nor042aa1n09x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nanp02aa1n12x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  aoai13aa1n03x5               g105(.a(new_n200), .b(new_n194), .c(new_n191), .d(new_n197), .o1(new_n201));
  nanp02aa1n06x5               g106(.a(new_n127), .b(new_n174), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n175), .o1(new_n203));
  oai112aa1n06x5               g108(.a(new_n202), .b(new_n203), .c(new_n163), .d(new_n180), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(\b[16] ), .b(new_n171), .out0(new_n205));
  oaoi03aa1n12x5               g110(.a(\a[18] ), .b(\b[17] ), .c(new_n205), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n197), .b(new_n206), .c(new_n204), .d(new_n187), .o1(new_n207));
  nona22aa1n02x4               g112(.a(new_n207), .b(new_n200), .c(new_n194), .out0(new_n208));
  nanp02aa1n03x5               g113(.a(new_n201), .b(new_n208), .o1(\s[20] ));
  nona23aa1d18x5               g114(.a(new_n199), .b(new_n195), .c(new_n194), .d(new_n198), .out0(new_n210));
  oa0012aa1n03x5               g115(.a(new_n199), .b(new_n198), .c(new_n194), .o(new_n211));
  inv040aa1n03x5               g116(.a(new_n211), .o1(new_n212));
  oai012aa1d24x5               g117(.a(new_n212), .b(new_n210), .c(new_n190), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  nano23aa1n09x5               g119(.a(new_n194), .b(new_n198), .c(new_n199), .d(new_n195), .out0(new_n215));
  nand22aa1n09x5               g120(.a(new_n187), .b(new_n215), .o1(new_n216));
  tech160nm_fioai012aa1n05x5   g121(.a(new_n214), .b(new_n182), .c(new_n216), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xnrc02aa1n12x5               g124(.a(\b[20] ), .b(\a[21] ), .out0(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  tech160nm_fixnrc02aa1n05x5   g126(.a(\b[21] ), .b(\a[22] ), .out0(new_n222));
  aoai13aa1n03x5               g127(.a(new_n222), .b(new_n219), .c(new_n217), .d(new_n221), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n216), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n221), .b(new_n213), .c(new_n204), .d(new_n224), .o1(new_n225));
  nona22aa1n02x4               g130(.a(new_n225), .b(new_n222), .c(new_n219), .out0(new_n226));
  nanp02aa1n03x5               g131(.a(new_n223), .b(new_n226), .o1(\s[22] ));
  nor042aa1n06x5               g132(.a(new_n222), .b(new_n220), .o1(new_n228));
  inv040aa1d32x5               g133(.a(\a[22] ), .o1(new_n229));
  inv040aa1d32x5               g134(.a(\b[21] ), .o1(new_n230));
  oao003aa1n09x5               g135(.a(new_n229), .b(new_n230), .c(new_n219), .carry(new_n231));
  aoi012aa1d24x5               g136(.a(new_n231), .b(new_n213), .c(new_n228), .o1(new_n232));
  nano22aa1n06x5               g137(.a(new_n188), .b(new_n228), .c(new_n215), .out0(new_n233));
  inv000aa1n02x5               g138(.a(new_n233), .o1(new_n234));
  tech160nm_fioai012aa1n05x5   g139(.a(new_n232), .b(new_n182), .c(new_n234), .o1(new_n235));
  xorb03aa1n02x5               g140(.a(new_n235), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g141(.a(\b[22] ), .b(\a[23] ), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  tech160nm_fixnrc02aa1n05x5   g143(.a(\b[23] ), .b(\a[24] ), .out0(new_n239));
  aoai13aa1n03x5               g144(.a(new_n239), .b(new_n237), .c(new_n235), .d(new_n238), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n232), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n238), .b(new_n241), .c(new_n204), .d(new_n233), .o1(new_n242));
  nona22aa1n02x4               g147(.a(new_n242), .b(new_n239), .c(new_n237), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n240), .b(new_n243), .o1(\s[24] ));
  norb02aa1n02x5               g149(.a(new_n238), .b(new_n239), .out0(new_n245));
  inv030aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  nano32aa1n02x4               g151(.a(new_n246), .b(new_n187), .c(new_n228), .d(new_n215), .out0(new_n247));
  inv020aa1n02x5               g152(.a(new_n247), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n228), .b(new_n211), .c(new_n215), .d(new_n206), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n231), .o1(new_n250));
  oai022aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n251));
  aob012aa1n02x5               g156(.a(new_n251), .b(\b[23] ), .c(\a[24] ), .out0(new_n252));
  aoai13aa1n04x5               g157(.a(new_n252), .b(new_n246), .c(new_n249), .d(new_n250), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  tech160nm_fioai012aa1n05x5   g159(.a(new_n254), .b(new_n182), .c(new_n248), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[25] ), .b(\a[26] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n258), .b(new_n253), .c(new_n204), .d(new_n247), .o1(new_n261));
  nona22aa1n02x4               g166(.a(new_n261), .b(new_n259), .c(new_n257), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n260), .b(new_n262), .o1(\s[26] ));
  nanp02aa1n02x5               g168(.a(\b[25] ), .b(\a[26] ), .o1(new_n264));
  norb02aa1n12x5               g169(.a(new_n258), .b(new_n259), .out0(new_n265));
  oai022aa1n02x5               g170(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n266));
  aoi022aa1n09x5               g171(.a(new_n253), .b(new_n265), .c(new_n264), .d(new_n266), .o1(new_n267));
  nano23aa1n06x5               g172(.a(new_n216), .b(new_n246), .c(new_n265), .d(new_n228), .out0(new_n268));
  inv020aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  oai012aa1n12x5               g174(.a(new_n267), .b(new_n182), .c(new_n269), .o1(new_n270));
  xorb03aa1n02x5               g175(.a(new_n270), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  xorc02aa1n02x5               g177(.a(\a[27] ), .b(\b[26] ), .out0(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[27] ), .b(\a[28] ), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .d(new_n273), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n245), .b(new_n231), .c(new_n213), .d(new_n228), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n265), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(new_n266), .b(new_n264), .o1(new_n278));
  aoai13aa1n04x5               g183(.a(new_n278), .b(new_n277), .c(new_n276), .d(new_n252), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n273), .b(new_n279), .c(new_n204), .d(new_n268), .o1(new_n280));
  nona22aa1n02x5               g185(.a(new_n280), .b(new_n274), .c(new_n272), .out0(new_n281));
  nanp02aa1n03x5               g186(.a(new_n275), .b(new_n281), .o1(\s[28] ));
  norb02aa1n02x5               g187(.a(new_n273), .b(new_n274), .out0(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n279), .c(new_n204), .d(new_n268), .o1(new_n284));
  inv000aa1n03x5               g189(.a(new_n272), .o1(new_n285));
  oaoi03aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .o1(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[28] ), .b(\a[29] ), .out0(new_n287));
  nona22aa1n02x4               g192(.a(new_n284), .b(new_n286), .c(new_n287), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n287), .b(new_n286), .c(new_n270), .d(new_n283), .o1(new_n289));
  nanp02aa1n03x5               g194(.a(new_n289), .b(new_n288), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g196(.a(new_n273), .b(new_n287), .c(new_n274), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[28] ), .b(\b[27] ), .c(new_n285), .carry(new_n293));
  oaoi03aa1n02x5               g198(.a(\a[29] ), .b(\b[28] ), .c(new_n293), .o1(new_n294));
  tech160nm_fixorc02aa1n03p5x5 g199(.a(\a[30] ), .b(\b[29] ), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n294), .c(new_n270), .d(new_n292), .o1(new_n297));
  aoai13aa1n02x5               g202(.a(new_n292), .b(new_n279), .c(new_n204), .d(new_n268), .o1(new_n298));
  nona22aa1n02x4               g203(.a(new_n298), .b(new_n294), .c(new_n296), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[30] ));
  nanp02aa1n02x5               g205(.a(new_n294), .b(new_n295), .o1(new_n301));
  oai012aa1n02x5               g206(.a(new_n301), .b(\b[29] ), .c(\a[30] ), .o1(new_n302));
  nano23aa1n03x5               g207(.a(new_n287), .b(new_n274), .c(new_n295), .d(new_n273), .out0(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n279), .c(new_n204), .d(new_n268), .o1(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[30] ), .b(\a[31] ), .out0(new_n305));
  nona22aa1n02x5               g210(.a(new_n304), .b(new_n305), .c(new_n302), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n305), .b(new_n302), .c(new_n270), .d(new_n303), .o1(new_n307));
  nanp02aa1n03x5               g212(.a(new_n307), .b(new_n306), .o1(\s[31] ));
  xobna2aa1n03x5               g213(.a(new_n122), .b(new_n117), .c(new_n114), .out0(\s[3] ));
  oai012aa1n02x5               g214(.a(new_n117), .b(new_n122), .c(new_n113), .o1(new_n310));
  xnrb03aa1n02x5               g215(.a(new_n310), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  nanp02aa1n02x5               g216(.a(new_n123), .b(new_n115), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g218(.a(new_n109), .b(new_n312), .c(new_n124), .o1(new_n314));
  xnrb03aa1n02x5               g219(.a(new_n314), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g220(.a(new_n110), .b(new_n312), .c(new_n125), .o(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g222(.a(new_n104), .b(new_n316), .c(new_n105), .o1(new_n318));
  xnrb03aa1n02x5               g223(.a(new_n318), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g224(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


