// Benchmark "adder" written by ABC on Thu Jul 18 08:04:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n334, new_n337, new_n339, new_n340, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  norb02aa1n06x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  xorc02aa1n12x5               g004(.a(\a[7] ), .b(\b[6] ), .out0(new_n100));
  nor002aa1n04x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  nand22aa1n04x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  nor002aa1n02x5               g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[4] ), .b(\a[5] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  nano22aa1n03x7               g010(.a(new_n105), .b(new_n100), .c(new_n99), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\a[2] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[1] ), .o1(new_n108));
  nand22aa1n02x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  tech160nm_fioaoi03aa1n03p5x5 g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  nor022aa1n06x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[2] ), .b(\a[3] ), .o1(new_n114));
  nona23aa1n02x4               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  oa0012aa1n02x5               g020(.a(new_n112), .b(new_n113), .c(new_n111), .o(new_n116));
  oabi12aa1n12x5               g021(.a(new_n116), .b(new_n110), .c(new_n115), .out0(new_n117));
  aoi112aa1n02x5               g022(.a(\b[6] ), .b(\a[7] ), .c(\a[8] ), .d(\b[7] ), .o1(new_n118));
  aoi112aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n119));
  oai112aa1n02x7               g024(.a(new_n100), .b(new_n99), .c(new_n101), .d(new_n119), .o1(new_n120));
  nona22aa1n03x5               g025(.a(new_n120), .b(new_n118), .c(new_n97), .out0(new_n121));
  tech160nm_fiaoi012aa1n04x5   g026(.a(new_n121), .b(new_n117), .c(new_n106), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[9] ), .b(\b[8] ), .c(new_n122), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1d18x5               g029(.a(\b[10] ), .b(\a[11] ), .o1(new_n125));
  nand42aa1d28x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  norb02aa1n06x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  nanb03aa1n02x5               g032(.a(new_n105), .b(new_n99), .c(new_n100), .out0(new_n128));
  oao003aa1n02x5               g033(.a(new_n107), .b(new_n108), .c(new_n109), .carry(new_n129));
  nano23aa1n02x4               g034(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n130));
  aoi012aa1n02x5               g035(.a(new_n116), .b(new_n130), .c(new_n129), .o1(new_n131));
  tech160nm_fiao0012aa1n02p5x5 g036(.a(new_n101), .b(new_n103), .c(new_n102), .o(new_n132));
  aoi113aa1n02x5               g037(.a(new_n118), .b(new_n97), .c(new_n132), .d(new_n100), .e(new_n98), .o1(new_n133));
  tech160nm_fioai012aa1n03p5x5 g038(.a(new_n133), .b(new_n128), .c(new_n131), .o1(new_n134));
  xorc02aa1n12x5               g039(.a(\a[9] ), .b(\b[8] ), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  xorc02aa1n12x5               g041(.a(\a[10] ), .b(\b[9] ), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  nona22aa1n02x4               g043(.a(new_n134), .b(new_n136), .c(new_n138), .out0(new_n139));
  inv000aa1d42x5               g044(.a(\a[10] ), .o1(new_n140));
  inv000aa1d42x5               g045(.a(\b[9] ), .o1(new_n141));
  norp02aa1n02x5               g046(.a(\b[8] ), .b(\a[9] ), .o1(new_n142));
  oao003aa1n02x5               g047(.a(new_n140), .b(new_n141), .c(new_n142), .carry(new_n143));
  inv000aa1d42x5               g048(.a(new_n143), .o1(new_n144));
  xnbna2aa1n03x5               g049(.a(new_n127), .b(new_n139), .c(new_n144), .out0(\s[11] ));
  aobi12aa1n02x5               g050(.a(new_n127), .b(new_n139), .c(new_n144), .out0(new_n146));
  nor002aa1n16x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand42aa1n16x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n06x4               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  norp03aa1n02x5               g054(.a(new_n146), .b(new_n149), .c(new_n125), .o1(new_n150));
  oai012aa1n02x5               g055(.a(new_n149), .b(new_n146), .c(new_n125), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(\s[12] ));
  aoi112aa1n02x7               g057(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n153));
  nor002aa1n02x5               g058(.a(\b[9] ), .b(\a[10] ), .o1(new_n154));
  aoi112aa1n09x5               g059(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n155));
  oai112aa1n06x5               g060(.a(new_n149), .b(new_n127), .c(new_n155), .d(new_n154), .o1(new_n156));
  nona22aa1d24x5               g061(.a(new_n156), .b(new_n153), .c(new_n147), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  nano23aa1d15x5               g063(.a(new_n125), .b(new_n147), .c(new_n148), .d(new_n126), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  nona32aa1n02x4               g065(.a(new_n134), .b(new_n160), .c(new_n138), .d(new_n136), .out0(new_n161));
  nor042aa1n06x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand02aa1n08x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  xobna2aa1n03x5               g069(.a(new_n164), .b(new_n161), .c(new_n158), .out0(\s[13] ));
  nanp02aa1n02x5               g070(.a(new_n161), .b(new_n158), .o1(new_n166));
  nor042aa1n04x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nand02aa1n10x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nanb02aa1n12x5               g073(.a(new_n167), .b(new_n168), .out0(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n162), .b(new_n170), .c(new_n166), .d(new_n163), .o1(new_n171));
  aoai13aa1n02x5               g076(.a(new_n170), .b(new_n162), .c(new_n166), .d(new_n163), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(\s[14] ));
  nano23aa1d18x5               g078(.a(new_n162), .b(new_n167), .c(new_n168), .d(new_n163), .out0(new_n174));
  tech160nm_fiaoi012aa1n04x5   g079(.a(new_n167), .b(new_n162), .c(new_n168), .o1(new_n175));
  aob012aa1n02x5               g080(.a(new_n175), .b(new_n157), .c(new_n174), .out0(new_n176));
  nand22aa1n12x5               g081(.a(new_n174), .b(new_n159), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  nano32aa1n03x7               g083(.a(new_n122), .b(new_n178), .c(new_n135), .d(new_n137), .out0(new_n179));
  norp02aa1n02x5               g084(.a(new_n179), .b(new_n176), .o1(new_n180));
  nor042aa1n12x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  nand42aa1n10x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  xnbna2aa1n03x5               g088(.a(new_n180), .b(new_n183), .c(new_n182), .out0(\s[15] ));
  oaoi13aa1n06x5               g089(.a(new_n181), .b(new_n183), .c(new_n179), .d(new_n176), .o1(new_n185));
  xnrb03aa1n02x5               g090(.a(new_n185), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor002aa1n04x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nand42aa1n04x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  nano23aa1d15x5               g093(.a(new_n181), .b(new_n187), .c(new_n188), .d(new_n183), .out0(new_n189));
  aoi112aa1n02x5               g094(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n190));
  inv000aa1n02x5               g095(.a(new_n175), .o1(new_n191));
  nand22aa1n02x5               g096(.a(new_n189), .b(new_n191), .o1(new_n192));
  nona22aa1n03x5               g097(.a(new_n192), .b(new_n190), .c(new_n187), .out0(new_n193));
  aoi013aa1n09x5               g098(.a(new_n193), .b(new_n157), .c(new_n174), .d(new_n189), .o1(new_n194));
  nano32aa1d12x5               g099(.a(new_n177), .b(new_n189), .c(new_n135), .d(new_n137), .out0(new_n195));
  aoai13aa1n12x5               g100(.a(new_n195), .b(new_n121), .c(new_n117), .d(new_n106), .o1(new_n196));
  xnrc02aa1n12x5               g101(.a(\b[16] ), .b(\a[17] ), .out0(new_n197));
  xobna2aa1n03x5               g102(.a(new_n197), .b(new_n194), .c(new_n196), .out0(\s[17] ));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  nanp02aa1n09x5               g104(.a(new_n194), .b(new_n196), .o1(new_n200));
  norp02aa1n02x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  aoib12aa1n06x5               g106(.a(new_n201), .b(new_n200), .c(new_n197), .out0(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[17] ), .c(new_n199), .out0(\s[18] ));
  xnrc02aa1n02x5               g108(.a(\b[17] ), .b(\a[18] ), .out0(new_n204));
  norp02aa1n02x5               g109(.a(new_n204), .b(new_n197), .o1(new_n205));
  inv000aa1n02x5               g110(.a(new_n205), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[17] ), .o1(new_n207));
  oao003aa1n02x5               g112(.a(new_n199), .b(new_n207), .c(new_n201), .carry(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n206), .c(new_n194), .d(new_n196), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nanp02aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  nor042aa1n04x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nanp02aa1n04x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  norb02aa1n06x4               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  aoi112aa1n03x4               g122(.a(new_n213), .b(new_n217), .c(new_n210), .d(new_n214), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n217), .b(new_n213), .c(new_n210), .d(new_n214), .o1(new_n219));
  norb02aa1n02x7               g124(.a(new_n219), .b(new_n218), .out0(\s[20] ));
  nano23aa1n03x7               g125(.a(new_n213), .b(new_n215), .c(new_n216), .d(new_n214), .out0(new_n221));
  nona22aa1n02x4               g126(.a(new_n221), .b(new_n204), .c(new_n197), .out0(new_n222));
  aoi112aa1n02x5               g127(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n223));
  norp02aa1n02x5               g128(.a(\b[17] ), .b(\a[18] ), .o1(new_n224));
  aoi112aa1n09x5               g129(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n225));
  norb02aa1n02x7               g130(.a(new_n214), .b(new_n213), .out0(new_n226));
  oai112aa1n06x5               g131(.a(new_n226), .b(new_n217), .c(new_n225), .d(new_n224), .o1(new_n227));
  nona22aa1d18x5               g132(.a(new_n227), .b(new_n223), .c(new_n215), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n04x5               g134(.a(new_n229), .b(new_n222), .c(new_n194), .d(new_n196), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n04x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nanp02aa1n04x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  nor022aa1n08x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  nanp02aa1n06x5               g140(.a(\b[21] ), .b(\a[22] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  aoi112aa1n02x5               g142(.a(new_n232), .b(new_n237), .c(new_n230), .d(new_n234), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n237), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n239));
  norb02aa1n02x7               g144(.a(new_n239), .b(new_n238), .out0(\s[22] ));
  nano23aa1n06x5               g145(.a(new_n232), .b(new_n235), .c(new_n236), .d(new_n233), .out0(new_n241));
  aoi012aa1n02x5               g146(.a(new_n235), .b(new_n232), .c(new_n236), .o1(new_n242));
  aobi12aa1n02x5               g147(.a(new_n242), .b(new_n228), .c(new_n241), .out0(new_n243));
  nona23aa1n02x4               g148(.a(new_n221), .b(new_n241), .c(new_n204), .d(new_n197), .out0(new_n244));
  aoai13aa1n04x5               g149(.a(new_n243), .b(new_n244), .c(new_n194), .d(new_n196), .o1(new_n245));
  xorb03aa1n02x5               g150(.a(new_n245), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n09x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  nand22aa1n04x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  nor042aa1n09x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  nand02aa1n03x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  aoi122aa1n03x5               g156(.a(new_n247), .b(new_n250), .c(new_n251), .d(new_n245), .e(new_n248), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n247), .o1(new_n253));
  nanb02aa1n12x5               g158(.a(new_n247), .b(new_n248), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  nand02aa1n02x5               g160(.a(new_n245), .b(new_n255), .o1(new_n256));
  nanb02aa1n02x5               g161(.a(new_n249), .b(new_n251), .out0(new_n257));
  tech160nm_fiaoi012aa1n03p5x5 g162(.a(new_n257), .b(new_n256), .c(new_n253), .o1(new_n258));
  nor002aa1n02x5               g163(.a(new_n258), .b(new_n252), .o1(\s[24] ));
  nona23aa1n09x5               g164(.a(new_n251), .b(new_n248), .c(new_n247), .d(new_n249), .out0(new_n260));
  inv040aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  nanb03aa1n02x5               g166(.a(new_n222), .b(new_n261), .c(new_n241), .out0(new_n262));
  nanp02aa1n02x5               g167(.a(new_n247), .b(new_n251), .o1(new_n263));
  oai112aa1n03x5               g168(.a(new_n263), .b(new_n250), .c(new_n260), .d(new_n242), .o1(new_n264));
  nano22aa1n06x5               g169(.a(new_n260), .b(new_n234), .c(new_n237), .out0(new_n265));
  aoi012aa1n02x5               g170(.a(new_n264), .b(new_n228), .c(new_n265), .o1(new_n266));
  aoai13aa1n04x5               g171(.a(new_n266), .b(new_n262), .c(new_n194), .d(new_n196), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  xorc02aa1n03x5               g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xorc02aa1n02x5               g175(.a(\a[26] ), .b(\b[25] ), .out0(new_n271));
  aoi112aa1n02x5               g176(.a(new_n269), .b(new_n271), .c(new_n267), .d(new_n270), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n270), .o1(new_n273));
  norb02aa1n02x7               g178(.a(new_n273), .b(new_n272), .out0(\s[26] ));
  inv000aa1n02x5               g179(.a(new_n193), .o1(new_n275));
  nona23aa1n02x4               g180(.a(new_n188), .b(new_n183), .c(new_n181), .d(new_n187), .out0(new_n276));
  nona32aa1n06x5               g181(.a(new_n157), .b(new_n276), .c(new_n169), .d(new_n164), .out0(new_n277));
  tech160nm_finand02aa1n03p5x5 g182(.a(new_n277), .b(new_n275), .o1(new_n278));
  nano32aa1n03x7               g183(.a(new_n244), .b(new_n271), .c(new_n261), .d(new_n270), .out0(new_n279));
  aoai13aa1n06x5               g184(.a(new_n279), .b(new_n278), .c(new_n134), .d(new_n195), .o1(new_n280));
  norp02aa1n02x5               g185(.a(\b[25] ), .b(\a[26] ), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n281), .o1(new_n282));
  aoi112aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n283));
  inv000aa1n02x5               g188(.a(new_n283), .o1(new_n284));
  nor043aa1n02x5               g189(.a(new_n242), .b(new_n254), .c(new_n257), .o1(new_n285));
  nano22aa1n02x5               g190(.a(new_n285), .b(new_n250), .c(new_n263), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n228), .b(new_n265), .o1(new_n287));
  and002aa1n09x5               g192(.a(new_n271), .b(new_n270), .o(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  tech160nm_fiaoi012aa1n04x5   g194(.a(new_n289), .b(new_n287), .c(new_n286), .o1(new_n290));
  nano22aa1n03x7               g195(.a(new_n290), .b(new_n282), .c(new_n284), .out0(new_n291));
  xorc02aa1n12x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  xnbna2aa1n03x5               g197(.a(new_n292), .b(new_n280), .c(new_n291), .out0(\s[27] ));
  norp02aa1n02x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv040aa1n03x5               g199(.a(new_n294), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n292), .o1(new_n296));
  aoi012aa1n02x5               g201(.a(new_n296), .b(new_n280), .c(new_n291), .o1(new_n297));
  tech160nm_fixnrc02aa1n04x5   g202(.a(\b[27] ), .b(\a[28] ), .out0(new_n298));
  nano22aa1n02x4               g203(.a(new_n297), .b(new_n295), .c(new_n298), .out0(new_n299));
  aoai13aa1n02x5               g204(.a(new_n288), .b(new_n264), .c(new_n228), .d(new_n265), .o1(new_n300));
  nona22aa1n03x5               g205(.a(new_n300), .b(new_n283), .c(new_n281), .out0(new_n301));
  aoai13aa1n03x5               g206(.a(new_n292), .b(new_n301), .c(new_n200), .d(new_n279), .o1(new_n302));
  aoi012aa1n03x5               g207(.a(new_n298), .b(new_n302), .c(new_n295), .o1(new_n303));
  norp02aa1n03x5               g208(.a(new_n303), .b(new_n299), .o1(\s[28] ));
  norb02aa1d21x5               g209(.a(new_n292), .b(new_n298), .out0(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n301), .c(new_n200), .d(new_n279), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[28] ), .b(\a[29] ), .out0(new_n308));
  aoi012aa1n03x5               g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n305), .o1(new_n310));
  aoi012aa1n06x5               g215(.a(new_n310), .b(new_n280), .c(new_n291), .o1(new_n311));
  nano22aa1n02x5               g216(.a(new_n311), .b(new_n307), .c(new_n308), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n309), .b(new_n312), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g219(.a(new_n292), .b(new_n308), .c(new_n298), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n301), .c(new_n200), .d(new_n279), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n307), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .out0(new_n318));
  aoi012aa1n03x5               g223(.a(new_n318), .b(new_n316), .c(new_n317), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n315), .o1(new_n320));
  tech160nm_fiaoi012aa1n02p5x5 g225(.a(new_n320), .b(new_n280), .c(new_n291), .o1(new_n321));
  nano22aa1n02x4               g226(.a(new_n321), .b(new_n317), .c(new_n318), .out0(new_n322));
  nor002aa1n02x5               g227(.a(new_n319), .b(new_n322), .o1(\s[30] ));
  norb02aa1n09x5               g228(.a(new_n315), .b(new_n318), .out0(new_n324));
  inv030aa1n02x5               g229(.a(new_n324), .o1(new_n325));
  aoi012aa1n02x7               g230(.a(new_n325), .b(new_n280), .c(new_n291), .o1(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n327));
  xnrc02aa1n02x5               g232(.a(\b[30] ), .b(\a[31] ), .out0(new_n328));
  nano22aa1n02x4               g233(.a(new_n326), .b(new_n327), .c(new_n328), .out0(new_n329));
  aoai13aa1n03x5               g234(.a(new_n324), .b(new_n301), .c(new_n200), .d(new_n279), .o1(new_n330));
  aoi012aa1n03x5               g235(.a(new_n328), .b(new_n330), .c(new_n327), .o1(new_n331));
  nor002aa1n02x5               g236(.a(new_n331), .b(new_n329), .o1(\s[31] ));
  xnrb03aa1n02x5               g237(.a(new_n110), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g238(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g240(.a(new_n117), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g241(.a(\a[5] ), .b(\b[4] ), .c(new_n131), .o1(new_n337));
  xorb03aa1n02x5               g242(.a(new_n337), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g243(.a(new_n100), .b(new_n101), .c(new_n337), .d(new_n102), .o1(new_n339));
  aoi112aa1n02x5               g244(.a(new_n100), .b(new_n101), .c(new_n337), .d(new_n102), .o1(new_n340));
  norb02aa1n02x5               g245(.a(new_n339), .b(new_n340), .out0(\s[7] ));
  orn002aa1n02x5               g246(.a(\a[7] ), .b(\b[6] ), .o(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n99), .b(new_n339), .c(new_n342), .out0(\s[8] ));
  xnrc02aa1n02x5               g248(.a(new_n122), .b(new_n135), .out0(\s[9] ));
endmodule


