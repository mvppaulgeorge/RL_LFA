// Benchmark "adder" written by ABC on Thu Jul 18 11:54:23 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n317,
    new_n318, new_n320, new_n321, new_n322, new_n324, new_n325, new_n326,
    new_n328, new_n330, new_n331, new_n332;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nand42aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[4] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[3] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  aoi012aa1n02x5               g007(.a(new_n102), .b(new_n100), .c(new_n101), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb02aa1n06x5               g009(.a(new_n102), .b(new_n104), .out0(new_n105));
  nanp02aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nand22aa1n04x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  nor042aa1n02x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  tech160nm_fioai012aa1n05x5   g013(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n109));
  tech160nm_fioai012aa1n05x5   g014(.a(new_n103), .b(new_n109), .c(new_n105), .o1(new_n110));
  aoi022aa1n02x7               g015(.a(\b[7] ), .b(\a[8] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n111));
  nor022aa1n08x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor022aa1n16x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n03x5               g019(.a(new_n111), .b(new_n114), .c(new_n113), .d(new_n112), .out0(new_n115));
  nanp02aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nor022aa1n16x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nor002aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand02aa1d04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nona23aa1n03x5               g024(.a(new_n116), .b(new_n119), .c(new_n118), .d(new_n117), .out0(new_n120));
  nona22aa1n06x5               g025(.a(new_n110), .b(new_n115), .c(new_n120), .out0(new_n121));
  inv000aa1d42x5               g026(.a(new_n113), .o1(new_n122));
  tech160nm_fioai012aa1n05x5   g027(.a(new_n119), .b(new_n117), .c(new_n112), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n123), .b(new_n122), .o1(new_n124));
  aoi022aa1n02x5               g029(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n125));
  tech160nm_fiaoi012aa1n04x5   g030(.a(new_n118), .b(new_n124), .c(new_n125), .o1(new_n126));
  tech160nm_fixnrc02aa1n04x5   g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n99), .b(new_n127), .c(new_n121), .d(new_n126), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n08x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nanb02aa1n12x5               g036(.a(new_n130), .b(new_n131), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  oaoi03aa1n03x5               g038(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanp02aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  aoai13aa1n06x5               g043(.a(new_n138), .b(new_n134), .c(new_n128), .d(new_n133), .o1(new_n139));
  aoi112aa1n02x5               g044(.a(new_n138), .b(new_n134), .c(new_n128), .d(new_n133), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(\s[11] ));
  inv040aa1n03x5               g046(.a(new_n135), .o1(new_n142));
  norp02aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanp02aa1n04x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n139), .c(new_n142), .out0(\s[12] ));
  nor002aa1n02x5               g051(.a(new_n120), .b(new_n115), .o1(new_n147));
  oaoi13aa1n06x5               g052(.a(new_n113), .b(new_n119), .c(new_n117), .d(new_n112), .o1(new_n148));
  obai22aa1n02x7               g053(.a(new_n125), .b(new_n148), .c(\a[8] ), .d(\b[7] ), .out0(new_n149));
  nona23aa1d18x5               g054(.a(new_n144), .b(new_n136), .c(new_n135), .d(new_n143), .out0(new_n150));
  norp03aa1n02x5               g055(.a(new_n150), .b(new_n132), .c(new_n127), .o1(new_n151));
  aoai13aa1n03x5               g056(.a(new_n151), .b(new_n149), .c(new_n147), .d(new_n110), .o1(new_n152));
  aoai13aa1n04x5               g057(.a(new_n131), .b(new_n130), .c(new_n97), .d(new_n98), .o1(new_n153));
  oaoi03aa1n09x5               g058(.a(\a[12] ), .b(\b[11] ), .c(new_n142), .o1(new_n154));
  oabi12aa1n18x5               g059(.a(new_n154), .b(new_n150), .c(new_n153), .out0(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nand22aa1n03x5               g061(.a(new_n152), .b(new_n156), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n03x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1n06x5               g069(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n165));
  tech160nm_fiaoi012aa1n04x5   g070(.a(new_n163), .b(new_n159), .c(new_n164), .o1(new_n166));
  inv000aa1n02x5               g071(.a(new_n166), .o1(new_n167));
  nor022aa1n04x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nanp02aa1n04x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n167), .c(new_n157), .d(new_n165), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n170), .b(new_n167), .c(new_n157), .d(new_n165), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[15] ));
  nor022aa1n06x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  tech160nm_fioai012aa1n03p5x5 g080(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .o1(new_n176));
  oaib12aa1n02x5               g081(.a(new_n176), .b(new_n174), .c(new_n175), .out0(new_n177));
  nona23aa1n02x4               g082(.a(new_n171), .b(new_n175), .c(new_n174), .d(new_n168), .out0(new_n178));
  nanp02aa1n02x5               g083(.a(new_n177), .b(new_n178), .o1(\s[16] ));
  inv000aa1d42x5               g084(.a(\a[17] ), .o1(new_n180));
  nona23aa1d18x5               g085(.a(new_n175), .b(new_n169), .c(new_n168), .d(new_n174), .out0(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  nor042aa1n02x5               g087(.a(new_n127), .b(new_n132), .o1(new_n183));
  nona23aa1n09x5               g088(.a(new_n165), .b(new_n183), .c(new_n181), .d(new_n150), .out0(new_n184));
  aoi012aa1n06x5               g089(.a(new_n184), .b(new_n121), .c(new_n126), .o1(new_n185));
  nano23aa1n03x5               g090(.a(new_n135), .b(new_n143), .c(new_n144), .d(new_n136), .out0(new_n186));
  aoai13aa1n02x5               g091(.a(new_n165), .b(new_n154), .c(new_n186), .d(new_n134), .o1(new_n187));
  nanp02aa1n03x5               g092(.a(new_n187), .b(new_n166), .o1(new_n188));
  oa0012aa1n06x5               g093(.a(new_n175), .b(new_n174), .c(new_n168), .o(new_n189));
  aoi112aa1n09x5               g094(.a(new_n185), .b(new_n189), .c(new_n188), .d(new_n182), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(new_n180), .out0(\s[17] ));
  oaoi03aa1n03x5               g096(.a(\a[17] ), .b(\b[16] ), .c(new_n190), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g098(.a(\a[18] ), .o1(new_n194));
  xroi22aa1d06x4               g099(.a(new_n180), .b(\b[16] ), .c(new_n194), .d(\b[17] ), .out0(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  oai022aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oaib12aa1n02x5               g102(.a(new_n197), .b(new_n194), .c(\b[17] ), .out0(new_n198));
  oai012aa1n06x5               g103(.a(new_n198), .b(new_n190), .c(new_n196), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand02aa1d04x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  nor042aa1n04x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand02aa1d04x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nanb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(new_n207));
  aoai13aa1n03x5               g112(.a(new_n207), .b(new_n202), .c(new_n199), .d(new_n204), .o1(new_n208));
  tech160nm_fiaoi012aa1n05x5   g113(.a(new_n149), .b(new_n147), .c(new_n110), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n182), .b(new_n167), .c(new_n155), .d(new_n165), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n189), .o1(new_n211));
  oai112aa1n06x5               g116(.a(new_n210), .b(new_n211), .c(new_n209), .d(new_n184), .o1(new_n212));
  nanb02aa1n02x5               g117(.a(\b[16] ), .b(new_n180), .out0(new_n213));
  oaoi03aa1n02x5               g118(.a(\a[18] ), .b(\b[17] ), .c(new_n213), .o1(new_n214));
  aoai13aa1n03x5               g119(.a(new_n204), .b(new_n214), .c(new_n212), .d(new_n195), .o1(new_n215));
  nona22aa1n02x4               g120(.a(new_n215), .b(new_n207), .c(new_n202), .out0(new_n216));
  nanp02aa1n03x5               g121(.a(new_n208), .b(new_n216), .o1(\s[20] ));
  nona23aa1n09x5               g122(.a(new_n206), .b(new_n203), .c(new_n202), .d(new_n205), .out0(new_n218));
  norb02aa1n02x5               g123(.a(new_n195), .b(new_n218), .out0(new_n219));
  inv020aa1n02x5               g124(.a(new_n219), .o1(new_n220));
  tech160nm_fiao0012aa1n02p5x5 g125(.a(new_n205), .b(new_n202), .c(new_n206), .o(new_n221));
  oabi12aa1n06x5               g126(.a(new_n221), .b(new_n218), .c(new_n198), .out0(new_n222));
  oabi12aa1n06x5               g127(.a(new_n222), .b(new_n190), .c(new_n220), .out0(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  tech160nm_fixnrc02aa1n05x5   g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  aoai13aa1n03x5               g133(.a(new_n228), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n227), .b(new_n222), .c(new_n212), .d(new_n219), .o1(new_n230));
  nona22aa1n02x4               g135(.a(new_n230), .b(new_n228), .c(new_n225), .out0(new_n231));
  nanp02aa1n03x5               g136(.a(new_n229), .b(new_n231), .o1(\s[22] ));
  nano23aa1d15x5               g137(.a(new_n202), .b(new_n205), .c(new_n206), .d(new_n203), .out0(new_n233));
  nor022aa1n08x5               g138(.a(new_n228), .b(new_n226), .o1(new_n234));
  nand23aa1d12x5               g139(.a(new_n195), .b(new_n234), .c(new_n233), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n234), .b(new_n221), .c(new_n233), .d(new_n214), .o1(new_n236));
  inv000aa1d42x5               g141(.a(\a[22] ), .o1(new_n237));
  inv000aa1d42x5               g142(.a(\b[21] ), .o1(new_n238));
  oao003aa1n06x5               g143(.a(new_n237), .b(new_n238), .c(new_n225), .carry(new_n239));
  inv000aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  nanp02aa1n02x5               g145(.a(new_n236), .b(new_n240), .o1(new_n241));
  oabi12aa1n06x5               g146(.a(new_n241), .b(new_n190), .c(new_n235), .out0(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  tech160nm_fixnrc02aa1n05x5   g150(.a(\b[23] ), .b(\a[24] ), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n244), .c(new_n242), .d(new_n245), .o1(new_n247));
  inv040aa1n03x5               g152(.a(new_n235), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n245), .b(new_n241), .c(new_n212), .d(new_n248), .o1(new_n249));
  nona22aa1n03x5               g154(.a(new_n249), .b(new_n246), .c(new_n244), .out0(new_n250));
  nanp02aa1n03x5               g155(.a(new_n247), .b(new_n250), .o1(\s[24] ));
  norb02aa1n02x5               g156(.a(new_n245), .b(new_n246), .out0(new_n252));
  inv030aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  nano32aa1n03x7               g158(.a(new_n253), .b(new_n195), .c(new_n234), .d(new_n233), .out0(new_n254));
  inv020aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  oai022aa1n02x5               g160(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n256));
  aob012aa1n02x5               g161(.a(new_n256), .b(\b[23] ), .c(\a[24] ), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n253), .c(new_n236), .d(new_n240), .o1(new_n258));
  oabi12aa1n06x5               g163(.a(new_n258), .b(new_n190), .c(new_n255), .out0(new_n259));
  xorb03aa1n02x5               g164(.a(new_n259), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  xorc02aa1n03x5               g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xorc02aa1n12x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n261), .c(new_n259), .d(new_n262), .o1(new_n265));
  aoai13aa1n02x5               g170(.a(new_n262), .b(new_n258), .c(new_n212), .d(new_n254), .o1(new_n266));
  nona22aa1n02x4               g171(.a(new_n266), .b(new_n264), .c(new_n261), .out0(new_n267));
  nanp02aa1n03x5               g172(.a(new_n265), .b(new_n267), .o1(\s[26] ));
  and002aa1n12x5               g173(.a(new_n263), .b(new_n262), .o(new_n269));
  nano22aa1d15x5               g174(.a(new_n235), .b(new_n269), .c(new_n252), .out0(new_n270));
  nand02aa1d08x5               g175(.a(new_n212), .b(new_n270), .o1(new_n271));
  nanp02aa1n02x5               g176(.a(\b[25] ), .b(\a[26] ), .o1(new_n272));
  oai022aa1n02x5               g177(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n273));
  aoi022aa1n06x5               g178(.a(new_n258), .b(new_n269), .c(new_n272), .d(new_n273), .o1(new_n274));
  xorc02aa1n12x5               g179(.a(\a[27] ), .b(\b[26] ), .out0(new_n275));
  xnbna2aa1n06x5               g180(.a(new_n275), .b(new_n271), .c(new_n274), .out0(\s[27] ));
  inv020aa1n03x5               g181(.a(new_n270), .o1(new_n277));
  tech160nm_fioai012aa1n03p5x5 g182(.a(new_n274), .b(new_n190), .c(new_n277), .o1(new_n278));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  norp02aa1n04x5               g184(.a(\b[27] ), .b(\a[28] ), .o1(new_n280));
  nanp02aa1n04x5               g185(.a(\b[27] ), .b(\a[28] ), .o1(new_n281));
  nanb02aa1n06x5               g186(.a(new_n280), .b(new_n281), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n282), .b(new_n279), .c(new_n278), .d(new_n275), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n252), .b(new_n239), .c(new_n222), .d(new_n234), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n269), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n273), .b(new_n272), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n286), .b(new_n285), .c(new_n284), .d(new_n257), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n275), .b(new_n287), .c(new_n212), .d(new_n270), .o1(new_n288));
  nona22aa1n02x5               g193(.a(new_n288), .b(new_n282), .c(new_n279), .out0(new_n289));
  nanp02aa1n03x5               g194(.a(new_n283), .b(new_n289), .o1(\s[28] ));
  norb02aa1n02x7               g195(.a(new_n275), .b(new_n282), .out0(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n287), .c(new_n212), .d(new_n270), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n291), .o1(new_n293));
  aoi012aa1n02x5               g198(.a(new_n280), .b(new_n279), .c(new_n281), .o1(new_n294));
  aoai13aa1n02x7               g199(.a(new_n294), .b(new_n293), .c(new_n271), .d(new_n274), .o1(new_n295));
  tech160nm_fixorc02aa1n03p5x5 g200(.a(\a[29] ), .b(\b[28] ), .out0(new_n296));
  norb02aa1n02x5               g201(.a(new_n294), .b(new_n296), .out0(new_n297));
  aoi022aa1n02x7               g202(.a(new_n295), .b(new_n296), .c(new_n292), .d(new_n297), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g204(.a(new_n282), .b(new_n275), .c(new_n296), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n287), .c(new_n212), .d(new_n270), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n300), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .carry(new_n303));
  aoai13aa1n02x7               g208(.a(new_n303), .b(new_n302), .c(new_n271), .d(new_n274), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .out0(new_n305));
  norb02aa1n02x5               g210(.a(new_n303), .b(new_n305), .out0(new_n306));
  aoi022aa1n02x7               g211(.a(new_n304), .b(new_n305), .c(new_n301), .d(new_n306), .o1(\s[30] ));
  nand03aa1n02x5               g212(.a(new_n291), .b(new_n296), .c(new_n305), .o1(new_n308));
  nanb02aa1n03x5               g213(.a(new_n308), .b(new_n278), .out0(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n303), .carry(new_n310));
  aoai13aa1n02x7               g215(.a(new_n310), .b(new_n308), .c(new_n271), .d(new_n274), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[31] ), .b(\b[30] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n309), .d(new_n313), .o1(\s[31] ));
  xnrb03aa1n02x5               g219(.a(new_n109), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  orn002aa1n02x5               g220(.a(new_n109), .b(new_n105), .o(new_n316));
  xorc02aa1n02x5               g221(.a(\a[4] ), .b(\b[3] ), .out0(new_n317));
  norp02aa1n02x5               g222(.a(new_n317), .b(new_n102), .o1(new_n318));
  aoi022aa1n02x5               g223(.a(new_n316), .b(new_n318), .c(new_n110), .d(new_n317), .o1(\s[4] ));
  norb02aa1n02x5               g224(.a(new_n116), .b(new_n117), .out0(new_n320));
  oaoi13aa1n02x5               g225(.a(new_n320), .b(new_n110), .c(new_n100), .d(new_n101), .o1(new_n321));
  oai112aa1n03x5               g226(.a(new_n110), .b(new_n320), .c(new_n101), .d(new_n100), .o1(new_n322));
  norb02aa1n02x5               g227(.a(new_n322), .b(new_n321), .out0(\s[5] ));
  nanb02aa1n02x5               g228(.a(new_n112), .b(new_n119), .out0(new_n324));
  oaoi13aa1n04x5               g229(.a(new_n324), .b(new_n322), .c(\a[5] ), .d(\b[4] ), .o1(new_n325));
  oai112aa1n02x5               g230(.a(new_n322), .b(new_n324), .c(\b[4] ), .d(\a[5] ), .o1(new_n326));
  norb02aa1n02x5               g231(.a(new_n326), .b(new_n325), .out0(\s[6] ));
  nanb02aa1n06x5               g232(.a(new_n325), .b(new_n123), .out0(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aob012aa1n02x5               g234(.a(new_n122), .b(new_n328), .c(new_n114), .out0(new_n330));
  xorc02aa1n02x5               g235(.a(\a[8] ), .b(\b[7] ), .out0(new_n331));
  aoi112aa1n02x5               g236(.a(new_n331), .b(new_n113), .c(new_n328), .d(new_n114), .o1(new_n332));
  aoi012aa1n03x5               g237(.a(new_n332), .b(new_n330), .c(new_n331), .o1(\s[8] ));
  xobna2aa1n03x5               g238(.a(new_n127), .b(new_n121), .c(new_n126), .out0(\s[9] ));
endmodule


