// Benchmark "adder" written by ABC on Thu Jul 18 12:01:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n318, new_n320, new_n321, new_n322, new_n324, new_n325,
    new_n327, new_n329, new_n330, new_n332, new_n333, new_n334, new_n335,
    new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  oa0022aa1n02x5               g003(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n99));
  tech160nm_fixnrc02aa1n04x5   g004(.a(\b[2] ), .b(\a[3] ), .out0(new_n100));
  nand42aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1d24x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  nor042aa1n09x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oaih12aa1n06x5               g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  oai012aa1n12x5               g009(.a(new_n99), .b(new_n100), .c(new_n104), .o1(new_n105));
  inv000aa1d42x5               g010(.a(\a[8] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[7] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  orn002aa1n03x5               g013(.a(\a[5] ), .b(\b[4] ), .o(new_n109));
  oai112aa1n03x5               g014(.a(new_n109), .b(new_n108), .c(new_n107), .d(new_n106), .o1(new_n110));
  nand02aa1n04x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  inv040aa1d32x5               g016(.a(\a[7] ), .o1(new_n112));
  inv030aa1d32x5               g017(.a(\b[6] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(new_n113), .b(new_n112), .o1(new_n114));
  nand22aa1n06x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand03aa1n02x5               g020(.a(new_n114), .b(new_n111), .c(new_n115), .o1(new_n116));
  nand42aa1n02x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  oai122aa1n02x5               g022(.a(new_n117), .b(\a[8] ), .c(\b[7] ), .d(\a[6] ), .e(\b[5] ), .o1(new_n118));
  nor043aa1n03x5               g023(.a(new_n110), .b(new_n116), .c(new_n118), .o1(new_n119));
  and002aa1n02x5               g024(.a(\b[7] ), .b(\a[8] ), .o(new_n120));
  nanp02aa1n02x5               g025(.a(new_n107), .b(new_n106), .o1(new_n121));
  oai022aa1d18x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  nanp03aa1n06x5               g027(.a(new_n122), .b(new_n111), .c(new_n115), .o1(new_n123));
  aoai13aa1n04x5               g028(.a(new_n121), .b(new_n120), .c(new_n123), .d(new_n114), .o1(new_n124));
  tech160nm_fixorc02aa1n05x5   g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n105), .d(new_n119), .o1(new_n126));
  nor002aa1n12x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand02aa1d08x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n06x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  nanp02aa1n02x5               g035(.a(new_n119), .b(new_n105), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n124), .b(new_n131), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n129), .b(new_n97), .c(new_n132), .d(new_n125), .o1(new_n133));
  oai012aa1d24x5               g038(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n134));
  nor002aa1d24x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanp02aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n136), .b(new_n135), .out0(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n137), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  inv000aa1d42x5               g043(.a(new_n137), .o1(new_n139));
  aoi012aa1n02x5               g044(.a(new_n139), .b(new_n133), .c(new_n134), .o1(new_n140));
  nor002aa1d32x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand02aa1d08x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanb02aa1n02x5               g047(.a(new_n141), .b(new_n142), .out0(new_n143));
  oai012aa1n02x5               g048(.a(new_n143), .b(new_n140), .c(new_n135), .o1(new_n144));
  norb03aa1n02x5               g049(.a(new_n142), .b(new_n135), .c(new_n141), .out0(new_n145));
  oaib12aa1n02x5               g050(.a(new_n144), .b(new_n140), .c(new_n145), .out0(\s[12] ));
  nona23aa1d18x5               g051(.a(new_n142), .b(new_n136), .c(new_n135), .d(new_n141), .out0(new_n147));
  nano22aa1n03x7               g052(.a(new_n147), .b(new_n125), .c(new_n129), .out0(new_n148));
  aoai13aa1n02x5               g053(.a(new_n148), .b(new_n124), .c(new_n105), .d(new_n119), .o1(new_n149));
  oai012aa1d24x5               g054(.a(new_n142), .b(new_n141), .c(new_n135), .o1(new_n150));
  oai012aa1d24x5               g055(.a(new_n150), .b(new_n147), .c(new_n134), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  xorc02aa1n02x5               g057(.a(\a[13] ), .b(\b[12] ), .out0(new_n153));
  xnbna2aa1n03x5               g058(.a(new_n153), .b(new_n149), .c(new_n152), .out0(\s[13] ));
  nor042aa1n09x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(new_n149), .b(new_n152), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(new_n157), .b(new_n153), .o1(new_n158));
  xorc02aa1n02x5               g063(.a(\a[14] ), .b(\b[13] ), .out0(new_n159));
  inv040aa1d32x5               g064(.a(\a[14] ), .o1(new_n160));
  inv000aa1d42x5               g065(.a(\b[13] ), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n155), .b(new_n160), .c(new_n161), .o1(new_n162));
  oai112aa1n02x5               g067(.a(new_n158), .b(new_n162), .c(new_n161), .d(new_n160), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n159), .c(new_n156), .d(new_n158), .o1(\s[14] ));
  inv000aa1d42x5               g069(.a(\a[13] ), .o1(new_n165));
  xroi22aa1d06x4               g070(.a(new_n165), .b(\b[12] ), .c(new_n160), .d(\b[13] ), .out0(new_n166));
  oaoi03aa1n12x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n167));
  xorc02aa1n12x5               g072(.a(\a[15] ), .b(\b[14] ), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n167), .c(new_n157), .d(new_n166), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n168), .b(new_n167), .c(new_n157), .d(new_n166), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n169), .b(new_n170), .out0(\s[15] ));
  nor042aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  xorc02aa1n12x5               g078(.a(\a[16] ), .b(\b[15] ), .out0(new_n174));
  inv000aa1d42x5               g079(.a(\a[16] ), .o1(new_n175));
  inv000aa1d42x5               g080(.a(\b[15] ), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n172), .b(new_n175), .c(new_n176), .o1(new_n177));
  oai112aa1n02x5               g082(.a(new_n169), .b(new_n177), .c(new_n176), .d(new_n175), .o1(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n174), .c(new_n173), .d(new_n169), .o1(\s[16] ));
  tech160nm_fiaoi012aa1n05x5   g084(.a(new_n124), .b(new_n105), .c(new_n119), .o1(new_n180));
  nanp02aa1n12x5               g085(.a(new_n174), .b(new_n168), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  nand23aa1n02x5               g087(.a(new_n148), .b(new_n182), .c(new_n166), .o1(new_n183));
  aoai13aa1n04x5               g088(.a(new_n182), .b(new_n167), .c(new_n151), .d(new_n166), .o1(new_n184));
  tech160nm_fioaoi03aa1n03p5x5 g089(.a(new_n175), .b(new_n176), .c(new_n172), .o1(new_n185));
  oai112aa1n06x5               g090(.a(new_n184), .b(new_n185), .c(new_n180), .d(new_n183), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g092(.a(\a[18] ), .o1(new_n188));
  nor002aa1n02x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  tech160nm_fiaoi012aa1n05x5   g095(.a(new_n189), .b(new_n186), .c(new_n190), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[17] ), .c(new_n188), .out0(\s[18] ));
  inv000aa1d42x5               g097(.a(\a[17] ), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n193), .b(\b[16] ), .c(new_n188), .d(\b[17] ), .out0(new_n194));
  aob012aa1n02x5               g099(.a(new_n189), .b(\b[17] ), .c(\a[18] ), .out0(new_n195));
  oaib12aa1n06x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n188), .out0(new_n196));
  nor042aa1n04x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  aoai13aa1n04x5               g104(.a(new_n199), .b(new_n196), .c(new_n186), .d(new_n194), .o1(new_n200));
  aoi112aa1n02x5               g105(.a(new_n199), .b(new_n196), .c(new_n186), .d(new_n194), .o1(new_n201));
  norb02aa1n03x4               g106(.a(new_n200), .b(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g108(.a(new_n197), .o1(new_n204));
  nor042aa1n02x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand02aa1n03x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  norb03aa1n02x5               g112(.a(new_n206), .b(new_n197), .c(new_n205), .out0(new_n208));
  nanp02aa1n03x5               g113(.a(new_n200), .b(new_n208), .o1(new_n209));
  aoai13aa1n03x5               g114(.a(new_n209), .b(new_n207), .c(new_n204), .d(new_n200), .o1(\s[20] ));
  nano23aa1n09x5               g115(.a(new_n197), .b(new_n205), .c(new_n206), .d(new_n198), .out0(new_n211));
  nand02aa1d04x5               g116(.a(new_n194), .b(new_n211), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  aoi112aa1n02x5               g118(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n214));
  aoib12aa1n02x5               g119(.a(new_n214), .b(new_n188), .c(\b[17] ), .out0(new_n215));
  nona23aa1n02x4               g120(.a(new_n206), .b(new_n198), .c(new_n197), .d(new_n205), .out0(new_n216));
  oaoi03aa1n02x5               g121(.a(\a[20] ), .b(\b[19] ), .c(new_n204), .o1(new_n217));
  oabi12aa1n06x5               g122(.a(new_n217), .b(new_n216), .c(new_n215), .out0(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n218), .c(new_n186), .d(new_n213), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(new_n220), .b(new_n218), .c(new_n186), .d(new_n213), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n221), .b(new_n222), .out0(\s[21] ));
  nor042aa1n06x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  inv020aa1n04x5               g129(.a(new_n224), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  and002aa1n02x5               g132(.a(\b[21] ), .b(\a[22] ), .o(new_n228));
  oai022aa1n02x5               g133(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n229));
  nona22aa1n03x5               g134(.a(new_n221), .b(new_n228), .c(new_n229), .out0(new_n230));
  aoai13aa1n03x5               g135(.a(new_n230), .b(new_n227), .c(new_n225), .d(new_n221), .o1(\s[22] ));
  nor042aa1n06x5               g136(.a(new_n226), .b(new_n219), .o1(new_n232));
  nanp03aa1d12x5               g137(.a(new_n194), .b(new_n232), .c(new_n211), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoai13aa1n06x5               g139(.a(new_n232), .b(new_n217), .c(new_n211), .d(new_n196), .o1(new_n235));
  oaoi03aa1n02x5               g140(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .o1(new_n236));
  inv000aa1n02x5               g141(.a(new_n236), .o1(new_n237));
  nanp02aa1n02x5               g142(.a(new_n235), .b(new_n237), .o1(new_n238));
  xorc02aa1n12x5               g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n238), .c(new_n186), .d(new_n234), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(new_n239), .b(new_n238), .c(new_n186), .d(new_n234), .o1(new_n241));
  norb02aa1n03x4               g146(.a(new_n240), .b(new_n241), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  tech160nm_fixorc02aa1n05x5   g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  and002aa1n02x5               g150(.a(\b[23] ), .b(\a[24] ), .o(new_n246));
  oai022aa1n02x5               g151(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n247));
  nona22aa1n03x5               g152(.a(new_n240), .b(new_n246), .c(new_n247), .out0(new_n248));
  aoai13aa1n03x5               g153(.a(new_n248), .b(new_n245), .c(new_n244), .d(new_n240), .o1(\s[24] ));
  nano32aa1n02x5               g154(.a(new_n212), .b(new_n245), .c(new_n232), .d(new_n239), .out0(new_n250));
  and002aa1n02x5               g155(.a(new_n245), .b(new_n239), .o(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  aob012aa1n02x5               g157(.a(new_n247), .b(\b[23] ), .c(\a[24] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n252), .c(new_n235), .d(new_n237), .o1(new_n254));
  tech160nm_fixorc02aa1n03p5x5 g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n186), .d(new_n250), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n255), .b(new_n254), .c(new_n186), .d(new_n250), .o1(new_n257));
  norb02aa1n03x4               g162(.a(new_n256), .b(new_n257), .out0(\s[25] ));
  norp02aa1n02x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  xorc02aa1n02x5               g165(.a(\a[26] ), .b(\b[25] ), .out0(new_n261));
  and002aa1n02x5               g166(.a(\b[25] ), .b(\a[26] ), .o(new_n262));
  oai022aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n263));
  nona22aa1n03x5               g168(.a(new_n256), .b(new_n262), .c(new_n263), .out0(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n261), .c(new_n260), .d(new_n256), .o1(\s[26] ));
  aoib12aa1n02x5               g170(.a(new_n183), .b(new_n131), .c(new_n124), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n167), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n134), .o1(new_n268));
  nano23aa1n02x4               g173(.a(new_n135), .b(new_n141), .c(new_n142), .d(new_n136), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n150), .o1(new_n270));
  aoai13aa1n02x5               g175(.a(new_n166), .b(new_n270), .c(new_n269), .d(new_n268), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n185), .b(new_n181), .c(new_n271), .d(new_n267), .o1(new_n272));
  and002aa1n06x5               g177(.a(new_n261), .b(new_n255), .o(new_n273));
  nano22aa1d15x5               g178(.a(new_n233), .b(new_n251), .c(new_n273), .out0(new_n274));
  tech160nm_fioai012aa1n05x5   g179(.a(new_n274), .b(new_n272), .c(new_n266), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n262), .o1(new_n276));
  aoi022aa1n06x5               g181(.a(new_n254), .b(new_n273), .c(new_n276), .d(new_n263), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnbna2aa1n06x5               g183(.a(new_n278), .b(new_n275), .c(new_n277), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n251), .b(new_n236), .c(new_n218), .d(new_n232), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n273), .o1(new_n283));
  aob012aa1n02x5               g188(.a(new_n263), .b(\b[25] ), .c(\a[26] ), .out0(new_n284));
  aoai13aa1n04x5               g189(.a(new_n284), .b(new_n283), .c(new_n282), .d(new_n253), .o1(new_n285));
  aoai13aa1n04x5               g190(.a(new_n278), .b(new_n285), .c(new_n186), .d(new_n274), .o1(new_n286));
  xorc02aa1n02x5               g191(.a(\a[28] ), .b(\b[27] ), .out0(new_n287));
  inv000aa1d42x5               g192(.a(new_n278), .o1(new_n288));
  oai022aa1n02x5               g193(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n289));
  aoi012aa1n02x5               g194(.a(new_n289), .b(\a[28] ), .c(\b[27] ), .o1(new_n290));
  aoai13aa1n04x5               g195(.a(new_n290), .b(new_n288), .c(new_n275), .d(new_n277), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n291), .b(new_n287), .c(new_n286), .d(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g197(.a(new_n287), .b(new_n278), .o(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n285), .c(new_n186), .d(new_n274), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n293), .o1(new_n295));
  aob012aa1n02x5               g200(.a(new_n289), .b(\b[27] ), .c(\a[28] ), .out0(new_n296));
  aoai13aa1n02x5               g201(.a(new_n296), .b(new_n295), .c(new_n275), .d(new_n277), .o1(new_n297));
  xorc02aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .out0(new_n298));
  norb02aa1n02x5               g203(.a(new_n296), .b(new_n298), .out0(new_n299));
  aoi022aa1n03x5               g204(.a(new_n297), .b(new_n298), .c(new_n294), .d(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g206(.a(new_n288), .b(new_n287), .c(new_n298), .out0(new_n302));
  aoai13aa1n02x5               g207(.a(new_n302), .b(new_n285), .c(new_n186), .d(new_n274), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n302), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n304), .c(new_n275), .d(new_n277), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[30] ));
  nano32aa1n03x7               g214(.a(new_n288), .b(new_n307), .c(new_n287), .d(new_n298), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n285), .c(new_n186), .d(new_n274), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n310), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n312), .c(new_n275), .d(new_n277), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[31] ), .b(\b[30] ), .out0(new_n315));
  norb02aa1n02x5               g220(.a(new_n313), .b(new_n315), .out0(new_n316));
  aoi022aa1n03x5               g221(.a(new_n314), .b(new_n315), .c(new_n311), .d(new_n316), .o1(\s[31] ));
  inv000aa1d42x5               g222(.a(\a[3] ), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n104), .b(\b[2] ), .c(new_n318), .out0(\s[3] ));
  norp02aa1n02x5               g224(.a(new_n100), .b(new_n104), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[4] ), .b(\b[3] ), .out0(new_n321));
  aoib12aa1n02x5               g226(.a(new_n321), .b(new_n318), .c(\b[2] ), .out0(new_n322));
  aboi22aa1n03x5               g227(.a(new_n320), .b(new_n322), .c(new_n105), .d(new_n321), .out0(\s[4] ));
  aoi022aa1n02x5               g228(.a(new_n105), .b(new_n117), .c(new_n108), .d(new_n109), .o1(new_n324));
  aoi022aa1n02x5               g229(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n325));
  aoi013aa1n02x4               g230(.a(new_n324), .b(new_n109), .c(new_n105), .d(new_n325), .o1(\s[5] ));
  aob012aa1n02x5               g231(.a(new_n109), .b(new_n105), .c(new_n325), .out0(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  xorc02aa1n02x5               g233(.a(\a[6] ), .b(\b[5] ), .out0(new_n329));
  ao0022aa1n03x5               g234(.a(new_n327), .b(new_n329), .c(new_n111), .d(new_n122), .o(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp03aa1n02x5               g236(.a(new_n330), .b(new_n114), .c(new_n115), .o1(new_n332));
  aob012aa1n02x5               g237(.a(new_n114), .b(new_n330), .c(new_n115), .out0(new_n333));
  xorc02aa1n02x5               g238(.a(\a[8] ), .b(\b[7] ), .out0(new_n334));
  aboi22aa1n03x5               g239(.a(new_n120), .b(new_n121), .c(new_n112), .d(new_n113), .out0(new_n335));
  aoi022aa1n02x5               g240(.a(new_n333), .b(new_n334), .c(new_n332), .d(new_n335), .o1(\s[8] ));
  norp02aa1n02x5               g241(.a(new_n124), .b(new_n125), .o1(new_n337));
  aoi022aa1n02x5               g242(.a(new_n132), .b(new_n125), .c(new_n131), .d(new_n337), .o1(\s[9] ));
endmodule


