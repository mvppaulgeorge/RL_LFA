// Benchmark "adder" written by ABC on Thu Jul 18 10:28:02 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n142, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n318, new_n319, new_n322, new_n324, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n20x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nor042aa1n04x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand02aa1d04x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oao003aa1n02x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .carry(new_n105));
  nor002aa1d32x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanp02aa1n04x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand42aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nano23aa1n02x4               g014(.a(new_n106), .b(new_n108), .c(new_n109), .d(new_n107), .out0(new_n110));
  inv000aa1d42x5               g015(.a(\a[3] ), .o1(new_n111));
  inv000aa1d42x5               g016(.a(\b[2] ), .o1(new_n112));
  aoai13aa1n03x5               g017(.a(new_n107), .b(new_n106), .c(new_n111), .d(new_n112), .o1(new_n113));
  aobi12aa1n03x7               g018(.a(new_n113), .b(new_n110), .c(new_n105), .out0(new_n114));
  nand22aa1n04x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor022aa1n16x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor002aa1n06x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nano23aa1n02x4               g023(.a(new_n117), .b(new_n116), .c(new_n118), .d(new_n115), .out0(new_n119));
  nand22aa1n03x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  orn002aa1n03x5               g025(.a(\a[8] ), .b(\b[7] ), .o(new_n121));
  nand42aa1n02x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  xnrc02aa1n12x5               g027(.a(\b[6] ), .b(\a[7] ), .out0(new_n123));
  nona22aa1n02x4               g028(.a(new_n119), .b(new_n123), .c(new_n122), .out0(new_n124));
  nona22aa1n02x4               g029(.a(new_n120), .b(\b[6] ), .c(\a[7] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n120), .b(new_n116), .c(new_n117), .d(new_n115), .o1(new_n126));
  nor002aa1n02x5               g031(.a(new_n126), .b(new_n123), .o1(new_n127));
  nano22aa1n03x7               g032(.a(new_n127), .b(new_n121), .c(new_n125), .out0(new_n128));
  oai012aa1n02x7               g033(.a(new_n128), .b(new_n114), .c(new_n124), .o1(new_n129));
  nanp02aa1n09x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n100), .b(new_n101), .c(new_n129), .d(new_n130), .o1(new_n131));
  tech160nm_fioaoi03aa1n04x5   g036(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n132));
  nona23aa1n03x5               g037(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n133));
  oai012aa1n04x7               g038(.a(new_n113), .b(new_n133), .c(new_n132), .o1(new_n134));
  nona23aa1n03x5               g039(.a(new_n115), .b(new_n118), .c(new_n117), .d(new_n116), .out0(new_n135));
  nor043aa1n03x5               g040(.a(new_n135), .b(new_n122), .c(new_n123), .o1(new_n136));
  oai112aa1n04x5               g041(.a(new_n121), .b(new_n125), .c(new_n126), .d(new_n123), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n130), .b(new_n101), .out0(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n137), .c(new_n134), .d(new_n136), .o1(new_n139));
  nona22aa1n02x4               g044(.a(new_n139), .b(new_n101), .c(new_n100), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n131), .b(new_n140), .o1(\s[10] ));
  xorc02aa1n12x5               g046(.a(\a[11] ), .b(\b[10] ), .out0(new_n142));
  xobna2aa1n03x5               g047(.a(new_n142), .b(new_n140), .c(new_n98), .out0(\s[11] ));
  orn002aa1n02x5               g048(.a(\a[11] ), .b(\b[10] ), .o(new_n144));
  nanp03aa1n02x5               g049(.a(new_n140), .b(new_n98), .c(new_n142), .o1(new_n145));
  xorc02aa1n12x5               g050(.a(\a[12] ), .b(\b[11] ), .out0(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n145), .c(new_n144), .out0(\s[12] ));
  nanp02aa1n03x5               g052(.a(new_n134), .b(new_n136), .o1(new_n148));
  nano23aa1n03x7               g053(.a(new_n97), .b(new_n101), .c(new_n130), .d(new_n98), .out0(new_n149));
  nand23aa1n03x5               g054(.a(new_n149), .b(new_n142), .c(new_n146), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\a[12] ), .o1(new_n151));
  inv000aa1d42x5               g056(.a(\b[11] ), .o1(new_n152));
  tech160nm_fioai012aa1n05x5   g057(.a(new_n98), .b(new_n101), .c(new_n97), .o1(new_n153));
  nanp02aa1n03x5               g058(.a(new_n153), .b(new_n144), .o1(new_n154));
  aoi022aa1n02x5               g059(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n155));
  aoi022aa1n02x5               g060(.a(new_n154), .b(new_n155), .c(new_n152), .d(new_n151), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n150), .c(new_n148), .d(new_n128), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand02aa1n08x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand22aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nona23aa1n09x5               g069(.a(new_n164), .b(new_n160), .c(new_n159), .d(new_n163), .out0(new_n165));
  inv040aa1n03x5               g070(.a(new_n165), .o1(new_n166));
  ao0012aa1n12x5               g071(.a(new_n163), .b(new_n159), .c(new_n164), .o(new_n167));
  nor022aa1n16x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n16x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nanb02aa1n12x5               g074(.a(new_n168), .b(new_n169), .out0(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  aoai13aa1n06x5               g076(.a(new_n171), .b(new_n167), .c(new_n157), .d(new_n166), .o1(new_n172));
  aoi112aa1n02x5               g077(.a(new_n171), .b(new_n167), .c(new_n157), .d(new_n166), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(\s[15] ));
  nor002aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand02aa1n03x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  oaoi13aa1n02x5               g082(.a(new_n177), .b(new_n172), .c(\a[15] ), .d(\b[14] ), .o1(new_n178));
  oai112aa1n02x5               g083(.a(new_n172), .b(new_n177), .c(\b[14] ), .d(\a[15] ), .o1(new_n179));
  norb02aa1n02x7               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  nano23aa1n06x5               g085(.a(new_n168), .b(new_n175), .c(new_n176), .d(new_n169), .out0(new_n181));
  nano22aa1n12x5               g086(.a(new_n150), .b(new_n166), .c(new_n181), .out0(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n137), .c(new_n134), .d(new_n136), .o1(new_n183));
  nanp02aa1n03x5               g088(.a(new_n154), .b(new_n155), .o1(new_n184));
  oaib12aa1n02x5               g089(.a(new_n184), .b(\b[11] ), .c(new_n151), .out0(new_n185));
  nor003aa1n03x5               g090(.a(new_n165), .b(new_n170), .c(new_n177), .o1(new_n186));
  aoi112aa1n02x5               g091(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n187));
  nand42aa1n02x5               g092(.a(new_n181), .b(new_n167), .o1(new_n188));
  nona22aa1n02x4               g093(.a(new_n188), .b(new_n187), .c(new_n175), .out0(new_n189));
  aoi012aa1n12x5               g094(.a(new_n189), .b(new_n185), .c(new_n186), .o1(new_n190));
  nand02aa1d06x5               g095(.a(new_n183), .b(new_n190), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g097(.a(\a[18] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  oaoi03aa1n03x5               g100(.a(new_n194), .b(new_n195), .c(new_n191), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  xroi22aa1d06x4               g102(.a(new_n194), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n198));
  nor042aa1n04x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  aoi112aa1n09x5               g104(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n200));
  nor042aa1n06x5               g105(.a(new_n200), .b(new_n199), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  nor002aa1n12x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nanp02aa1n09x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  norb02aa1n12x5               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n202), .c(new_n191), .d(new_n198), .o1(new_n206));
  aoi112aa1n02x5               g111(.a(new_n205), .b(new_n202), .c(new_n191), .d(new_n198), .o1(new_n207));
  norb02aa1n02x7               g112(.a(new_n206), .b(new_n207), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nand02aa1d28x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  norb02aa1n15x5               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  oaoi13aa1n06x5               g118(.a(new_n213), .b(new_n206), .c(\a[19] ), .d(\b[18] ), .o1(new_n214));
  nona22aa1n02x5               g119(.a(new_n206), .b(new_n212), .c(new_n203), .out0(new_n215));
  norb02aa1n03x4               g120(.a(new_n215), .b(new_n214), .out0(\s[20] ));
  nona23aa1n09x5               g121(.a(new_n211), .b(new_n204), .c(new_n203), .d(new_n210), .out0(new_n217));
  inv040aa1n02x5               g122(.a(new_n217), .o1(new_n218));
  nanp02aa1n02x5               g123(.a(new_n198), .b(new_n218), .o1(new_n219));
  oaih12aa1n06x5               g124(.a(new_n211), .b(new_n210), .c(new_n203), .o1(new_n220));
  oai012aa1n18x5               g125(.a(new_n220), .b(new_n217), .c(new_n201), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n222), .b(new_n219), .c(new_n183), .d(new_n190), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xorc02aa1n12x5               g130(.a(\a[21] ), .b(\b[20] ), .out0(new_n226));
  xorc02aa1n12x5               g131(.a(\a[22] ), .b(\b[21] ), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n225), .c(new_n223), .d(new_n226), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n225), .b(new_n227), .c(new_n223), .d(new_n226), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n228), .b(new_n229), .out0(\s[22] ));
  nand22aa1n12x5               g135(.a(new_n227), .b(new_n226), .o1(new_n231));
  nanb03aa1n06x5               g136(.a(new_n231), .b(new_n198), .c(new_n218), .out0(new_n232));
  oai112aa1n06x5               g137(.a(new_n205), .b(new_n212), .c(new_n200), .d(new_n199), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\a[22] ), .o1(new_n234));
  inv040aa1d32x5               g139(.a(\b[21] ), .o1(new_n235));
  oao003aa1n03x5               g140(.a(new_n234), .b(new_n235), .c(new_n225), .carry(new_n236));
  inv030aa1n02x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n12x5               g142(.a(new_n237), .b(new_n231), .c(new_n233), .d(new_n220), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  aoai13aa1n04x5               g144(.a(new_n239), .b(new_n232), .c(new_n183), .d(new_n190), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  xorc02aa1n02x5               g147(.a(\a[23] ), .b(\b[22] ), .out0(new_n243));
  xorc02aa1n02x5               g148(.a(\a[24] ), .b(\b[23] ), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n242), .c(new_n240), .d(new_n243), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n242), .b(new_n244), .c(new_n240), .d(new_n243), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n245), .b(new_n246), .out0(\s[24] ));
  and002aa1n06x5               g152(.a(new_n244), .b(new_n243), .o(new_n248));
  nona23aa1n02x4               g153(.a(new_n248), .b(new_n198), .c(new_n231), .d(new_n217), .out0(new_n249));
  inv000aa1d42x5               g154(.a(\a[24] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[23] ), .o1(new_n251));
  oao003aa1n02x5               g156(.a(new_n250), .b(new_n251), .c(new_n242), .carry(new_n252));
  tech160nm_fiaoi012aa1n05x5   g157(.a(new_n252), .b(new_n238), .c(new_n248), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n249), .c(new_n183), .d(new_n190), .o1(new_n254));
  xorb03aa1n02x5               g159(.a(new_n254), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g160(.a(\b[24] ), .b(\a[25] ), .o1(new_n256));
  tech160nm_fixorc02aa1n05x5   g161(.a(\a[25] ), .b(\b[24] ), .out0(new_n257));
  xorc02aa1n12x5               g162(.a(\a[26] ), .b(\b[25] ), .out0(new_n258));
  aoai13aa1n04x5               g163(.a(new_n258), .b(new_n256), .c(new_n254), .d(new_n257), .o1(new_n259));
  aoi112aa1n02x7               g164(.a(new_n256), .b(new_n258), .c(new_n254), .d(new_n257), .o1(new_n260));
  norb02aa1n03x4               g165(.a(new_n259), .b(new_n260), .out0(\s[26] ));
  aoi112aa1n02x5               g166(.a(new_n187), .b(new_n175), .c(new_n181), .d(new_n167), .o1(new_n262));
  oaib12aa1n02x5               g167(.a(new_n262), .b(new_n156), .c(new_n186), .out0(new_n263));
  and002aa1n09x5               g168(.a(new_n258), .b(new_n257), .o(new_n264));
  nano22aa1n03x7               g169(.a(new_n232), .b(new_n248), .c(new_n264), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n263), .c(new_n129), .d(new_n182), .o1(new_n266));
  aoai13aa1n09x5               g171(.a(new_n264), .b(new_n252), .c(new_n238), .d(new_n248), .o1(new_n267));
  oai022aa1n02x5               g172(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n268));
  aob012aa1n02x5               g173(.a(new_n268), .b(\b[25] ), .c(\a[26] ), .out0(new_n269));
  xorc02aa1n12x5               g174(.a(\a[27] ), .b(\b[26] ), .out0(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  aoi013aa1n03x5               g176(.a(new_n271), .b(new_n266), .c(new_n267), .d(new_n269), .o1(new_n272));
  inv020aa1n02x5               g177(.a(new_n265), .o1(new_n273));
  aoi012aa1n06x5               g178(.a(new_n273), .b(new_n183), .c(new_n190), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n231), .o1(new_n275));
  aoai13aa1n06x5               g180(.a(new_n248), .b(new_n236), .c(new_n221), .d(new_n275), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n252), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n264), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n269), .b(new_n278), .c(new_n276), .d(new_n277), .o1(new_n279));
  norp03aa1n02x5               g184(.a(new_n279), .b(new_n274), .c(new_n270), .o1(new_n280));
  nor002aa1n02x5               g185(.a(new_n272), .b(new_n280), .o1(\s[27] ));
  norp02aa1n02x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  inv040aa1n03x5               g187(.a(new_n282), .o1(new_n283));
  oaih12aa1n02x5               g188(.a(new_n270), .b(new_n279), .c(new_n274), .o1(new_n284));
  xnrc02aa1n12x5               g189(.a(\b[27] ), .b(\a[28] ), .out0(new_n285));
  tech160nm_fiaoi012aa1n02p5x5 g190(.a(new_n285), .b(new_n284), .c(new_n283), .o1(new_n286));
  nano22aa1n03x5               g191(.a(new_n272), .b(new_n283), .c(new_n285), .out0(new_n287));
  norp02aa1n03x5               g192(.a(new_n286), .b(new_n287), .o1(\s[28] ));
  norb02aa1n02x5               g193(.a(new_n270), .b(new_n285), .out0(new_n289));
  oaih12aa1n02x5               g194(.a(new_n289), .b(new_n279), .c(new_n274), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n283), .carry(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[28] ), .b(\a[29] ), .out0(new_n292));
  aoi012aa1n02x5               g197(.a(new_n292), .b(new_n290), .c(new_n291), .o1(new_n293));
  inv000aa1n02x5               g198(.a(new_n289), .o1(new_n294));
  aoi013aa1n02x5               g199(.a(new_n294), .b(new_n266), .c(new_n267), .d(new_n269), .o1(new_n295));
  nano22aa1n03x5               g200(.a(new_n295), .b(new_n291), .c(new_n292), .out0(new_n296));
  norp02aa1n03x5               g201(.a(new_n293), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g202(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g203(.a(new_n270), .b(new_n292), .c(new_n285), .out0(new_n299));
  tech160nm_fioai012aa1n03p5x5 g204(.a(new_n299), .b(new_n279), .c(new_n274), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .carry(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[29] ), .b(\a[30] ), .out0(new_n302));
  tech160nm_fiaoi012aa1n03p5x5 g207(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n299), .o1(new_n304));
  aoi013aa1n02x5               g209(.a(new_n304), .b(new_n266), .c(new_n267), .d(new_n269), .o1(new_n305));
  nano22aa1n03x5               g210(.a(new_n305), .b(new_n301), .c(new_n302), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n303), .b(new_n306), .o1(\s[30] ));
  norb02aa1n02x5               g212(.a(new_n299), .b(new_n302), .out0(new_n308));
  oaih12aa1n02x5               g213(.a(new_n308), .b(new_n279), .c(new_n274), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n301), .carry(new_n310));
  xnrc02aa1n02x5               g215(.a(\b[30] ), .b(\a[31] ), .out0(new_n311));
  aoi012aa1n02x5               g216(.a(new_n311), .b(new_n309), .c(new_n310), .o1(new_n312));
  inv000aa1n02x5               g217(.a(new_n308), .o1(new_n313));
  aoi013aa1n02x5               g218(.a(new_n313), .b(new_n266), .c(new_n267), .d(new_n269), .o1(new_n314));
  nano22aa1n03x5               g219(.a(new_n314), .b(new_n310), .c(new_n311), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n312), .b(new_n315), .o1(\s[31] ));
  xorb03aa1n02x5               g221(.a(new_n132), .b(\b[2] ), .c(new_n111), .out0(\s[3] ));
  nanb03aa1n02x5               g222(.a(new_n108), .b(new_n105), .c(new_n109), .out0(new_n318));
  aboi22aa1n03x5               g223(.a(new_n106), .b(new_n107), .c(new_n111), .d(new_n112), .out0(new_n319));
  aboi22aa1n03x5               g224(.a(new_n106), .b(new_n134), .c(new_n318), .d(new_n319), .out0(\s[4] ));
  xorb03aa1n02x5               g225(.a(new_n134), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g226(.a(\a[5] ), .b(\b[4] ), .c(new_n114), .o1(new_n322));
  xorb03aa1n02x5               g227(.a(new_n322), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g228(.a(\a[7] ), .o1(new_n324));
  oai012aa1n02x5               g229(.a(new_n115), .b(new_n322), .c(new_n116), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[6] ), .c(new_n324), .out0(\s[7] ));
  oaoi03aa1n02x5               g231(.a(\a[7] ), .b(\b[6] ), .c(new_n325), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g233(.a(new_n138), .b(new_n148), .c(new_n128), .out0(\s[9] ));
endmodule


