// Benchmark "adder" written by ABC on Thu Jul 18 07:23:26 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n308, new_n309, new_n310,
    new_n311, new_n314, new_n315, new_n316, new_n318, new_n319, new_n321,
    new_n322, new_n323, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d28x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand42aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nor022aa1n04x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nor002aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  oai012aa1n02x5               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  inv000aa1d42x5               g008(.a(\a[2] ), .o1(new_n104));
  inv000aa1d42x5               g009(.a(\b[1] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  oaoi03aa1n02x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nona23aa1n03x5               g013(.a(new_n100), .b(new_n108), .c(new_n102), .d(new_n101), .out0(new_n109));
  oai012aa1n02x7               g014(.a(new_n103), .b(new_n109), .c(new_n107), .o1(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .out0(new_n111));
  tech160nm_finor002aa1n05x5   g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nona23aa1n02x4               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .out0(new_n117));
  nor003aa1n02x5               g022(.a(new_n116), .b(new_n117), .c(new_n111), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(new_n110), .b(new_n118), .o1(new_n119));
  orn002aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .o(new_n120));
  inv000aa1n03x5               g025(.a(new_n112), .o1(new_n121));
  oai022aa1n06x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  aob012aa1n06x5               g027(.a(new_n122), .b(\b[5] ), .c(\a[6] ), .out0(new_n123));
  aob012aa1n02x5               g028(.a(new_n113), .b(\b[7] ), .c(\a[8] ), .out0(new_n124));
  aoai13aa1n09x5               g029(.a(new_n120), .b(new_n124), .c(new_n123), .d(new_n121), .o1(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  aoai13aa1n02x5               g033(.a(new_n99), .b(new_n128), .c(new_n119), .d(new_n126), .o1(new_n129));
  xorb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1d32x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nand42aa1d28x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nanb02aa1n06x5               g037(.a(new_n131), .b(new_n132), .out0(new_n133));
  inv040aa1d30x5               g038(.a(new_n133), .o1(new_n134));
  aoai13aa1n12x5               g039(.a(new_n132), .b(new_n131), .c(new_n97), .d(new_n98), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nor042aa1n09x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nanp02aa1n04x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n136), .c(new_n129), .d(new_n134), .o1(new_n140));
  aoi112aa1n02x5               g045(.a(new_n139), .b(new_n136), .c(new_n129), .d(new_n134), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n140), .b(new_n141), .out0(\s[11] ));
  inv000aa1d42x5               g047(.a(new_n137), .o1(new_n143));
  nor042aa1n09x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanp02aa1n04x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nanb02aa1n02x5               g050(.a(new_n144), .b(new_n145), .out0(new_n146));
  nanp03aa1n02x5               g051(.a(new_n140), .b(new_n143), .c(new_n146), .o1(new_n147));
  aoi012aa1n02x5               g052(.a(new_n146), .b(new_n140), .c(new_n143), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n147), .b(new_n148), .out0(\s[12] ));
  nona23aa1n09x5               g054(.a(new_n145), .b(new_n138), .c(new_n137), .d(new_n144), .out0(new_n150));
  norb03aa1n02x5               g055(.a(new_n127), .b(new_n150), .c(new_n133), .out0(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n125), .c(new_n110), .d(new_n118), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n144), .o1(new_n153));
  nand42aa1n03x5               g058(.a(new_n137), .b(new_n145), .o1(new_n154));
  oai112aa1n06x5               g059(.a(new_n154), .b(new_n153), .c(new_n150), .d(new_n135), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(new_n152), .b(new_n156), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n02x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nanp02aa1n02x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n02x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nona23aa1n02x4               g069(.a(new_n164), .b(new_n160), .c(new_n159), .d(new_n163), .out0(new_n165));
  oai012aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n159), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n165), .c(new_n152), .d(new_n156), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n169), .b(new_n167), .c(new_n170), .o1(new_n171));
  nor022aa1n12x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  nanp02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n171), .b(new_n174), .c(new_n173), .out0(\s[16] ));
  nano23aa1n02x4               g080(.a(new_n137), .b(new_n144), .c(new_n145), .d(new_n138), .out0(new_n176));
  nano23aa1n02x4               g081(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n177));
  nanb02aa1n02x5               g082(.a(new_n169), .b(new_n170), .out0(new_n178));
  nanb02aa1n02x5               g083(.a(new_n172), .b(new_n174), .out0(new_n179));
  nona22aa1n02x4               g084(.a(new_n177), .b(new_n178), .c(new_n179), .out0(new_n180));
  nano32aa1n02x4               g085(.a(new_n180), .b(new_n176), .c(new_n134), .d(new_n127), .out0(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n125), .c(new_n110), .d(new_n118), .o1(new_n182));
  norp03aa1n02x5               g087(.a(new_n165), .b(new_n178), .c(new_n179), .o1(new_n183));
  aoi112aa1n02x5               g088(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n184));
  oai013aa1n02x4               g089(.a(new_n173), .b(new_n166), .c(new_n178), .d(new_n179), .o1(new_n185));
  aoi112aa1n06x5               g090(.a(new_n185), .b(new_n184), .c(new_n155), .d(new_n183), .o1(new_n186));
  nand02aa1d10x5               g091(.a(new_n186), .b(new_n182), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g093(.a(\a[18] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(\a[17] ), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[16] ), .o1(new_n191));
  oaoi03aa1n02x5               g096(.a(new_n190), .b(new_n191), .c(new_n187), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[17] ), .c(new_n189), .out0(\s[18] ));
  xroi22aa1d06x4               g098(.a(new_n190), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n194));
  nanp02aa1n02x5               g099(.a(new_n191), .b(new_n190), .o1(new_n195));
  oaoi03aa1n02x5               g100(.a(\a[18] ), .b(\b[17] ), .c(new_n195), .o1(new_n196));
  nor042aa1n02x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanp02aa1n03x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  norb02aa1n02x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n196), .c(new_n187), .d(new_n194), .o1(new_n200));
  aoi112aa1n02x5               g105(.a(new_n199), .b(new_n196), .c(new_n187), .d(new_n194), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n200), .b(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n02x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand42aa1n06x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  norb02aa1n02x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  nona22aa1n03x5               g111(.a(new_n200), .b(new_n206), .c(new_n197), .out0(new_n207));
  inv000aa1n03x5               g112(.a(new_n206), .o1(new_n208));
  oaoi13aa1n04x5               g113(.a(new_n208), .b(new_n200), .c(\a[19] ), .d(\b[18] ), .o1(new_n209));
  norb02aa1n03x4               g114(.a(new_n207), .b(new_n209), .out0(\s[20] ));
  nona23aa1n12x5               g115(.a(new_n194), .b(new_n198), .c(new_n208), .d(new_n197), .out0(new_n211));
  oai022aa1n02x5               g116(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n212));
  oaib12aa1n02x5               g117(.a(new_n212), .b(new_n189), .c(\b[17] ), .out0(new_n213));
  tech160nm_fiao0012aa1n02p5x5 g118(.a(new_n204), .b(new_n197), .c(new_n205), .o(new_n214));
  nona23aa1n06x5               g119(.a(new_n205), .b(new_n198), .c(new_n197), .d(new_n204), .out0(new_n215));
  oabi12aa1n12x5               g120(.a(new_n214), .b(new_n215), .c(new_n213), .out0(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n03x5               g122(.a(new_n217), .b(new_n211), .c(new_n186), .d(new_n182), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  xorc02aa1n02x5               g125(.a(\a[21] ), .b(\b[20] ), .out0(new_n221));
  xorc02aa1n02x5               g126(.a(\a[22] ), .b(\b[21] ), .out0(new_n222));
  aoi112aa1n02x5               g127(.a(new_n220), .b(new_n222), .c(new_n218), .d(new_n221), .o1(new_n223));
  aoai13aa1n03x5               g128(.a(new_n222), .b(new_n220), .c(new_n218), .d(new_n221), .o1(new_n224));
  norb02aa1n03x4               g129(.a(new_n224), .b(new_n223), .out0(\s[22] ));
  inv000aa1d42x5               g130(.a(\a[21] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  nanb02aa1n03x5               g133(.a(new_n211), .b(new_n228), .out0(new_n229));
  inv000aa1d42x5               g134(.a(\b[21] ), .o1(new_n230));
  tech160nm_fioaoi03aa1n03p5x5 g135(.a(new_n227), .b(new_n230), .c(new_n220), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n216), .c(new_n228), .o1(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n229), .c(new_n186), .d(new_n182), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  xorc02aa1n02x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  xorc02aa1n02x5               g142(.a(\a[24] ), .b(\b[23] ), .out0(new_n238));
  aoi112aa1n03x5               g143(.a(new_n236), .b(new_n238), .c(new_n234), .d(new_n237), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n238), .b(new_n236), .c(new_n234), .d(new_n237), .o1(new_n240));
  norb02aa1n03x4               g145(.a(new_n240), .b(new_n239), .out0(\s[24] ));
  nanp02aa1n03x5               g146(.a(new_n238), .b(new_n237), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  nano22aa1n03x7               g148(.a(new_n211), .b(new_n228), .c(new_n243), .out0(new_n244));
  nano23aa1n02x4               g149(.a(new_n197), .b(new_n204), .c(new_n205), .d(new_n198), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n228), .b(new_n214), .c(new_n245), .d(new_n196), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n247));
  oab012aa1n02x4               g152(.a(new_n247), .b(\a[24] ), .c(\b[23] ), .out0(new_n248));
  aoai13aa1n04x5               g153(.a(new_n248), .b(new_n242), .c(new_n246), .d(new_n231), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[25] ), .b(\b[24] ), .out0(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n249), .c(new_n187), .d(new_n244), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(new_n250), .b(new_n249), .c(new_n187), .d(new_n244), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n251), .b(new_n252), .out0(\s[25] ));
  norp02aa1n02x5               g158(.a(\b[24] ), .b(\a[25] ), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[26] ), .b(\b[25] ), .out0(new_n255));
  nona22aa1n03x5               g160(.a(new_n251), .b(new_n255), .c(new_n254), .out0(new_n256));
  inv000aa1n02x5               g161(.a(new_n254), .o1(new_n257));
  aobi12aa1n03x5               g162(.a(new_n255), .b(new_n251), .c(new_n257), .out0(new_n258));
  norb02aa1n03x4               g163(.a(new_n256), .b(new_n258), .out0(\s[26] ));
  and002aa1n02x5               g164(.a(new_n255), .b(new_n250), .o(new_n260));
  nano32aa1d12x5               g165(.a(new_n211), .b(new_n260), .c(new_n228), .d(new_n243), .out0(new_n261));
  nand02aa1d08x5               g166(.a(new_n187), .b(new_n261), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[26] ), .b(\b[25] ), .c(new_n257), .carry(new_n263));
  aobi12aa1n12x5               g168(.a(new_n263), .b(new_n249), .c(new_n260), .out0(new_n264));
  xorc02aa1n02x5               g169(.a(\a[27] ), .b(\b[26] ), .out0(new_n265));
  xnbna2aa1n03x5               g170(.a(new_n265), .b(new_n262), .c(new_n264), .out0(\s[27] ));
  norp02aa1n02x5               g171(.a(\b[26] ), .b(\a[27] ), .o1(new_n267));
  inv040aa1n03x5               g172(.a(new_n267), .o1(new_n268));
  aobi12aa1n02x7               g173(.a(new_n265), .b(new_n262), .c(new_n264), .out0(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[27] ), .b(\a[28] ), .out0(new_n270));
  nano22aa1n03x5               g175(.a(new_n269), .b(new_n268), .c(new_n270), .out0(new_n271));
  inv000aa1d42x5               g176(.a(new_n211), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n228), .o1(new_n273));
  inv000aa1n02x5               g178(.a(new_n260), .o1(new_n274));
  nona32aa1n02x4               g179(.a(new_n272), .b(new_n274), .c(new_n242), .d(new_n273), .out0(new_n275));
  tech160nm_fiaoi012aa1n05x5   g180(.a(new_n275), .b(new_n186), .c(new_n182), .o1(new_n276));
  aoai13aa1n02x7               g181(.a(new_n243), .b(new_n232), .c(new_n216), .d(new_n228), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n263), .b(new_n274), .c(new_n277), .d(new_n248), .o1(new_n278));
  oai012aa1n02x5               g183(.a(new_n265), .b(new_n278), .c(new_n276), .o1(new_n279));
  aoi012aa1n03x5               g184(.a(new_n270), .b(new_n279), .c(new_n268), .o1(new_n280));
  norp02aa1n03x5               g185(.a(new_n280), .b(new_n271), .o1(\s[28] ));
  norb02aa1n02x5               g186(.a(new_n265), .b(new_n270), .out0(new_n282));
  oaih12aa1n02x5               g187(.a(new_n282), .b(new_n278), .c(new_n276), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .c(new_n268), .carry(new_n284));
  xnrc02aa1n02x5               g189(.a(\b[28] ), .b(\a[29] ), .out0(new_n285));
  tech160nm_fiaoi012aa1n02p5x5 g190(.a(new_n285), .b(new_n283), .c(new_n284), .o1(new_n286));
  aobi12aa1n06x5               g191(.a(new_n282), .b(new_n262), .c(new_n264), .out0(new_n287));
  nano22aa1n03x7               g192(.a(new_n287), .b(new_n284), .c(new_n285), .out0(new_n288));
  norp02aa1n03x5               g193(.a(new_n286), .b(new_n288), .o1(\s[29] ));
  xorb03aa1n02x5               g194(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g195(.a(new_n265), .b(new_n285), .c(new_n270), .out0(new_n291));
  oai012aa1n02x5               g196(.a(new_n291), .b(new_n278), .c(new_n276), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .carry(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[29] ), .b(\a[30] ), .out0(new_n294));
  aoi012aa1n03x5               g199(.a(new_n294), .b(new_n292), .c(new_n293), .o1(new_n295));
  aobi12aa1n03x5               g200(.a(new_n291), .b(new_n262), .c(new_n264), .out0(new_n296));
  nano22aa1n03x5               g201(.a(new_n296), .b(new_n293), .c(new_n294), .out0(new_n297));
  norp02aa1n03x5               g202(.a(new_n295), .b(new_n297), .o1(\s[30] ));
  xnrc02aa1n02x5               g203(.a(\b[30] ), .b(\a[31] ), .out0(new_n299));
  norb02aa1n02x5               g204(.a(new_n291), .b(new_n294), .out0(new_n300));
  oai012aa1n02x5               g205(.a(new_n300), .b(new_n278), .c(new_n276), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n302));
  aoi012aa1n03x5               g207(.a(new_n299), .b(new_n301), .c(new_n302), .o1(new_n303));
  aobi12aa1n06x5               g208(.a(new_n300), .b(new_n262), .c(new_n264), .out0(new_n304));
  nano22aa1n03x7               g209(.a(new_n304), .b(new_n299), .c(new_n302), .out0(new_n305));
  norp02aa1n03x5               g210(.a(new_n303), .b(new_n305), .o1(\s[31] ));
  xnrb03aa1n02x5               g211(.a(new_n107), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanb02aa1n02x5               g212(.a(new_n102), .b(new_n100), .out0(new_n308));
  norp02aa1n02x5               g213(.a(new_n109), .b(new_n107), .o1(new_n309));
  oao003aa1n02x5               g214(.a(new_n104), .b(new_n105), .c(new_n106), .carry(new_n310));
  oai112aa1n02x5               g215(.a(new_n108), .b(new_n308), .c(new_n310), .d(new_n101), .o1(new_n311));
  oai013aa1n02x4               g216(.a(new_n311), .b(new_n309), .c(new_n101), .d(new_n308), .o1(\s[4] ));
  xorb03aa1n02x5               g217(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nano23aa1n02x4               g218(.a(new_n102), .b(new_n101), .c(new_n108), .d(new_n100), .out0(new_n314));
  aobi12aa1n02x5               g219(.a(new_n103), .b(new_n314), .c(new_n310), .out0(new_n315));
  oaoi03aa1n02x5               g220(.a(\a[5] ), .b(\b[4] ), .c(new_n315), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g222(.a(new_n113), .b(new_n112), .out0(new_n318));
  nanb02aa1n02x5               g223(.a(new_n117), .b(new_n316), .out0(new_n319));
  xnbna2aa1n03x5               g224(.a(new_n318), .b(new_n319), .c(new_n123), .out0(\s[7] ));
  norb02aa1n02x5               g225(.a(new_n316), .b(new_n117), .out0(new_n321));
  oaib12aa1n02x5               g226(.a(new_n318), .b(new_n321), .c(new_n123), .out0(new_n322));
  aoi012aa1n02x5               g227(.a(new_n111), .b(new_n322), .c(new_n121), .o1(new_n323));
  nanp03aa1n02x5               g228(.a(new_n322), .b(new_n111), .c(new_n121), .o1(new_n324));
  norb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(\s[8] ));
  xnbna2aa1n03x5               g230(.a(new_n127), .b(new_n119), .c(new_n126), .out0(\s[9] ));
endmodule


