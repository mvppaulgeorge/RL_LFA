// Benchmark "adder" written by ABC on Wed Jul 17 14:46:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n148, new_n149,
    new_n150, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n316, new_n319,
    new_n321, new_n322, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d32x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d28x5               g002(.a(\b[8] ), .o1(new_n98));
  and002aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n12x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  xorc02aa1n12x5               g005(.a(\a[4] ), .b(\b[3] ), .out0(new_n101));
  nor042aa1n02x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  norb02aa1n06x5               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  nanp03aa1d12x5               g009(.a(new_n100), .b(new_n101), .c(new_n104), .o1(new_n105));
  orn002aa1n06x5               g010(.a(\a[3] ), .b(\b[2] ), .o(new_n106));
  oao003aa1n03x5               g011(.a(\a[4] ), .b(\b[3] ), .c(new_n106), .carry(new_n107));
  nand42aa1d28x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nor042aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor002aa1n06x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n24x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nano23aa1n09x5               g016(.a(new_n110), .b(new_n109), .c(new_n111), .d(new_n108), .out0(new_n112));
  tech160nm_fixorc02aa1n05x5   g017(.a(\a[6] ), .b(\b[5] ), .out0(new_n113));
  xorc02aa1n12x5               g018(.a(\a[5] ), .b(\b[4] ), .out0(new_n114));
  nand03aa1n02x5               g019(.a(new_n112), .b(new_n113), .c(new_n114), .o1(new_n115));
  nor042aa1d18x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  inv030aa1n04x5               g021(.a(new_n116), .o1(new_n117));
  oaoi03aa1n03x5               g022(.a(\a[6] ), .b(\b[5] ), .c(new_n117), .o1(new_n118));
  oai022aa1n02x5               g023(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n119));
  aoi022aa1n06x5               g024(.a(new_n112), .b(new_n118), .c(new_n108), .d(new_n119), .o1(new_n120));
  aoai13aa1n12x5               g025(.a(new_n120), .b(new_n115), .c(new_n105), .d(new_n107), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(new_n97), .b(new_n98), .c(new_n121), .o1(new_n122));
  xnrb03aa1n03x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1d18x5               g028(.a(\b[9] ), .b(\a[10] ), .o1(new_n124));
  nand02aa1n04x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nanb02aa1n03x5               g030(.a(new_n124), .b(new_n125), .out0(new_n126));
  xnrc02aa1n06x5               g031(.a(\b[8] ), .b(\a[9] ), .out0(new_n127));
  norp02aa1n02x5               g032(.a(new_n127), .b(new_n126), .o1(new_n128));
  aoai13aa1n06x5               g033(.a(new_n125), .b(new_n124), .c(new_n97), .d(new_n98), .o1(new_n129));
  aob012aa1n03x5               g034(.a(new_n129), .b(new_n121), .c(new_n128), .out0(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand42aa1d28x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  tech160nm_fiaoi012aa1n05x5   g038(.a(new_n132), .b(new_n130), .c(new_n133), .o1(new_n134));
  xnrb03aa1n03x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1d32x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand42aa1d28x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nano23aa1n09x5               g042(.a(new_n132), .b(new_n136), .c(new_n137), .d(new_n133), .out0(new_n138));
  nona22aa1n09x5               g043(.a(new_n138), .b(new_n127), .c(new_n126), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  nand22aa1n03x5               g045(.a(new_n121), .b(new_n140), .o1(new_n141));
  nona23aa1n09x5               g046(.a(new_n137), .b(new_n133), .c(new_n132), .d(new_n136), .out0(new_n142));
  ao0012aa1n03x7               g047(.a(new_n136), .b(new_n132), .c(new_n137), .o(new_n143));
  oabi12aa1n18x5               g048(.a(new_n143), .b(new_n142), .c(new_n129), .out0(new_n144));
  inv000aa1d42x5               g049(.a(new_n144), .o1(new_n145));
  nanp02aa1n06x5               g050(.a(new_n141), .b(new_n145), .o1(new_n146));
  xorb03aa1n02x5               g051(.a(new_n146), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  nand42aa1d28x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  aoi012aa1n06x5               g054(.a(new_n148), .b(new_n146), .c(new_n149), .o1(new_n150));
  xnrb03aa1n03x5               g055(.a(new_n150), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n09x5               g056(.a(\b[13] ), .b(\a[14] ), .o1(new_n152));
  nand42aa1d28x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nano23aa1d15x5               g058(.a(new_n148), .b(new_n152), .c(new_n153), .d(new_n149), .out0(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n144), .c(new_n121), .d(new_n140), .o1(new_n155));
  oai012aa1d24x5               g060(.a(new_n153), .b(new_n152), .c(new_n148), .o1(new_n156));
  nor042aa1n06x5               g061(.a(\b[14] ), .b(\a[15] ), .o1(new_n157));
  nanp02aa1n04x5               g062(.a(\b[14] ), .b(\a[15] ), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n157), .b(new_n158), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n155), .c(new_n156), .out0(\s[15] ));
  nand22aa1n03x5               g066(.a(new_n155), .b(new_n156), .o1(new_n162));
  nor042aa1n04x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nand02aa1n08x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  aoai13aa1n03x5               g070(.a(new_n165), .b(new_n157), .c(new_n162), .d(new_n160), .o1(new_n166));
  aoi112aa1n03x4               g071(.a(new_n157), .b(new_n165), .c(new_n162), .d(new_n158), .o1(new_n167));
  nanb02aa1n03x5               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  inv000aa1d42x5               g073(.a(\a[17] ), .o1(new_n169));
  nano23aa1n06x5               g074(.a(new_n157), .b(new_n163), .c(new_n164), .d(new_n158), .out0(new_n170));
  nano22aa1n12x5               g075(.a(new_n139), .b(new_n154), .c(new_n170), .out0(new_n171));
  inv000aa1n02x5               g076(.a(new_n170), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(new_n98), .b(new_n97), .o1(new_n173));
  tech160nm_fioaoi03aa1n03p5x5 g078(.a(\a[10] ), .b(\b[9] ), .c(new_n173), .o1(new_n174));
  aoai13aa1n03x5               g079(.a(new_n154), .b(new_n143), .c(new_n138), .d(new_n174), .o1(new_n175));
  tech160nm_fiaoi012aa1n04x5   g080(.a(new_n172), .b(new_n175), .c(new_n156), .o1(new_n176));
  aoi012aa1d24x5               g081(.a(new_n163), .b(new_n157), .c(new_n164), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  aoi112aa1n09x5               g083(.a(new_n176), .b(new_n178), .c(new_n121), .d(new_n171), .o1(new_n179));
  xorb03aa1n03x5               g084(.a(new_n179), .b(\b[16] ), .c(new_n169), .out0(\s[17] ));
  nanb02aa1n02x5               g085(.a(\b[16] ), .b(new_n169), .out0(new_n181));
  aoai13aa1n02x7               g086(.a(new_n177), .b(new_n172), .c(new_n175), .d(new_n156), .o1(new_n182));
  xorc02aa1n12x5               g087(.a(\a[17] ), .b(\b[16] ), .out0(new_n183));
  aoai13aa1n03x5               g088(.a(new_n183), .b(new_n182), .c(new_n121), .d(new_n171), .o1(new_n184));
  tech160nm_fixnrc02aa1n04x5   g089(.a(\b[17] ), .b(\a[18] ), .out0(new_n185));
  xobna2aa1n03x5               g090(.a(new_n185), .b(new_n184), .c(new_n181), .out0(\s[18] ));
  inv000aa1d42x5               g091(.a(\a[18] ), .o1(new_n187));
  xroi22aa1d06x4               g092(.a(new_n169), .b(\b[16] ), .c(new_n187), .d(\b[17] ), .out0(new_n188));
  inv000aa1n02x5               g093(.a(new_n188), .o1(new_n189));
  oaih22aa1d12x5               g094(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n190));
  oaib12aa1n18x5               g095(.a(new_n190), .b(new_n187), .c(\b[17] ), .out0(new_n191));
  tech160nm_fioai012aa1n05x5   g096(.a(new_n191), .b(new_n179), .c(new_n189), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g098(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand42aa1d28x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nanb02aa1d36x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  nor002aa1d32x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand42aa1d28x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nanb02aa1n12x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  aoai13aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n192), .d(new_n198), .o1(new_n202));
  nanp02aa1n06x5               g107(.a(new_n121), .b(new_n171), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n156), .o1(new_n204));
  aoai13aa1n04x5               g109(.a(new_n170), .b(new_n204), .c(new_n144), .d(new_n154), .o1(new_n205));
  nand23aa1n06x5               g110(.a(new_n203), .b(new_n205), .c(new_n177), .o1(new_n206));
  tech160nm_fioaoi03aa1n02p5x5 g111(.a(\a[18] ), .b(\b[17] ), .c(new_n181), .o1(new_n207));
  aoai13aa1n02x5               g112(.a(new_n198), .b(new_n207), .c(new_n206), .d(new_n188), .o1(new_n208));
  nona22aa1n02x4               g113(.a(new_n208), .b(new_n201), .c(new_n195), .out0(new_n209));
  nanp02aa1n03x5               g114(.a(new_n202), .b(new_n209), .o1(\s[20] ));
  nano23aa1d15x5               g115(.a(new_n195), .b(new_n199), .c(new_n200), .d(new_n196), .out0(new_n211));
  nanb03aa1d18x5               g116(.a(new_n185), .b(new_n211), .c(new_n183), .out0(new_n212));
  aoi012aa1n06x5               g117(.a(new_n199), .b(new_n195), .c(new_n200), .o1(new_n213));
  oai013aa1d12x5               g118(.a(new_n213), .b(new_n191), .c(new_n197), .d(new_n201), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  tech160nm_fioai012aa1n05x5   g120(.a(new_n215), .b(new_n179), .c(new_n212), .o1(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n04x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  xnrc02aa1n12x5               g125(.a(\b[21] ), .b(\a[22] ), .out0(new_n221));
  aoai13aa1n03x5               g126(.a(new_n221), .b(new_n218), .c(new_n216), .d(new_n220), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n212), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n220), .b(new_n214), .c(new_n206), .d(new_n223), .o1(new_n224));
  nona22aa1n02x4               g129(.a(new_n224), .b(new_n221), .c(new_n218), .out0(new_n225));
  nanp02aa1n03x5               g130(.a(new_n222), .b(new_n225), .o1(\s[22] ));
  nor042aa1n06x5               g131(.a(new_n221), .b(new_n219), .o1(new_n227));
  nano22aa1n03x7               g132(.a(new_n189), .b(new_n227), .c(new_n211), .out0(new_n228));
  inv000aa1n02x5               g133(.a(new_n228), .o1(new_n229));
  inv000aa1d42x5               g134(.a(\a[22] ), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\b[21] ), .o1(new_n231));
  oaoi03aa1n09x5               g136(.a(new_n230), .b(new_n231), .c(new_n218), .o1(new_n232));
  inv000aa1n02x5               g137(.a(new_n232), .o1(new_n233));
  aoi012aa1n09x5               g138(.a(new_n233), .b(new_n214), .c(new_n227), .o1(new_n234));
  tech160nm_fioai012aa1n05x5   g139(.a(new_n234), .b(new_n179), .c(new_n229), .o1(new_n235));
  xorb03aa1n02x5               g140(.a(new_n235), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g141(.a(\b[22] ), .b(\a[23] ), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  tech160nm_fixnrc02aa1n05x5   g143(.a(\b[23] ), .b(\a[24] ), .out0(new_n239));
  aoai13aa1n03x5               g144(.a(new_n239), .b(new_n237), .c(new_n235), .d(new_n238), .o1(new_n240));
  inv000aa1n02x5               g145(.a(new_n234), .o1(new_n241));
  aoai13aa1n02x5               g146(.a(new_n238), .b(new_n241), .c(new_n206), .d(new_n228), .o1(new_n242));
  nona22aa1n02x4               g147(.a(new_n242), .b(new_n239), .c(new_n237), .out0(new_n243));
  nanp02aa1n03x5               g148(.a(new_n240), .b(new_n243), .o1(\s[24] ));
  norb02aa1n03x4               g149(.a(new_n238), .b(new_n239), .out0(new_n245));
  inv030aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  nano32aa1n03x7               g151(.a(new_n246), .b(new_n188), .c(new_n227), .d(new_n211), .out0(new_n247));
  inv000aa1n02x5               g152(.a(new_n247), .o1(new_n248));
  inv000aa1n02x5               g153(.a(new_n213), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n227), .b(new_n249), .c(new_n211), .d(new_n207), .o1(new_n250));
  orn002aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .o(new_n251));
  oao003aa1n02x5               g156(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .carry(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n246), .c(new_n250), .d(new_n232), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  tech160nm_fioai012aa1n05x5   g159(.a(new_n254), .b(new_n179), .c(new_n248), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n03x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[25] ), .b(\a[26] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n260));
  aoai13aa1n02x5               g165(.a(new_n258), .b(new_n253), .c(new_n206), .d(new_n247), .o1(new_n261));
  nona22aa1n02x4               g166(.a(new_n261), .b(new_n259), .c(new_n257), .out0(new_n262));
  nanp02aa1n03x5               g167(.a(new_n260), .b(new_n262), .o1(\s[26] ));
  norb02aa1n06x5               g168(.a(new_n258), .b(new_n259), .out0(new_n264));
  nano23aa1n06x5               g169(.a(new_n212), .b(new_n246), .c(new_n264), .d(new_n227), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n182), .c(new_n121), .d(new_n171), .o1(new_n266));
  inv000aa1d42x5               g171(.a(\a[26] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(\b[25] ), .o1(new_n268));
  tech160nm_fioaoi03aa1n04x5   g173(.a(new_n267), .b(new_n268), .c(new_n257), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  aoi012aa1n06x5               g175(.a(new_n270), .b(new_n253), .c(new_n264), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[27] ), .b(\b[26] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n266), .c(new_n271), .out0(\s[27] ));
  inv000aa1n02x5               g178(.a(new_n265), .o1(new_n274));
  tech160nm_fioai012aa1n05x5   g179(.a(new_n271), .b(new_n179), .c(new_n274), .o1(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  nor002aa1n04x5               g181(.a(\b[27] ), .b(\a[28] ), .o1(new_n277));
  nand02aa1n06x5               g182(.a(\b[27] ), .b(\a[28] ), .o1(new_n278));
  nanb02aa1n06x5               g183(.a(new_n277), .b(new_n278), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n276), .c(new_n275), .d(new_n272), .o1(new_n280));
  aoai13aa1n02x5               g185(.a(new_n245), .b(new_n233), .c(new_n214), .d(new_n227), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n264), .o1(new_n282));
  aoai13aa1n04x5               g187(.a(new_n269), .b(new_n282), .c(new_n281), .d(new_n252), .o1(new_n283));
  aoai13aa1n02x5               g188(.a(new_n272), .b(new_n283), .c(new_n206), .d(new_n265), .o1(new_n284));
  nona22aa1n02x4               g189(.a(new_n284), .b(new_n279), .c(new_n276), .out0(new_n285));
  nanp02aa1n03x5               g190(.a(new_n280), .b(new_n285), .o1(\s[28] ));
  norb02aa1n03x5               g191(.a(new_n272), .b(new_n279), .out0(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n283), .c(new_n206), .d(new_n265), .o1(new_n288));
  nor002aa1n02x5               g193(.a(\b[28] ), .b(\a[29] ), .o1(new_n289));
  nand42aa1n08x5               g194(.a(\b[28] ), .b(\a[29] ), .o1(new_n290));
  norb02aa1n02x7               g195(.a(new_n290), .b(new_n289), .out0(new_n291));
  oai022aa1n02x5               g196(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n292));
  aboi22aa1n03x5               g197(.a(new_n289), .b(new_n290), .c(new_n292), .d(new_n278), .out0(new_n293));
  inv000aa1d42x5               g198(.a(new_n287), .o1(new_n294));
  oai012aa1n02x5               g199(.a(new_n278), .b(new_n277), .c(new_n276), .o1(new_n295));
  aoai13aa1n02x7               g200(.a(new_n295), .b(new_n294), .c(new_n266), .d(new_n271), .o1(new_n296));
  aoi022aa1n03x5               g201(.a(new_n296), .b(new_n291), .c(new_n288), .d(new_n293), .o1(\s[29] ));
  xnrb03aa1n02x5               g202(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g203(.a(new_n279), .b(new_n272), .c(new_n291), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n283), .c(new_n206), .d(new_n265), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  aoi113aa1n02x5               g206(.a(new_n301), .b(new_n289), .c(new_n290), .d(new_n292), .e(new_n278), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n299), .o1(new_n303));
  aoi013aa1n02x4               g208(.a(new_n289), .b(new_n292), .c(new_n290), .d(new_n278), .o1(new_n304));
  aoai13aa1n02x7               g209(.a(new_n304), .b(new_n303), .c(new_n266), .d(new_n271), .o1(new_n305));
  aoi022aa1n03x5               g210(.a(new_n305), .b(new_n301), .c(new_n300), .d(new_n302), .o1(\s[30] ));
  nand03aa1n02x5               g211(.a(new_n287), .b(new_n291), .c(new_n301), .o1(new_n307));
  nanb02aa1n03x5               g212(.a(new_n307), .b(new_n275), .out0(new_n308));
  xorc02aa1n02x5               g213(.a(\a[31] ), .b(\b[30] ), .out0(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n304), .carry(new_n310));
  norb02aa1n02x5               g215(.a(new_n310), .b(new_n309), .out0(new_n311));
  aoai13aa1n02x5               g216(.a(new_n310), .b(new_n307), .c(new_n266), .d(new_n271), .o1(new_n312));
  aoi022aa1n03x5               g217(.a(new_n312), .b(new_n309), .c(new_n308), .d(new_n311), .o1(\s[31] ));
  xorb03aa1n02x5               g218(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g219(.a(new_n105), .b(new_n107), .o1(new_n315));
  aoi112aa1n02x5               g220(.a(new_n102), .b(new_n101), .c(new_n100), .d(new_n103), .o1(new_n316));
  oaoi13aa1n02x5               g221(.a(new_n316), .b(new_n315), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g222(.a(new_n114), .b(new_n105), .c(new_n107), .out0(\s[5] ));
  nanp02aa1n03x5               g223(.a(new_n315), .b(new_n114), .o1(new_n319));
  xnbna2aa1n03x5               g224(.a(new_n113), .b(new_n319), .c(new_n117), .out0(\s[6] ));
  norb02aa1n02x5               g225(.a(new_n113), .b(new_n116), .out0(new_n321));
  ao0022aa1n03x5               g226(.a(new_n319), .b(new_n321), .c(\b[5] ), .d(\a[6] ), .o(new_n322));
  xnrb03aa1n02x5               g227(.a(new_n322), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n03x5               g228(.a(\a[7] ), .b(\b[6] ), .c(new_n322), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g230(.a(new_n121), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


