// Benchmark "adder" written by ABC on Thu Jul 18 10:38:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n348, new_n351, new_n352, new_n354, new_n355,
    new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1n08x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n03x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  nor042aa1n06x5               g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  nor002aa1n02x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  xnrc02aa1n12x5               g009(.a(\b[7] ), .b(\a[8] ), .out0(new_n105));
  nand42aa1d28x5               g010(.a(\b[5] ), .b(\a[6] ), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand42aa1n06x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nanb03aa1n03x5               g013(.a(new_n107), .b(new_n108), .c(new_n106), .out0(new_n109));
  inv000aa1d42x5               g014(.a(new_n107), .o1(new_n110));
  oao003aa1n02x5               g015(.a(\a[8] ), .b(\b[7] ), .c(new_n110), .carry(new_n111));
  oai013aa1n03x5               g016(.a(new_n111), .b(new_n109), .c(new_n105), .d(new_n104), .o1(new_n112));
  nor042aa1n02x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand02aa1d08x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nand02aa1n06x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  aoi012aa1n06x5               g020(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[4] ), .o1(new_n117));
  nanb02aa1n03x5               g022(.a(\b[3] ), .b(new_n117), .out0(new_n118));
  nanp02aa1n02x5               g023(.a(\b[3] ), .b(\a[4] ), .o1(new_n119));
  nanp02aa1n03x5               g024(.a(new_n118), .b(new_n119), .o1(new_n120));
  inv040aa1d32x5               g025(.a(\a[3] ), .o1(new_n121));
  inv030aa1d32x5               g026(.a(\b[2] ), .o1(new_n122));
  nanp02aa1n06x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  nand42aa1n04x5               g028(.a(\b[2] ), .b(\a[3] ), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(new_n123), .b(new_n124), .o1(new_n125));
  aob012aa1n02x5               g030(.a(new_n119), .b(new_n118), .c(new_n123), .out0(new_n126));
  oai013aa1n06x5               g031(.a(new_n126), .b(new_n116), .c(new_n120), .d(new_n125), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n107), .b(new_n108), .out0(new_n128));
  nand22aa1n03x5               g033(.a(\b[4] ), .b(\a[5] ), .o1(new_n129));
  nona23aa1n02x4               g034(.a(new_n106), .b(new_n129), .c(new_n103), .d(new_n102), .out0(new_n130));
  nor043aa1n03x5               g035(.a(new_n130), .b(new_n128), .c(new_n105), .o1(new_n131));
  nand42aa1n02x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  norb02aa1n06x5               g037(.a(new_n132), .b(new_n100), .out0(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n112), .c(new_n127), .d(new_n131), .o1(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n99), .b(new_n134), .c(new_n101), .out0(\s[10] ));
  oaoi03aa1n02x5               g040(.a(\a[10] ), .b(\b[9] ), .c(new_n101), .o1(new_n136));
  inv000aa1d42x5               g041(.a(new_n136), .o1(new_n137));
  norp03aa1n02x5               g042(.a(new_n109), .b(new_n105), .c(new_n104), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n111), .b(new_n138), .out0(new_n139));
  nanp02aa1n03x5               g044(.a(new_n127), .b(new_n131), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(new_n140), .b(new_n139), .o1(new_n141));
  nanp03aa1n03x5               g046(.a(new_n141), .b(new_n99), .c(new_n133), .o1(new_n142));
  norp02aa1n06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nand42aa1n06x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n142), .c(new_n137), .out0(\s[11] ));
  inv040aa1d32x5               g051(.a(\a[11] ), .o1(new_n147));
  inv000aa1d42x5               g052(.a(\b[10] ), .o1(new_n148));
  nand02aa1d12x5               g053(.a(new_n148), .b(new_n147), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n149), .b(new_n144), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n149), .b(new_n150), .c(new_n142), .d(new_n137), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv040aa1d32x5               g057(.a(\a[12] ), .o1(new_n153));
  inv000aa1d42x5               g058(.a(\b[11] ), .o1(new_n154));
  nand42aa1n08x5               g059(.a(new_n154), .b(new_n153), .o1(new_n155));
  nand42aa1n06x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  nand42aa1n02x5               g061(.a(new_n155), .b(new_n156), .o1(new_n157));
  nano32aa1n03x7               g062(.a(new_n157), .b(new_n145), .c(new_n133), .d(new_n99), .out0(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n112), .c(new_n127), .d(new_n131), .o1(new_n159));
  oai112aa1n06x5               g064(.a(new_n155), .b(new_n156), .c(new_n100), .d(new_n97), .o1(new_n160));
  nanb03aa1n09x5               g065(.a(new_n143), .b(new_n144), .c(new_n98), .out0(new_n161));
  oaoi03aa1n09x5               g066(.a(\a[12] ), .b(\b[11] ), .c(new_n149), .o1(new_n162));
  inv040aa1n02x5               g067(.a(new_n162), .o1(new_n163));
  oai012aa1d24x5               g068(.a(new_n163), .b(new_n160), .c(new_n161), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nor002aa1d32x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  nand42aa1n03x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  xobna2aa1n03x5               g073(.a(new_n168), .b(new_n159), .c(new_n165), .out0(\s[13] ));
  inv040aa1n08x5               g074(.a(new_n166), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n170), .b(new_n168), .c(new_n159), .d(new_n165), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nand02aa1n02x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nano23aa1n09x5               g079(.a(new_n166), .b(new_n173), .c(new_n174), .d(new_n167), .out0(new_n175));
  oaoi03aa1n09x5               g080(.a(\a[14] ), .b(\b[13] ), .c(new_n170), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n176), .b(new_n164), .c(new_n175), .o1(new_n177));
  nano23aa1n06x5               g082(.a(new_n97), .b(new_n100), .c(new_n132), .d(new_n98), .out0(new_n178));
  nona22aa1n09x5               g083(.a(new_n178), .b(new_n157), .c(new_n150), .out0(new_n179));
  nona23aa1n03x5               g084(.a(new_n174), .b(new_n167), .c(new_n166), .d(new_n173), .out0(new_n180));
  nona22aa1n02x4               g085(.a(new_n141), .b(new_n179), .c(new_n180), .out0(new_n181));
  nor002aa1d32x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nand42aa1d28x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n181), .c(new_n177), .out0(\s[15] ));
  inv040aa1n02x5               g090(.a(new_n182), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n184), .o1(new_n187));
  aoai13aa1n02x5               g092(.a(new_n186), .b(new_n187), .c(new_n181), .d(new_n177), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor042aa1n03x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nanp02aa1n12x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nano23aa1d15x5               g096(.a(new_n182), .b(new_n190), .c(new_n191), .d(new_n183), .out0(new_n192));
  aoai13aa1n06x5               g097(.a(new_n192), .b(new_n176), .c(new_n164), .d(new_n175), .o1(new_n193));
  oaoi03aa1n12x5               g098(.a(\a[16] ), .b(\b[15] ), .c(new_n186), .o1(new_n194));
  inv000aa1d42x5               g099(.a(new_n194), .o1(new_n195));
  nano22aa1d15x5               g100(.a(new_n179), .b(new_n175), .c(new_n192), .out0(new_n196));
  aoai13aa1n12x5               g101(.a(new_n196), .b(new_n112), .c(new_n127), .d(new_n131), .o1(new_n197));
  nand23aa1d12x5               g102(.a(new_n197), .b(new_n193), .c(new_n195), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  oaoi13aa1n06x5               g104(.a(new_n180), .b(new_n163), .c(new_n160), .d(new_n161), .o1(new_n200));
  oaoi13aa1n09x5               g105(.a(new_n194), .b(new_n192), .c(new_n200), .d(new_n176), .o1(new_n201));
  orn002aa1n02x5               g106(.a(\a[17] ), .b(\b[16] ), .o(new_n202));
  xnrc02aa1n02x5               g107(.a(\b[16] ), .b(\a[17] ), .out0(new_n203));
  aoai13aa1n03x5               g108(.a(new_n202), .b(new_n203), .c(new_n201), .d(new_n197), .o1(new_n204));
  xorb03aa1n02x5               g109(.a(new_n204), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  xorc02aa1n12x5               g110(.a(\a[18] ), .b(\b[17] ), .out0(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n203), .out0(new_n207));
  inv000aa1n02x5               g112(.a(new_n207), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  aoai13aa1n04x5               g115(.a(new_n210), .b(new_n208), .c(new_n201), .d(new_n197), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g118(.a(\a[19] ), .o1(new_n214));
  inv040aa1d28x5               g119(.a(\b[18] ), .o1(new_n215));
  nand02aa1d16x5               g120(.a(new_n215), .b(new_n214), .o1(new_n216));
  xorc02aa1n02x5               g121(.a(\a[19] ), .b(\b[18] ), .out0(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n209), .c(new_n198), .d(new_n207), .o1(new_n218));
  nor002aa1d32x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand42aa1n10x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  norb02aa1n02x5               g125(.a(new_n220), .b(new_n219), .out0(new_n221));
  aobi12aa1n06x5               g126(.a(new_n221), .b(new_n218), .c(new_n216), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n216), .o1(new_n223));
  nand42aa1n03x5               g128(.a(\b[18] ), .b(\a[19] ), .o1(new_n224));
  aoi112aa1n02x5               g129(.a(new_n223), .b(new_n221), .c(new_n211), .d(new_n224), .o1(new_n225));
  nor002aa1n02x5               g130(.a(new_n222), .b(new_n225), .o1(\s[20] ));
  nano22aa1n03x7               g131(.a(new_n219), .b(new_n224), .c(new_n220), .out0(new_n227));
  nona23aa1d18x5               g132(.a(new_n227), .b(new_n206), .c(new_n203), .d(new_n223), .out0(new_n228));
  nanb03aa1n06x5               g133(.a(new_n219), .b(new_n220), .c(new_n224), .out0(new_n229));
  nanp02aa1n02x5               g134(.a(\b[17] ), .b(\a[18] ), .o1(new_n230));
  oaih22aa1d12x5               g135(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n231));
  nand03aa1n04x5               g136(.a(new_n231), .b(new_n216), .c(new_n230), .o1(new_n232));
  aoai13aa1n12x5               g137(.a(new_n220), .b(new_n219), .c(new_n214), .d(new_n215), .o1(new_n233));
  oai012aa1d24x5               g138(.a(new_n233), .b(new_n232), .c(new_n229), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n228), .c(new_n201), .d(new_n197), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  inv000aa1n03x5               g143(.a(new_n238), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n228), .o1(new_n240));
  xnrc02aa1n12x5               g145(.a(\b[20] ), .b(\a[21] ), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n234), .c(new_n198), .d(new_n240), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[21] ), .b(\a[22] ), .out0(new_n244));
  tech160nm_fiaoi012aa1n02p5x5 g149(.a(new_n244), .b(new_n243), .c(new_n239), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n244), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n238), .b(new_n246), .c(new_n236), .d(new_n242), .o1(new_n247));
  norp02aa1n03x5               g152(.a(new_n245), .b(new_n247), .o1(\s[22] ));
  nor042aa1n06x5               g153(.a(new_n244), .b(new_n241), .o1(new_n249));
  norb02aa1n06x4               g154(.a(new_n249), .b(new_n228), .out0(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  oaoi03aa1n02x5               g156(.a(\a[22] ), .b(\b[21] ), .c(new_n239), .o1(new_n252));
  aoi012aa1n09x5               g157(.a(new_n252), .b(new_n234), .c(new_n249), .o1(new_n253));
  aoai13aa1n04x5               g158(.a(new_n253), .b(new_n251), .c(new_n201), .d(new_n197), .o1(new_n254));
  xorb03aa1n02x5               g159(.a(new_n254), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  inv000aa1n03x5               g161(.a(new_n256), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n253), .o1(new_n258));
  tech160nm_fixorc02aa1n05x5   g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n258), .c(new_n198), .d(new_n250), .o1(new_n260));
  tech160nm_fixorc02aa1n05x5   g165(.a(\a[24] ), .b(\b[23] ), .out0(new_n261));
  aobi12aa1n06x5               g166(.a(new_n261), .b(new_n260), .c(new_n257), .out0(new_n262));
  aoi112aa1n03x4               g167(.a(new_n256), .b(new_n261), .c(new_n254), .d(new_n259), .o1(new_n263));
  nor002aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(\s[24] ));
  oai012aa1n02x5               g169(.a(new_n230), .b(\b[18] ), .c(\a[19] ), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n231), .b(new_n265), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n233), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n249), .b(new_n267), .c(new_n266), .d(new_n227), .o1(new_n268));
  inv040aa1n02x5               g173(.a(new_n252), .o1(new_n269));
  and002aa1n06x5               g174(.a(new_n261), .b(new_n259), .o(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  oaoi03aa1n02x5               g176(.a(\a[24] ), .b(\b[23] ), .c(new_n257), .o1(new_n272));
  inv040aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n271), .c(new_n268), .d(new_n269), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nano32aa1n03x7               g180(.a(new_n228), .b(new_n261), .c(new_n249), .d(new_n259), .out0(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  aoai13aa1n04x5               g182(.a(new_n275), .b(new_n277), .c(new_n201), .d(new_n197), .o1(new_n278));
  xorb03aa1n02x5               g183(.a(new_n278), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  tech160nm_fixorc02aa1n05x5   g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n282), .b(new_n274), .c(new_n198), .d(new_n276), .o1(new_n283));
  tech160nm_fixorc02aa1n05x5   g188(.a(\a[26] ), .b(\b[25] ), .out0(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n283), .c(new_n281), .out0(new_n285));
  aoi112aa1n03x4               g190(.a(new_n280), .b(new_n284), .c(new_n278), .d(new_n282), .o1(new_n286));
  nor042aa1n03x5               g191(.a(new_n285), .b(new_n286), .o1(\s[26] ));
  norp02aa1n02x5               g192(.a(new_n100), .b(new_n97), .o1(new_n288));
  nano22aa1n02x4               g193(.a(new_n288), .b(new_n155), .c(new_n156), .out0(new_n289));
  nano22aa1n02x4               g194(.a(new_n143), .b(new_n98), .c(new_n144), .out0(new_n290));
  aoai13aa1n02x5               g195(.a(new_n175), .b(new_n162), .c(new_n289), .d(new_n290), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n176), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n192), .o1(new_n293));
  aoai13aa1n02x5               g198(.a(new_n195), .b(new_n293), .c(new_n291), .d(new_n292), .o1(new_n294));
  nona22aa1n02x4               g199(.a(new_n158), .b(new_n293), .c(new_n180), .out0(new_n295));
  aoi012aa1n06x5               g200(.a(new_n295), .b(new_n140), .c(new_n139), .o1(new_n296));
  and002aa1n02x5               g201(.a(new_n284), .b(new_n282), .o(new_n297));
  inv020aa1n02x5               g202(.a(new_n297), .o1(new_n298));
  nano23aa1n06x5               g203(.a(new_n298), .b(new_n228), .c(new_n270), .d(new_n249), .out0(new_n299));
  oai012aa1n06x5               g204(.a(new_n299), .b(new_n294), .c(new_n296), .o1(new_n300));
  nanp02aa1n02x5               g205(.a(\b[25] ), .b(\a[26] ), .o1(new_n301));
  oai022aa1n02x5               g206(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n302));
  aoi022aa1n06x5               g207(.a(new_n274), .b(new_n297), .c(new_n301), .d(new_n302), .o1(new_n303));
  xorc02aa1n12x5               g208(.a(\a[27] ), .b(\b[26] ), .out0(new_n304));
  xnbna2aa1n03x5               g209(.a(new_n304), .b(new_n300), .c(new_n303), .out0(\s[27] ));
  nor042aa1n03x5               g210(.a(\b[26] ), .b(\a[27] ), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n306), .o1(new_n307));
  aoai13aa1n04x5               g212(.a(new_n270), .b(new_n252), .c(new_n234), .d(new_n249), .o1(new_n308));
  nanp02aa1n02x5               g213(.a(new_n302), .b(new_n301), .o1(new_n309));
  aoai13aa1n06x5               g214(.a(new_n309), .b(new_n298), .c(new_n308), .d(new_n273), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n304), .b(new_n310), .c(new_n198), .d(new_n299), .o1(new_n311));
  xnrc02aa1n12x5               g216(.a(\b[27] ), .b(\a[28] ), .out0(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n312), .b(new_n311), .c(new_n307), .o1(new_n313));
  inv000aa1d42x5               g218(.a(new_n304), .o1(new_n314));
  tech160nm_fiaoi012aa1n02p5x5 g219(.a(new_n314), .b(new_n300), .c(new_n303), .o1(new_n315));
  nano22aa1n02x4               g220(.a(new_n315), .b(new_n307), .c(new_n312), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n313), .b(new_n316), .o1(\s[28] ));
  xnrc02aa1n02x5               g222(.a(\b[28] ), .b(\a[29] ), .out0(new_n318));
  norb02aa1n02x5               g223(.a(new_n304), .b(new_n312), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n310), .c(new_n198), .d(new_n299), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[28] ), .b(\b[27] ), .c(new_n307), .carry(new_n321));
  aoi012aa1n03x5               g226(.a(new_n318), .b(new_n320), .c(new_n321), .o1(new_n322));
  inv000aa1n02x5               g227(.a(new_n319), .o1(new_n323));
  tech160nm_fiaoi012aa1n02p5x5 g228(.a(new_n323), .b(new_n300), .c(new_n303), .o1(new_n324));
  nano22aa1n02x4               g229(.a(new_n324), .b(new_n318), .c(new_n321), .out0(new_n325));
  norp02aa1n03x5               g230(.a(new_n322), .b(new_n325), .o1(\s[29] ));
  xorb03aa1n02x5               g231(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g232(.a(\b[29] ), .b(\a[30] ), .out0(new_n328));
  norb03aa1d15x5               g233(.a(new_n304), .b(new_n318), .c(new_n312), .out0(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n310), .c(new_n198), .d(new_n299), .o1(new_n330));
  oao003aa1n02x5               g235(.a(\a[29] ), .b(\b[28] ), .c(new_n321), .carry(new_n331));
  tech160nm_fiaoi012aa1n02p5x5 g236(.a(new_n328), .b(new_n330), .c(new_n331), .o1(new_n332));
  inv000aa1d42x5               g237(.a(new_n329), .o1(new_n333));
  tech160nm_fiaoi012aa1n02p5x5 g238(.a(new_n333), .b(new_n300), .c(new_n303), .o1(new_n334));
  nano22aa1n02x4               g239(.a(new_n334), .b(new_n328), .c(new_n331), .out0(new_n335));
  norp02aa1n03x5               g240(.a(new_n332), .b(new_n335), .o1(\s[30] ));
  nanb02aa1n02x5               g241(.a(\b[30] ), .b(\a[31] ), .out0(new_n337));
  nanb02aa1n02x5               g242(.a(\a[31] ), .b(\b[30] ), .out0(new_n338));
  norb02aa1n02x5               g243(.a(new_n329), .b(new_n328), .out0(new_n339));
  aoai13aa1n06x5               g244(.a(new_n339), .b(new_n310), .c(new_n198), .d(new_n299), .o1(new_n340));
  oao003aa1n02x5               g245(.a(\a[30] ), .b(\b[29] ), .c(new_n331), .carry(new_n341));
  aoi022aa1n02x7               g246(.a(new_n340), .b(new_n341), .c(new_n338), .d(new_n337), .o1(new_n342));
  nanp02aa1n02x5               g247(.a(new_n338), .b(new_n337), .o1(new_n343));
  inv000aa1n02x5               g248(.a(new_n341), .o1(new_n344));
  nona22aa1n02x5               g249(.a(new_n340), .b(new_n344), .c(new_n343), .out0(new_n345));
  norb02aa1n03x4               g250(.a(new_n345), .b(new_n342), .out0(\s[31] ));
  xnbna2aa1n03x5               g251(.a(new_n116), .b(new_n124), .c(new_n123), .out0(\s[3] ));
  oaoi03aa1n02x5               g252(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g254(.a(new_n127), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g255(.a(new_n102), .o1(new_n351));
  tech160nm_fiaoi012aa1n05x5   g256(.a(new_n103), .b(new_n127), .c(new_n129), .o1(new_n352));
  xnbna2aa1n03x5               g257(.a(new_n352), .b(new_n351), .c(new_n106), .out0(\s[6] ));
  nano22aa1n02x4               g258(.a(new_n352), .b(new_n351), .c(new_n106), .out0(new_n354));
  tech160nm_fiao0012aa1n02p5x5 g259(.a(new_n109), .b(new_n352), .c(new_n351), .o(new_n355));
  oaib12aa1n02x5               g260(.a(new_n351), .b(new_n107), .c(new_n108), .out0(new_n356));
  oa0012aa1n02x5               g261(.a(new_n355), .b(new_n356), .c(new_n354), .o(\s[7] ));
  xobna2aa1n03x5               g262(.a(new_n105), .b(new_n355), .c(new_n110), .out0(\s[8] ));
  xnbna2aa1n03x5               g263(.a(new_n133), .b(new_n140), .c(new_n139), .out0(\s[9] ));
endmodule


