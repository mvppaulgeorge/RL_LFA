// Benchmark "adder" written by ABC on Thu Jul 11 12:52:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n179, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n304, new_n306, new_n308, new_n310, new_n312;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  norp02aa1n02x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  norp02aa1n02x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nano23aa1n02x4               g006(.a(new_n98), .b(new_n100), .c(new_n101), .d(new_n99), .out0(new_n102));
  norp02aa1n02x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  160nm_fiao0012aa1n02p5x5     g010(.a(new_n103), .b(new_n105), .c(new_n104), .o(new_n106));
  160nm_fiao0012aa1n02p5x5     g011(.a(new_n98), .b(new_n100), .c(new_n99), .o(new_n107));
  aoi012aa1n02x5               g012(.a(new_n107), .b(new_n102), .c(new_n106), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  160nm_ficinv00aa1n08x5       g014(.clk(new_n109), .clkout(new_n110));
  oao003aa1n02x5               g015(.a(\a[4] ), .b(\b[3] ), .c(new_n110), .carry(new_n111));
  xorc02aa1n02x5               g016(.a(\a[4] ), .b(\b[3] ), .out0(new_n112));
  nanp02aa1n02x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  norb02aa1n02x5               g018(.a(new_n113), .b(new_n109), .out0(new_n114));
  and002aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o(new_n115));
  nanp02aa1n02x5               g020(.a(\b[0] ), .b(\a[1] ), .o1(new_n116));
  norp02aa1n02x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  oab012aa1n02x4               g022(.a(new_n115), .b(new_n117), .c(new_n116), .out0(new_n118));
  nanp03aa1n02x5               g023(.a(new_n118), .b(new_n112), .c(new_n114), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nano23aa1n02x4               g025(.a(new_n103), .b(new_n105), .c(new_n120), .d(new_n104), .out0(new_n121));
  nanp02aa1n02x5               g026(.a(new_n121), .b(new_n102), .o1(new_n122));
  aoai13aa1n02x5               g027(.a(new_n108), .b(new_n122), .c(new_n119), .d(new_n111), .o1(new_n123));
  xorc02aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoi012aa1n02x5               g029(.a(new_n97), .b(new_n123), .c(new_n124), .o1(new_n125));
  160nm_ficinv00aa1n08x5       g030(.clk(\b[9] ), .clkout(new_n126));
  nanb02aa1n02x5               g031(.a(\a[10] ), .b(new_n126), .out0(new_n127));
  nanp02aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n125), .b(new_n128), .c(new_n127), .out0(\s[10] ));
  nanp02aa1n02x5               g034(.a(new_n127), .b(new_n128), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n124), .b(new_n130), .out0(new_n131));
  aob012aa1n02x5               g036(.a(new_n127), .b(new_n97), .c(new_n128), .out0(new_n132));
  norp02aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n132), .c(new_n123), .d(new_n131), .o1(new_n136));
  aoi112aa1n02x5               g041(.a(new_n135), .b(new_n132), .c(new_n123), .d(new_n131), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n136), .b(new_n137), .out0(\s[11] ));
  160nm_ficinv00aa1n08x5       g043(.clk(new_n133), .clkout(new_n139));
  norp02aa1n02x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n02x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n136), .c(new_n139), .out0(\s[12] ));
  nano23aa1n02x4               g048(.a(new_n133), .b(new_n140), .c(new_n141), .d(new_n134), .out0(new_n144));
  oaoi03aa1n02x5               g049(.a(\a[12] ), .b(\b[11] ), .c(new_n139), .o1(new_n145));
  160nm_fiao0012aa1n02p5x5     g050(.a(new_n145), .b(new_n144), .c(new_n132), .o(new_n146));
  nanb03aa1n02x5               g051(.a(new_n130), .b(new_n144), .c(new_n124), .out0(new_n147));
  160nm_ficinv00aa1n08x5       g052(.clk(new_n147), .clkout(new_n148));
  xnrc02aa1n02x5               g053(.a(\b[12] ), .b(\a[13] ), .out0(new_n149));
  160nm_ficinv00aa1n08x5       g054(.clk(new_n149), .clkout(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n146), .c(new_n123), .d(new_n148), .o1(new_n151));
  aoi112aa1n02x5               g056(.a(new_n146), .b(new_n150), .c(new_n123), .d(new_n148), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n151), .b(new_n152), .out0(\s[13] ));
  orn002aa1n02x5               g058(.a(\a[13] ), .b(\b[12] ), .o(new_n154));
  xnrc02aa1n02x5               g059(.a(\b[13] ), .b(\a[14] ), .out0(new_n155));
  xobna2aa1n03x5               g060(.a(new_n155), .b(new_n151), .c(new_n154), .out0(\s[14] ));
  norp02aa1n02x5               g061(.a(new_n155), .b(new_n149), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n145), .c(new_n144), .d(new_n132), .o1(new_n158));
  oao003aa1n02x5               g063(.a(\a[14] ), .b(\b[13] ), .c(new_n154), .carry(new_n159));
  nanp02aa1n02x5               g064(.a(new_n158), .b(new_n159), .o1(new_n160));
  160nm_ficinv00aa1n08x5       g065(.clk(new_n160), .clkout(new_n161));
  nona32aa1n02x4               g066(.a(new_n123), .b(new_n155), .c(new_n149), .d(new_n147), .out0(new_n162));
  xnrc02aa1n02x5               g067(.a(\b[14] ), .b(\a[15] ), .out0(new_n163));
  xobna2aa1n03x5               g068(.a(new_n163), .b(new_n162), .c(new_n161), .out0(\s[15] ));
  norp02aa1n02x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  160nm_ficinv00aa1n08x5       g070(.clk(new_n165), .clkout(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n163), .c(new_n162), .d(new_n161), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  160nm_ficinv00aa1n08x5       g073(.clk(\a[17] ), .clkout(new_n169));
  xnrc02aa1n02x5               g074(.a(\b[15] ), .b(\a[16] ), .out0(new_n170));
  norp02aa1n02x5               g075(.a(new_n170), .b(new_n163), .o1(new_n171));
  nano22aa1n02x4               g076(.a(new_n147), .b(new_n157), .c(new_n171), .out0(new_n172));
  160nm_ficinv00aa1n08x5       g077(.clk(new_n171), .clkout(new_n173));
  aoi012aa1n02x5               g078(.a(new_n173), .b(new_n158), .c(new_n159), .o1(new_n174));
  oao003aa1n02x5               g079(.a(\a[16] ), .b(\b[15] ), .c(new_n166), .carry(new_n175));
  160nm_ficinv00aa1n08x5       g080(.clk(new_n175), .clkout(new_n176));
  aoi112aa1n02x5               g081(.a(new_n174), .b(new_n176), .c(new_n123), .d(new_n172), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[16] ), .c(new_n169), .out0(\s[17] ));
  oaoi03aa1n02x5               g083(.a(\a[17] ), .b(\b[16] ), .c(new_n177), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  160nm_ficinv00aa1n08x5       g085(.clk(\a[18] ), .clkout(new_n181));
  xroi22aa1d04x5               g086(.a(new_n169), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n182));
  160nm_ficinv00aa1n08x5       g087(.clk(new_n182), .clkout(new_n183));
  aoi112aa1n02x5               g088(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n184));
  aoib12aa1n02x5               g089(.a(new_n184), .b(new_n181), .c(\b[17] ), .out0(new_n185));
  oai012aa1n02x5               g090(.a(new_n185), .b(new_n177), .c(new_n183), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g092(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g093(.a(\b[18] ), .b(\a[19] ), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(\b[18] ), .b(\a[19] ), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n190), .b(new_n189), .out0(new_n191));
  norp02aa1n02x5               g096(.a(\b[19] ), .b(\a[20] ), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(\b[19] ), .b(\a[20] ), .o1(new_n193));
  nanb02aa1n02x5               g098(.a(new_n192), .b(new_n193), .out0(new_n194));
  aoai13aa1n02x5               g099(.a(new_n194), .b(new_n189), .c(new_n186), .d(new_n191), .o1(new_n195));
  nanp02aa1n02x5               g100(.a(new_n123), .b(new_n172), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n160), .b(new_n171), .o1(new_n197));
  nanp03aa1n02x5               g102(.a(new_n196), .b(new_n197), .c(new_n175), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  aob012aa1n02x5               g104(.a(new_n199), .b(\b[17] ), .c(\a[18] ), .out0(new_n200));
  oaib12aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n181), .out0(new_n201));
  aoai13aa1n02x5               g106(.a(new_n191), .b(new_n201), .c(new_n198), .d(new_n182), .o1(new_n202));
  nona22aa1n02x4               g107(.a(new_n202), .b(new_n194), .c(new_n189), .out0(new_n203));
  nanp02aa1n02x5               g108(.a(new_n195), .b(new_n203), .o1(\s[20] ));
  nona23aa1n02x4               g109(.a(new_n193), .b(new_n190), .c(new_n189), .d(new_n192), .out0(new_n205));
  160nm_fiao0012aa1n02p5x5     g110(.a(new_n192), .b(new_n189), .c(new_n193), .o(new_n206));
  oabi12aa1n02x5               g111(.a(new_n206), .b(new_n205), .c(new_n185), .out0(new_n207));
  160nm_ficinv00aa1n08x5       g112(.clk(new_n207), .clkout(new_n208));
  norb02aa1n02x5               g113(.a(new_n182), .b(new_n205), .out0(new_n209));
  160nm_ficinv00aa1n08x5       g114(.clk(new_n209), .clkout(new_n210));
  oai012aa1n02x5               g115(.a(new_n208), .b(new_n177), .c(new_n210), .o1(new_n211));
  xorb03aa1n02x5               g116(.a(new_n211), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g117(.a(\b[20] ), .b(\a[21] ), .o1(new_n213));
  xnrc02aa1n02x5               g118(.a(\b[20] ), .b(\a[21] ), .out0(new_n214));
  160nm_ficinv00aa1n08x5       g119(.clk(new_n214), .clkout(new_n215));
  xnrc02aa1n02x5               g120(.a(\b[21] ), .b(\a[22] ), .out0(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n213), .c(new_n211), .d(new_n215), .o1(new_n217));
  aoai13aa1n02x5               g122(.a(new_n215), .b(new_n207), .c(new_n198), .d(new_n209), .o1(new_n218));
  nona22aa1n02x4               g123(.a(new_n218), .b(new_n216), .c(new_n213), .out0(new_n219));
  nanp02aa1n02x5               g124(.a(new_n217), .b(new_n219), .o1(\s[22] ));
  norp02aa1n02x5               g125(.a(new_n216), .b(new_n214), .o1(new_n221));
  160nm_ficinv00aa1n08x5       g126(.clk(\a[22] ), .clkout(new_n222));
  160nm_ficinv00aa1n08x5       g127(.clk(\b[21] ), .clkout(new_n223));
  oaoi03aa1n02x5               g128(.a(new_n222), .b(new_n223), .c(new_n213), .o1(new_n224));
  160nm_ficinv00aa1n08x5       g129(.clk(new_n224), .clkout(new_n225));
  aoi012aa1n02x5               g130(.a(new_n225), .b(new_n207), .c(new_n221), .o1(new_n226));
  nano23aa1n02x4               g131(.a(new_n189), .b(new_n192), .c(new_n193), .d(new_n190), .out0(new_n227));
  nano22aa1n02x4               g132(.a(new_n183), .b(new_n221), .c(new_n227), .out0(new_n228));
  160nm_ficinv00aa1n08x5       g133(.clk(new_n228), .clkout(new_n229));
  oai012aa1n02x5               g134(.a(new_n226), .b(new_n177), .c(new_n229), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  xnrc02aa1n02x5               g138(.a(\b[23] ), .b(\a[24] ), .out0(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n232), .c(new_n230), .d(new_n233), .o1(new_n235));
  160nm_ficinv00aa1n08x5       g140(.clk(new_n226), .clkout(new_n236));
  aoai13aa1n02x5               g141(.a(new_n233), .b(new_n236), .c(new_n198), .d(new_n228), .o1(new_n237));
  nona22aa1n02x4               g142(.a(new_n237), .b(new_n234), .c(new_n232), .out0(new_n238));
  nanp02aa1n02x5               g143(.a(new_n235), .b(new_n238), .o1(\s[24] ));
  norb02aa1n02x5               g144(.a(new_n233), .b(new_n234), .out0(new_n240));
  160nm_ficinv00aa1n08x5       g145(.clk(new_n240), .clkout(new_n241));
  nano32aa1n02x4               g146(.a(new_n241), .b(new_n182), .c(new_n221), .d(new_n227), .out0(new_n242));
  160nm_ficinv00aa1n08x5       g147(.clk(new_n242), .clkout(new_n243));
  aoai13aa1n02x5               g148(.a(new_n221), .b(new_n206), .c(new_n227), .d(new_n201), .o1(new_n244));
  orn002aa1n02x5               g149(.a(\a[23] ), .b(\b[22] ), .o(new_n245));
  oao003aa1n02x5               g150(.a(\a[24] ), .b(\b[23] ), .c(new_n245), .carry(new_n246));
  aoai13aa1n02x5               g151(.a(new_n246), .b(new_n241), .c(new_n244), .d(new_n224), .o1(new_n247));
  160nm_ficinv00aa1n08x5       g152(.clk(new_n247), .clkout(new_n248));
  oai012aa1n02x5               g153(.a(new_n248), .b(new_n177), .c(new_n243), .o1(new_n249));
  xorb03aa1n02x5               g154(.a(new_n249), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g155(.a(\b[24] ), .b(\a[25] ), .o1(new_n251));
  xorc02aa1n02x5               g156(.a(\a[25] ), .b(\b[24] ), .out0(new_n252));
  xnrc02aa1n02x5               g157(.a(\b[25] ), .b(\a[26] ), .out0(new_n253));
  aoai13aa1n02x5               g158(.a(new_n253), .b(new_n251), .c(new_n249), .d(new_n252), .o1(new_n254));
  aoai13aa1n02x5               g159(.a(new_n252), .b(new_n247), .c(new_n198), .d(new_n242), .o1(new_n255));
  nona22aa1n02x4               g160(.a(new_n255), .b(new_n253), .c(new_n251), .out0(new_n256));
  nanp02aa1n02x5               g161(.a(new_n254), .b(new_n256), .o1(\s[26] ));
  norb02aa1n02x5               g162(.a(new_n252), .b(new_n253), .out0(new_n258));
  160nm_ficinv00aa1n08x5       g163(.clk(\a[26] ), .clkout(new_n259));
  160nm_ficinv00aa1n08x5       g164(.clk(\b[25] ), .clkout(new_n260));
  oaoi03aa1n02x5               g165(.a(new_n259), .b(new_n260), .c(new_n251), .o1(new_n261));
  160nm_ficinv00aa1n08x5       g166(.clk(new_n261), .clkout(new_n262));
  aoi012aa1n02x5               g167(.a(new_n262), .b(new_n247), .c(new_n258), .o1(new_n263));
  160nm_ficinv00aa1n08x5       g168(.clk(new_n258), .clkout(new_n264));
  nona22aa1n02x4               g169(.a(new_n228), .b(new_n264), .c(new_n241), .out0(new_n265));
  oai012aa1n02x5               g170(.a(new_n263), .b(new_n177), .c(new_n265), .o1(new_n266));
  xorb03aa1n02x5               g171(.a(new_n266), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  xorc02aa1n02x5               g173(.a(\a[27] ), .b(\b[26] ), .out0(new_n269));
  xnrc02aa1n02x5               g174(.a(\b[27] ), .b(\a[28] ), .out0(new_n270));
  aoai13aa1n02x5               g175(.a(new_n270), .b(new_n268), .c(new_n266), .d(new_n269), .o1(new_n271));
  aoai13aa1n02x5               g176(.a(new_n240), .b(new_n225), .c(new_n207), .d(new_n221), .o1(new_n272));
  aoai13aa1n02x5               g177(.a(new_n261), .b(new_n264), .c(new_n272), .d(new_n246), .o1(new_n273));
  160nm_ficinv00aa1n08x5       g178(.clk(new_n265), .clkout(new_n274));
  aoai13aa1n02x5               g179(.a(new_n269), .b(new_n273), .c(new_n198), .d(new_n274), .o1(new_n275));
  nona22aa1n02x4               g180(.a(new_n275), .b(new_n270), .c(new_n268), .out0(new_n276));
  nanp02aa1n02x5               g181(.a(new_n271), .b(new_n276), .o1(\s[28] ));
  norb02aa1n02x5               g182(.a(new_n269), .b(new_n270), .out0(new_n278));
  aoai13aa1n02x5               g183(.a(new_n278), .b(new_n273), .c(new_n198), .d(new_n274), .o1(new_n279));
  aob012aa1n02x5               g184(.a(new_n268), .b(\b[27] ), .c(\a[28] ), .out0(new_n280));
  oa0012aa1n02x5               g185(.a(new_n280), .b(\b[27] ), .c(\a[28] ), .o(new_n281));
  160nm_ficinv00aa1n08x5       g186(.clk(new_n281), .clkout(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[28] ), .b(\a[29] ), .out0(new_n283));
  nona22aa1n02x4               g188(.a(new_n279), .b(new_n282), .c(new_n283), .out0(new_n284));
  aoai13aa1n02x5               g189(.a(new_n283), .b(new_n282), .c(new_n266), .d(new_n278), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n285), .b(new_n284), .o1(\s[29] ));
  xorb03aa1n02x5               g191(.a(new_n116), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g192(.a(new_n269), .b(new_n283), .c(new_n270), .out0(new_n288));
  oaoi03aa1n02x5               g193(.a(\a[29] ), .b(\b[28] ), .c(new_n281), .o1(new_n289));
  xnrc02aa1n02x5               g194(.a(\b[29] ), .b(\a[30] ), .out0(new_n290));
  aoai13aa1n02x5               g195(.a(new_n290), .b(new_n289), .c(new_n266), .d(new_n288), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n288), .b(new_n273), .c(new_n198), .d(new_n274), .o1(new_n292));
  nona22aa1n02x4               g197(.a(new_n292), .b(new_n289), .c(new_n290), .out0(new_n293));
  nanp02aa1n02x5               g198(.a(new_n291), .b(new_n293), .o1(\s[30] ));
  nanb02aa1n02x5               g199(.a(new_n290), .b(new_n289), .out0(new_n295));
  oai012aa1n02x5               g200(.a(new_n295), .b(\b[29] ), .c(\a[30] ), .o1(new_n296));
  norb02aa1n02x5               g201(.a(new_n288), .b(new_n290), .out0(new_n297));
  aoai13aa1n02x5               g202(.a(new_n297), .b(new_n273), .c(new_n198), .d(new_n274), .o1(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[30] ), .b(\a[31] ), .out0(new_n299));
  nona22aa1n02x4               g204(.a(new_n298), .b(new_n299), .c(new_n296), .out0(new_n300));
  aoai13aa1n02x5               g205(.a(new_n299), .b(new_n296), .c(new_n266), .d(new_n297), .o1(new_n301));
  nanp02aa1n02x5               g206(.a(new_n301), .b(new_n300), .o1(\s[31] ));
  xobna2aa1n03x5               g207(.a(new_n118), .b(new_n113), .c(new_n110), .out0(\s[3] ));
  oai012aa1n02x5               g208(.a(new_n113), .b(new_n118), .c(new_n109), .o1(new_n304));
  xnrb03aa1n02x5               g209(.a(new_n304), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  nanp02aa1n02x5               g210(.a(new_n119), .b(new_n111), .o1(new_n306));
  xorb03aa1n02x5               g211(.a(new_n306), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g212(.a(new_n105), .b(new_n306), .c(new_n120), .o1(new_n308));
  xnrb03aa1n02x5               g213(.a(new_n308), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  160nm_fiao0012aa1n02p5x5     g214(.a(new_n106), .b(new_n306), .c(new_n121), .o(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g216(.a(new_n100), .b(new_n310), .c(new_n101), .o1(new_n312));
  xnrb03aa1n02x5               g217(.a(new_n312), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g218(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


