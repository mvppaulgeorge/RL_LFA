// Benchmark "adder" written by ABC on Wed Jul 17 18:15:03 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n338,
    new_n339, new_n340, new_n342, new_n343, new_n344, new_n346, new_n348,
    new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n04x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nand42aa1n20x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nano23aa1d12x5               g005(.a(new_n97), .b(new_n99), .c(new_n100), .d(new_n98), .out0(new_n101));
  nona23aa1n02x4               g006(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n102));
  nor022aa1n04x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nanp02aa1n03x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nor042aa1n04x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  tech160nm_fiaoi012aa1n04x5   g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  ao0012aa1n03x5               g011(.a(new_n97), .b(new_n99), .c(new_n98), .o(new_n107));
  oabi12aa1n03x5               g012(.a(new_n107), .b(new_n102), .c(new_n106), .out0(new_n108));
  oa0022aa1n09x5               g013(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n109));
  inv040aa1d32x5               g014(.a(\a[3] ), .o1(new_n110));
  inv040aa1d28x5               g015(.a(\b[2] ), .o1(new_n111));
  nand02aa1n04x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nand42aa1n02x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nand22aa1n04x5               g018(.a(new_n112), .b(new_n113), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand22aa1n12x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  oai012aa1n12x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  oai012aa1n18x5               g023(.a(new_n109), .b(new_n118), .c(new_n114), .o1(new_n119));
  nanp02aa1n04x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nand02aa1n06x5               g025(.a(\b[3] ), .b(\a[4] ), .o1(new_n121));
  tech160nm_fioai012aa1n04x5   g026(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .o1(new_n122));
  nano23aa1n06x5               g027(.a(new_n122), .b(new_n103), .c(new_n104), .d(new_n120), .out0(new_n123));
  aoi013aa1n06x4               g028(.a(new_n108), .b(new_n119), .c(new_n101), .d(new_n123), .o1(new_n124));
  tech160nm_fioaoi03aa1n03p5x5 g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  xorb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n03x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  aoib12aa1n06x5               g032(.a(new_n107), .b(new_n101), .c(new_n106), .out0(new_n128));
  nand23aa1n06x5               g033(.a(new_n119), .b(new_n101), .c(new_n123), .o1(new_n129));
  nanp02aa1n12x5               g034(.a(new_n129), .b(new_n128), .o1(new_n130));
  xorc02aa1n12x5               g035(.a(\a[9] ), .b(\b[8] ), .out0(new_n131));
  nor022aa1n12x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nand22aa1n04x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norb02aa1n09x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  aoai13aa1n02x5               g039(.a(new_n134), .b(new_n127), .c(new_n130), .d(new_n131), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n132), .b(new_n127), .c(new_n133), .o1(new_n136));
  nor002aa1n16x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand42aa1d28x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n135), .c(new_n136), .out0(\s[11] ));
  nor042aa1n03x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nand42aa1n08x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  inv000aa1n02x5               g048(.a(new_n143), .o1(new_n144));
  inv020aa1n02x5               g049(.a(new_n136), .o1(new_n145));
  aoi112aa1n03x5               g050(.a(new_n137), .b(new_n145), .c(new_n125), .d(new_n134), .o1(new_n146));
  nano22aa1n03x5               g051(.a(new_n146), .b(new_n138), .c(new_n144), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n138), .o1(new_n148));
  oai012aa1n03x5               g053(.a(new_n143), .b(new_n146), .c(new_n148), .o1(new_n149));
  nanb02aa1n03x5               g054(.a(new_n147), .b(new_n149), .out0(\s[12] ));
  nano23aa1n03x7               g055(.a(new_n137), .b(new_n141), .c(new_n142), .d(new_n138), .out0(new_n151));
  nand23aa1n03x5               g056(.a(new_n151), .b(new_n131), .c(new_n134), .o1(new_n152));
  nanp02aa1n03x5               g057(.a(new_n127), .b(new_n133), .o1(new_n153));
  nona22aa1n03x5               g058(.a(new_n153), .b(new_n137), .c(new_n132), .out0(new_n154));
  aoai13aa1n09x5               g059(.a(new_n142), .b(new_n141), .c(new_n154), .d(new_n138), .o1(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n152), .c(new_n129), .d(new_n128), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n08x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nanp02aa1n04x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  aoi012aa1n02x5               g064(.a(new_n158), .b(new_n156), .c(new_n159), .o1(new_n160));
  xnrb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand22aa1n09x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nano23aa1n06x5               g068(.a(new_n158), .b(new_n162), .c(new_n163), .d(new_n159), .out0(new_n164));
  nanp02aa1n03x5               g069(.a(new_n156), .b(new_n164), .o1(new_n165));
  aoi012aa1n02x5               g070(.a(new_n162), .b(new_n158), .c(new_n163), .o1(new_n166));
  orn002aa1n24x5               g071(.a(\a[15] ), .b(\b[14] ), .o(new_n167));
  nand22aa1n09x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand02aa1d28x5               g073(.a(new_n167), .b(new_n168), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  xnbna2aa1n03x5               g075(.a(new_n170), .b(new_n165), .c(new_n166), .out0(\s[15] ));
  nand22aa1n03x5               g076(.a(new_n165), .b(new_n166), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n167), .o1(new_n173));
  xnrc02aa1n12x5               g078(.a(\b[15] ), .b(\a[16] ), .out0(new_n174));
  aoai13aa1n03x5               g079(.a(new_n174), .b(new_n173), .c(new_n172), .d(new_n168), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n172), .b(new_n170), .o1(new_n176));
  nona22aa1n02x4               g081(.a(new_n176), .b(new_n174), .c(new_n173), .out0(new_n177));
  nanp02aa1n02x5               g082(.a(new_n177), .b(new_n175), .o1(\s[16] ));
  nona22aa1n09x5               g083(.a(new_n164), .b(new_n174), .c(new_n169), .out0(new_n179));
  nor042aa1n06x5               g084(.a(new_n179), .b(new_n152), .o1(new_n180));
  nand02aa1d06x5               g085(.a(new_n130), .b(new_n180), .o1(new_n181));
  aoi112aa1n03x4               g086(.a(new_n132), .b(new_n137), .c(new_n127), .d(new_n133), .o1(new_n182));
  oai022aa1n03x5               g087(.a(new_n182), .b(new_n148), .c(\b[11] ), .d(\a[12] ), .o1(new_n183));
  nona23aa1n09x5               g088(.a(new_n163), .b(new_n159), .c(new_n158), .d(new_n162), .out0(new_n184));
  nor043aa1n06x5               g089(.a(new_n184), .b(new_n169), .c(new_n174), .o1(new_n185));
  orn002aa1n02x5               g090(.a(\a[16] ), .b(\b[15] ), .o(new_n186));
  and002aa1n02x5               g091(.a(\b[15] ), .b(\a[16] ), .o(new_n187));
  aoai13aa1n06x5               g092(.a(new_n168), .b(new_n162), .c(new_n158), .d(new_n163), .o1(new_n188));
  aoai13aa1n06x5               g093(.a(new_n186), .b(new_n187), .c(new_n188), .d(new_n167), .o1(new_n189));
  aoi013aa1n06x4               g094(.a(new_n189), .b(new_n185), .c(new_n183), .d(new_n142), .o1(new_n190));
  xorc02aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n181), .c(new_n190), .out0(\s[17] ));
  inv040aa1d32x5               g097(.a(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[16] ), .o1(new_n194));
  nand42aa1n02x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  oabi12aa1n12x5               g100(.a(new_n189), .b(new_n155), .c(new_n179), .out0(new_n196));
  aoai13aa1n02x5               g101(.a(new_n191), .b(new_n196), .c(new_n130), .d(new_n180), .o1(new_n197));
  nor002aa1d32x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nand22aa1n12x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nanb02aa1n06x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  xobna2aa1n03x5               g105(.a(new_n200), .b(new_n197), .c(new_n195), .out0(\s[18] ));
  nanp02aa1n02x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  nano22aa1n12x5               g107(.a(new_n200), .b(new_n195), .c(new_n202), .out0(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n196), .c(new_n130), .d(new_n180), .o1(new_n204));
  aoi013aa1n09x5               g109(.a(new_n198), .b(new_n199), .c(new_n193), .d(new_n194), .o1(new_n205));
  nor002aa1d32x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand22aa1n09x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  norb02aa1n06x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n204), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n04x5               g115(.a(new_n204), .b(new_n205), .o1(new_n211));
  nor002aa1d32x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand02aa1d28x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n15x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n02x5               g120(.a(new_n215), .b(new_n206), .c(new_n211), .d(new_n207), .o1(new_n216));
  nanb02aa1n06x5               g121(.a(new_n152), .b(new_n185), .out0(new_n217));
  oai012aa1n06x5               g122(.a(new_n190), .b(new_n124), .c(new_n217), .o1(new_n218));
  oaoi03aa1n02x5               g123(.a(\a[18] ), .b(\b[17] ), .c(new_n195), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n208), .b(new_n219), .c(new_n218), .d(new_n203), .o1(new_n220));
  nona22aa1n03x5               g125(.a(new_n220), .b(new_n215), .c(new_n206), .out0(new_n221));
  nanp02aa1n03x5               g126(.a(new_n216), .b(new_n221), .o1(\s[20] ));
  nano23aa1n06x5               g127(.a(new_n206), .b(new_n212), .c(new_n213), .d(new_n207), .out0(new_n223));
  nand02aa1d06x5               g128(.a(new_n203), .b(new_n223), .o1(new_n224));
  nona23aa1n09x5               g129(.a(new_n213), .b(new_n207), .c(new_n206), .d(new_n212), .out0(new_n225));
  oai012aa1d24x5               g130(.a(new_n213), .b(new_n212), .c(new_n206), .o1(new_n226));
  oai012aa1n18x5               g131(.a(new_n226), .b(new_n225), .c(new_n205), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n04x5               g133(.a(new_n228), .b(new_n224), .c(new_n181), .d(new_n190), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv040aa1n02x5               g135(.a(new_n230), .o1(new_n231));
  inv040aa1n03x5               g136(.a(new_n224), .o1(new_n232));
  aoi112aa1n02x5               g137(.a(new_n231), .b(new_n227), .c(new_n218), .d(new_n232), .o1(new_n233));
  aoi012aa1n02x5               g138(.a(new_n233), .b(new_n229), .c(new_n231), .o1(\s[21] ));
  nor042aa1d18x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[21] ), .b(\a[22] ), .out0(new_n236));
  aoai13aa1n03x5               g141(.a(new_n236), .b(new_n235), .c(new_n229), .d(new_n231), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n231), .b(new_n227), .c(new_n218), .d(new_n232), .o1(new_n238));
  nona22aa1n03x5               g143(.a(new_n238), .b(new_n236), .c(new_n235), .out0(new_n239));
  nanp02aa1n03x5               g144(.a(new_n237), .b(new_n239), .o1(\s[22] ));
  nanb02aa1n06x5               g145(.a(new_n236), .b(new_n231), .out0(new_n241));
  nano22aa1n02x4               g146(.a(new_n241), .b(new_n203), .c(new_n223), .out0(new_n242));
  aoai13aa1n06x5               g147(.a(new_n242), .b(new_n196), .c(new_n130), .d(new_n180), .o1(new_n243));
  aoi112aa1n09x5               g148(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n244));
  oai112aa1n06x5               g149(.a(new_n208), .b(new_n214), .c(new_n244), .d(new_n198), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oao003aa1n03x5               g152(.a(new_n246), .b(new_n247), .c(new_n235), .carry(new_n248));
  inv040aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n241), .c(new_n245), .d(new_n226), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  xorc02aa1n12x5               g156(.a(\a[23] ), .b(\b[22] ), .out0(new_n252));
  xnbna2aa1n03x5               g157(.a(new_n252), .b(new_n243), .c(new_n251), .out0(\s[23] ));
  tech160nm_finand02aa1n03p5x5 g158(.a(new_n243), .b(new_n251), .o1(new_n254));
  nor042aa1n03x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  xnrc02aa1n02x5               g160(.a(\b[23] ), .b(\a[24] ), .out0(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n255), .c(new_n254), .d(new_n252), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n252), .b(new_n250), .c(new_n218), .d(new_n242), .o1(new_n258));
  nona22aa1n03x5               g163(.a(new_n258), .b(new_n256), .c(new_n255), .out0(new_n259));
  nanp02aa1n03x5               g164(.a(new_n257), .b(new_n259), .o1(\s[24] ));
  norp02aa1n04x5               g165(.a(new_n236), .b(new_n230), .o1(new_n261));
  norb02aa1n02x7               g166(.a(new_n252), .b(new_n256), .out0(new_n262));
  nanb03aa1n02x5               g167(.a(new_n224), .b(new_n262), .c(new_n261), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n226), .o1(new_n264));
  aoai13aa1n06x5               g169(.a(new_n261), .b(new_n264), .c(new_n223), .d(new_n219), .o1(new_n265));
  nanb02aa1n12x5               g170(.a(new_n256), .b(new_n252), .out0(new_n266));
  inv000aa1d42x5               g171(.a(\a[24] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(\b[23] ), .o1(new_n268));
  oao003aa1n02x5               g173(.a(new_n267), .b(new_n268), .c(new_n255), .carry(new_n269));
  inv030aa1n02x5               g174(.a(new_n269), .o1(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n266), .c(new_n265), .d(new_n249), .o1(new_n271));
  inv040aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n263), .c(new_n181), .d(new_n190), .o1(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  xnrc02aa1n12x5               g181(.a(\b[25] ), .b(\a[26] ), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n275), .c(new_n273), .d(new_n276), .o1(new_n278));
  nand42aa1n02x5               g183(.a(new_n273), .b(new_n276), .o1(new_n279));
  nona22aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n280), .b(new_n278), .o1(\s[26] ));
  norb02aa1n12x5               g186(.a(new_n276), .b(new_n277), .out0(new_n282));
  nano23aa1n06x5               g187(.a(new_n224), .b(new_n266), .c(new_n282), .d(new_n261), .out0(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n196), .c(new_n130), .d(new_n180), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n282), .b(new_n269), .c(new_n250), .d(new_n262), .o1(new_n285));
  inv000aa1d42x5               g190(.a(\a[26] ), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\b[25] ), .o1(new_n287));
  oao003aa1n02x5               g192(.a(new_n286), .b(new_n287), .c(new_n275), .carry(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  nanp03aa1n03x5               g194(.a(new_n284), .b(new_n285), .c(new_n289), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  aoi112aa1n02x5               g196(.a(new_n291), .b(new_n288), .c(new_n271), .d(new_n282), .o1(new_n292));
  aoi022aa1n02x5               g197(.a(new_n290), .b(new_n291), .c(new_n292), .d(new_n284), .o1(\s[27] ));
  nor042aa1n03x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  xnrc02aa1n12x5               g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n290), .d(new_n291), .o1(new_n296));
  nona23aa1n09x5               g201(.a(new_n232), .b(new_n282), .c(new_n241), .d(new_n266), .out0(new_n297));
  oaoi13aa1n12x5               g202(.a(new_n297), .b(new_n190), .c(new_n124), .d(new_n217), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n262), .b(new_n248), .c(new_n227), .d(new_n261), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n282), .o1(new_n300));
  aoai13aa1n04x5               g205(.a(new_n289), .b(new_n300), .c(new_n299), .d(new_n270), .o1(new_n301));
  oaih12aa1n02x5               g206(.a(new_n291), .b(new_n301), .c(new_n298), .o1(new_n302));
  nona22aa1n02x4               g207(.a(new_n302), .b(new_n295), .c(new_n294), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n296), .b(new_n303), .o1(\s[28] ));
  norb02aa1n03x5               g209(.a(new_n291), .b(new_n295), .out0(new_n305));
  oaih12aa1n02x5               g210(.a(new_n305), .b(new_n301), .c(new_n298), .o1(new_n306));
  xorc02aa1n12x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  inv000aa1d42x5               g212(.a(\a[28] ), .o1(new_n308));
  inv000aa1d42x5               g213(.a(\b[27] ), .o1(new_n309));
  aoi112aa1n02x5               g214(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n310));
  aoi112aa1n02x5               g215(.a(new_n307), .b(new_n310), .c(new_n308), .d(new_n309), .o1(new_n311));
  aoi012aa1n03x5               g216(.a(new_n288), .b(new_n271), .c(new_n282), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n305), .o1(new_n313));
  oao003aa1n06x5               g218(.a(new_n308), .b(new_n309), .c(new_n294), .carry(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n02x7               g220(.a(new_n315), .b(new_n313), .c(new_n312), .d(new_n284), .o1(new_n316));
  aoi022aa1n03x5               g221(.a(new_n316), .b(new_n307), .c(new_n306), .d(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g222(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g223(.a(new_n295), .b(new_n291), .c(new_n307), .out0(new_n319));
  oaih12aa1n02x5               g224(.a(new_n319), .b(new_n301), .c(new_n298), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .out0(new_n321));
  inv000aa1d42x5               g226(.a(\a[29] ), .o1(new_n322));
  inv000aa1d42x5               g227(.a(\b[28] ), .o1(new_n323));
  oabi12aa1n02x5               g228(.a(new_n321), .b(\a[29] ), .c(\b[28] ), .out0(new_n324));
  oaoi13aa1n02x5               g229(.a(new_n324), .b(new_n314), .c(new_n322), .d(new_n323), .o1(new_n325));
  inv000aa1n02x5               g230(.a(new_n319), .o1(new_n326));
  tech160nm_fioaoi03aa1n03p5x5 g231(.a(new_n322), .b(new_n323), .c(new_n314), .o1(new_n327));
  aoai13aa1n02x7               g232(.a(new_n327), .b(new_n326), .c(new_n312), .d(new_n284), .o1(new_n328));
  aoi022aa1n03x5               g233(.a(new_n328), .b(new_n321), .c(new_n320), .d(new_n325), .o1(\s[30] ));
  nanp03aa1n02x5               g234(.a(new_n305), .b(new_n307), .c(new_n321), .o1(new_n330));
  oabi12aa1n02x5               g235(.a(new_n330), .b(new_n301), .c(new_n298), .out0(new_n331));
  xorc02aa1n02x5               g236(.a(\a[31] ), .b(\b[30] ), .out0(new_n332));
  oao003aa1n02x5               g237(.a(\a[30] ), .b(\b[29] ), .c(new_n327), .carry(new_n333));
  norb02aa1n02x5               g238(.a(new_n333), .b(new_n332), .out0(new_n334));
  aoai13aa1n02x7               g239(.a(new_n333), .b(new_n330), .c(new_n312), .d(new_n284), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n335), .b(new_n332), .c(new_n331), .d(new_n334), .o1(\s[31] ));
  xnbna2aa1n03x5               g241(.a(new_n118), .b(new_n112), .c(new_n113), .out0(\s[3] ));
  orn002aa1n02x5               g242(.a(new_n118), .b(new_n114), .o(new_n338));
  xorc02aa1n02x5               g243(.a(\a[4] ), .b(\b[3] ), .out0(new_n339));
  norb02aa1n02x5               g244(.a(new_n112), .b(new_n339), .out0(new_n340));
  aoi022aa1n02x5               g245(.a(new_n338), .b(new_n340), .c(new_n119), .d(new_n339), .o1(\s[4] ));
  nano22aa1n02x4               g246(.a(new_n105), .b(new_n120), .c(new_n121), .out0(new_n342));
  nanb02aa1n02x5               g247(.a(new_n105), .b(new_n120), .out0(new_n343));
  nanp02aa1n02x5               g248(.a(new_n119), .b(new_n121), .o1(new_n344));
  aoi022aa1n02x5               g249(.a(new_n344), .b(new_n343), .c(new_n119), .d(new_n342), .o1(\s[5] ));
  aoi012aa1n02x5               g250(.a(new_n105), .b(new_n119), .c(new_n342), .o1(new_n346));
  xnrb03aa1n02x5               g251(.a(new_n346), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aob012aa1n02x5               g252(.a(new_n106), .b(new_n119), .c(new_n123), .out0(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g254(.a(new_n99), .b(new_n348), .c(new_n100), .o1(new_n350));
  xnrb03aa1n02x5               g255(.a(new_n350), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g256(.a(new_n131), .b(new_n129), .c(new_n128), .out0(\s[9] ));
endmodule


