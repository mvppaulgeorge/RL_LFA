// Benchmark "adder" written by ABC on Thu Jul 18 08:13:17 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n338, new_n340, new_n343, new_n344, new_n347, new_n348, new_n349,
    new_n351, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv030aa1d32x5               g003(.a(\a[2] ), .o1(new_n99));
  inv020aa1d32x5               g004(.a(\b[1] ), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(new_n100), .b(new_n99), .o1(new_n101));
  nand42aa1n08x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nand42aa1d28x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  aob012aa1n12x5               g008(.a(new_n101), .b(new_n102), .c(new_n103), .out0(new_n104));
  xorc02aa1n12x5               g009(.a(\a[4] ), .b(\b[3] ), .out0(new_n105));
  xorc02aa1n12x5               g010(.a(\a[3] ), .b(\b[2] ), .out0(new_n106));
  nand03aa1n06x5               g011(.a(new_n104), .b(new_n105), .c(new_n106), .o1(new_n107));
  nor042aa1n06x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  inv040aa1n03x5               g013(.a(new_n108), .o1(new_n109));
  oao003aa1n09x5               g014(.a(\a[4] ), .b(\b[3] ), .c(new_n109), .carry(new_n110));
  nanp02aa1n03x5               g015(.a(new_n107), .b(new_n110), .o1(new_n111));
  nor022aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand02aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  norb02aa1n03x5               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  xnrc02aa1n12x5               g019(.a(\b[4] ), .b(\a[5] ), .out0(new_n115));
  inv000aa1d42x5               g020(.a(new_n115), .o1(new_n116));
  xorc02aa1n12x5               g021(.a(\a[8] ), .b(\b[7] ), .out0(new_n117));
  xorc02aa1n12x5               g022(.a(\a[7] ), .b(\b[6] ), .out0(new_n118));
  nanp02aa1n02x5               g023(.a(new_n118), .b(new_n117), .o1(new_n119));
  nano22aa1n03x7               g024(.a(new_n119), .b(new_n116), .c(new_n114), .out0(new_n120));
  inv000aa1n04x5               g025(.a(new_n112), .o1(new_n121));
  nor042aa1n03x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  aob012aa1n06x5               g027(.a(new_n121), .b(new_n122), .c(new_n113), .out0(new_n123));
  orn002aa1n03x5               g028(.a(\a[7] ), .b(\b[6] ), .o(new_n124));
  oaoi03aa1n09x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  aoi013aa1n06x4               g030(.a(new_n125), .b(new_n123), .c(new_n118), .d(new_n117), .o1(new_n126));
  inv020aa1n02x5               g031(.a(new_n126), .o1(new_n127));
  tech160nm_fixorc02aa1n02p5x5 g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n111), .d(new_n120), .o1(new_n129));
  xorc02aa1n02x5               g034(.a(\a[10] ), .b(\b[9] ), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  xnrc02aa1n02x5               g036(.a(\b[6] ), .b(\a[7] ), .out0(new_n132));
  nona23aa1n09x5               g037(.a(new_n117), .b(new_n114), .c(new_n132), .d(new_n115), .out0(new_n133));
  aoai13aa1n06x5               g038(.a(new_n126), .b(new_n133), .c(new_n107), .d(new_n110), .o1(new_n134));
  inv000aa1d42x5               g039(.a(\a[10] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(\b[8] ), .o1(new_n136));
  xroi22aa1d04x5               g041(.a(new_n135), .b(\b[9] ), .c(new_n136), .d(\a[9] ), .out0(new_n137));
  aoi112aa1n09x5               g042(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n138));
  aoib12aa1n06x5               g043(.a(new_n138), .b(new_n135), .c(\b[9] ), .out0(new_n139));
  inv000aa1n02x5               g044(.a(new_n139), .o1(new_n140));
  xnrc02aa1n12x5               g045(.a(\b[10] ), .b(\a[11] ), .out0(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  aoai13aa1n03x5               g047(.a(new_n142), .b(new_n140), .c(new_n134), .d(new_n137), .o1(new_n143));
  aoi112aa1n02x5               g048(.a(new_n142), .b(new_n140), .c(new_n134), .d(new_n137), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(\s[11] ));
  nor002aa1n04x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nanp02aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nanb02aa1n06x5               g052(.a(new_n146), .b(new_n147), .out0(new_n148));
  nor002aa1n02x5               g053(.a(\b[10] ), .b(\a[11] ), .o1(new_n149));
  aoib12aa1n02x5               g054(.a(new_n149), .b(new_n147), .c(new_n146), .out0(new_n150));
  oai012aa1n03x5               g055(.a(new_n143), .b(\b[10] ), .c(\a[11] ), .o1(new_n151));
  aboi22aa1n03x5               g056(.a(new_n148), .b(new_n151), .c(new_n143), .d(new_n150), .out0(\s[12] ));
  nano23aa1n02x4               g057(.a(new_n148), .b(new_n141), .c(new_n130), .d(new_n128), .out0(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n127), .c(new_n111), .d(new_n120), .o1(new_n154));
  nor042aa1n04x5               g059(.a(new_n141), .b(new_n148), .o1(new_n155));
  oai012aa1n02x5               g060(.a(new_n147), .b(new_n146), .c(new_n149), .o1(new_n156));
  aobi12aa1n06x5               g061(.a(new_n156), .b(new_n155), .c(new_n140), .out0(new_n157));
  nanp02aa1n06x5               g062(.a(new_n154), .b(new_n157), .o1(new_n158));
  tech160nm_fixnrc02aa1n05x5   g063(.a(\b[12] ), .b(\a[13] ), .out0(new_n159));
  nanp02aa1n02x5               g064(.a(new_n159), .b(new_n156), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n160), .b(new_n155), .c(new_n140), .o1(new_n161));
  aboi22aa1n03x5               g066(.a(new_n159), .b(new_n158), .c(new_n161), .d(new_n154), .out0(\s[13] ));
  nanb02aa1n06x5               g067(.a(new_n159), .b(new_n158), .out0(new_n163));
  xnrc02aa1n12x5               g068(.a(\b[13] ), .b(\a[14] ), .out0(new_n164));
  nor002aa1d32x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  tech160nm_fioai012aa1n03p5x5 g071(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .o1(new_n167));
  aboi22aa1n03x5               g072(.a(new_n164), .b(new_n167), .c(new_n163), .d(new_n166), .out0(\s[14] ));
  oai013aa1n03x5               g073(.a(new_n156), .b(new_n139), .c(new_n141), .d(new_n148), .o1(new_n169));
  nor042aa1n02x5               g074(.a(new_n164), .b(new_n159), .o1(new_n170));
  aoai13aa1n03x5               g075(.a(new_n170), .b(new_n169), .c(new_n134), .d(new_n153), .o1(new_n171));
  inv000aa1d42x5               g076(.a(\a[14] ), .o1(new_n172));
  inv040aa1d32x5               g077(.a(\b[13] ), .o1(new_n173));
  oaoi03aa1n12x5               g078(.a(new_n172), .b(new_n173), .c(new_n165), .o1(new_n174));
  xnrc02aa1n12x5               g079(.a(\b[14] ), .b(\a[15] ), .out0(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n171), .c(new_n174), .out0(\s[15] ));
  inv000aa1d42x5               g082(.a(new_n174), .o1(new_n178));
  aoai13aa1n03x5               g083(.a(new_n176), .b(new_n178), .c(new_n158), .d(new_n170), .o1(new_n179));
  xnrc02aa1n12x5               g084(.a(\b[15] ), .b(\a[16] ), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  nor042aa1d18x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n180), .b(new_n182), .out0(new_n183));
  inv000aa1n02x5               g088(.a(new_n182), .o1(new_n184));
  aoai13aa1n03x5               g089(.a(new_n184), .b(new_n175), .c(new_n171), .d(new_n174), .o1(new_n185));
  aoi022aa1n03x5               g090(.a(new_n185), .b(new_n181), .c(new_n179), .d(new_n183), .o1(\s[16] ));
  nona22aa1n09x5               g091(.a(new_n170), .b(new_n175), .c(new_n180), .out0(new_n187));
  nano22aa1n12x5               g092(.a(new_n187), .b(new_n137), .c(new_n155), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n127), .c(new_n120), .d(new_n111), .o1(new_n189));
  oao003aa1n02x5               g094(.a(\a[16] ), .b(\b[15] ), .c(new_n184), .carry(new_n190));
  oai013aa1n02x4               g095(.a(new_n190), .b(new_n174), .c(new_n175), .d(new_n180), .o1(new_n191));
  aoib12aa1n06x5               g096(.a(new_n191), .b(new_n169), .c(new_n187), .out0(new_n192));
  nanp02aa1n09x5               g097(.a(new_n189), .b(new_n192), .o1(new_n193));
  xorc02aa1n12x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  norb02aa1n02x5               g099(.a(new_n190), .b(new_n194), .out0(new_n195));
  oai013aa1n02x4               g100(.a(new_n195), .b(new_n175), .c(new_n174), .d(new_n180), .o1(new_n196));
  aoib12aa1n02x5               g101(.a(new_n196), .b(new_n169), .c(new_n187), .out0(new_n197));
  aoi022aa1n02x5               g102(.a(new_n193), .b(new_n194), .c(new_n189), .d(new_n197), .o1(\s[17] ));
  inv040aa1d32x5               g103(.a(\a[17] ), .o1(new_n199));
  inv040aa1d28x5               g104(.a(\b[16] ), .o1(new_n200));
  nand42aa1n02x5               g105(.a(new_n200), .b(new_n199), .o1(new_n201));
  oabi12aa1n06x5               g106(.a(new_n191), .b(new_n157), .c(new_n187), .out0(new_n202));
  aoai13aa1n03x5               g107(.a(new_n194), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n203));
  nor002aa1n03x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nand02aa1d08x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  norb02aa1n06x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n203), .c(new_n201), .out0(\s[18] ));
  and002aa1n02x5               g112(.a(new_n194), .b(new_n206), .o(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n209));
  aoi013aa1n09x5               g114(.a(new_n204), .b(new_n205), .c(new_n199), .d(new_n200), .o1(new_n210));
  nor002aa1d32x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand42aa1n16x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n12x5               g120(.a(\a[18] ), .b(\b[17] ), .c(new_n201), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n213), .b(new_n216), .c(new_n193), .d(new_n208), .o1(new_n217));
  nor002aa1d32x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanp02aa1n12x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  inv000aa1d42x5               g125(.a(\a[19] ), .o1(new_n221));
  inv000aa1d42x5               g126(.a(\b[18] ), .o1(new_n222));
  aboi22aa1n03x5               g127(.a(new_n218), .b(new_n219), .c(new_n221), .d(new_n222), .out0(new_n223));
  inv000aa1n06x5               g128(.a(new_n211), .o1(new_n224));
  inv000aa1d42x5               g129(.a(new_n213), .o1(new_n225));
  aoai13aa1n02x7               g130(.a(new_n224), .b(new_n225), .c(new_n209), .d(new_n210), .o1(new_n226));
  aoi022aa1n02x7               g131(.a(new_n226), .b(new_n220), .c(new_n217), .d(new_n223), .o1(\s[20] ));
  nano23aa1n06x5               g132(.a(new_n211), .b(new_n218), .c(new_n219), .d(new_n212), .out0(new_n228));
  nand23aa1n06x5               g133(.a(new_n228), .b(new_n194), .c(new_n206), .o1(new_n229));
  tech160nm_fiaoi012aa1n05x5   g134(.a(new_n229), .b(new_n189), .c(new_n192), .o1(new_n230));
  nona23aa1n09x5               g135(.a(new_n219), .b(new_n212), .c(new_n211), .d(new_n218), .out0(new_n231));
  oaoi03aa1n09x5               g136(.a(\a[20] ), .b(\b[19] ), .c(new_n224), .o1(new_n232));
  inv040aa1n03x5               g137(.a(new_n232), .o1(new_n233));
  oai012aa1d24x5               g138(.a(new_n233), .b(new_n231), .c(new_n210), .o1(new_n234));
  tech160nm_fixnrc02aa1n05x5   g139(.a(\b[20] ), .b(\a[21] ), .out0(new_n235));
  oabi12aa1n03x5               g140(.a(new_n235), .b(new_n230), .c(new_n234), .out0(new_n236));
  oai112aa1n02x5               g141(.a(new_n233), .b(new_n235), .c(new_n231), .d(new_n210), .o1(new_n237));
  oa0012aa1n03x5               g142(.a(new_n236), .b(new_n230), .c(new_n237), .o(\s[21] ));
  xnrc02aa1n12x5               g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nor042aa1n03x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n239), .b(new_n241), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n229), .o1(new_n243));
  aoai13aa1n02x5               g148(.a(new_n243), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n234), .o1(new_n245));
  inv000aa1n03x5               g150(.a(new_n241), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n235), .c(new_n244), .d(new_n245), .o1(new_n247));
  aoi022aa1n03x5               g152(.a(new_n247), .b(new_n240), .c(new_n236), .d(new_n242), .o1(\s[22] ));
  nor042aa1n06x5               g153(.a(new_n239), .b(new_n235), .o1(new_n249));
  norb02aa1n03x5               g154(.a(new_n249), .b(new_n229), .out0(new_n250));
  aoai13aa1n03x5               g155(.a(new_n250), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n251));
  oao003aa1n02x5               g156(.a(\a[22] ), .b(\b[21] ), .c(new_n246), .carry(new_n252));
  inv000aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  aoi012aa1n02x5               g158(.a(new_n253), .b(new_n234), .c(new_n249), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n254), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n255), .c(new_n193), .d(new_n250), .o1(new_n257));
  aoi112aa1n02x5               g162(.a(new_n256), .b(new_n253), .c(new_n234), .d(new_n249), .o1(new_n258));
  aobi12aa1n02x7               g163(.a(new_n257), .b(new_n258), .c(new_n251), .out0(\s[23] ));
  tech160nm_fixorc02aa1n04x5   g164(.a(\a[24] ), .b(\b[23] ), .out0(new_n260));
  nor042aa1n06x5               g165(.a(\b[22] ), .b(\a[23] ), .o1(new_n261));
  norp02aa1n02x5               g166(.a(new_n260), .b(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n261), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n256), .o1(new_n264));
  aoai13aa1n02x7               g169(.a(new_n263), .b(new_n264), .c(new_n251), .d(new_n254), .o1(new_n265));
  aoi022aa1n02x7               g170(.a(new_n265), .b(new_n260), .c(new_n257), .d(new_n262), .o1(\s[24] ));
  nano32aa1n03x7               g171(.a(new_n229), .b(new_n260), .c(new_n249), .d(new_n256), .out0(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n268));
  aoai13aa1n09x5               g173(.a(new_n249), .b(new_n232), .c(new_n228), .d(new_n216), .o1(new_n269));
  and002aa1n06x5               g174(.a(new_n260), .b(new_n256), .o(new_n270));
  inv020aa1n04x5               g175(.a(new_n270), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[24] ), .b(\b[23] ), .c(new_n263), .carry(new_n272));
  aoai13aa1n12x5               g177(.a(new_n272), .b(new_n271), .c(new_n269), .d(new_n252), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n193), .d(new_n267), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n270), .b(new_n253), .c(new_n234), .d(new_n249), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n274), .o1(new_n277));
  and003aa1n02x5               g182(.a(new_n276), .b(new_n277), .c(new_n272), .o(new_n278));
  aobi12aa1n02x7               g183(.a(new_n275), .b(new_n278), .c(new_n268), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g184(.a(\a[26] ), .b(\b[25] ), .out0(new_n280));
  norp02aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .o1(new_n281));
  norp02aa1n02x5               g186(.a(new_n280), .b(new_n281), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n273), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n281), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n277), .c(new_n268), .d(new_n283), .o1(new_n285));
  aoi022aa1n02x7               g190(.a(new_n285), .b(new_n280), .c(new_n275), .d(new_n282), .o1(\s[26] ));
  and002aa1n12x5               g191(.a(new_n280), .b(new_n274), .o(new_n287));
  inv000aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nano23aa1n06x5               g193(.a(new_n288), .b(new_n229), .c(new_n270), .d(new_n249), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n202), .c(new_n134), .d(new_n188), .o1(new_n290));
  nanp02aa1n02x5               g195(.a(\b[25] ), .b(\a[26] ), .o1(new_n291));
  oai022aa1n02x5               g196(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n292));
  nanp02aa1n02x5               g197(.a(new_n292), .b(new_n291), .o1(new_n293));
  aoai13aa1n04x5               g198(.a(new_n293), .b(new_n288), .c(new_n276), .d(new_n272), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n193), .d(new_n289), .o1(new_n296));
  aoi122aa1n02x7               g201(.a(new_n295), .b(new_n291), .c(new_n292), .d(new_n273), .e(new_n287), .o1(new_n297));
  aobi12aa1n02x7               g202(.a(new_n296), .b(new_n297), .c(new_n290), .out0(\s[27] ));
  xorc02aa1n02x5               g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  nor042aa1d18x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  norp02aa1n02x5               g205(.a(new_n299), .b(new_n300), .o1(new_n301));
  aoi022aa1n09x5               g206(.a(new_n273), .b(new_n287), .c(new_n291), .d(new_n292), .o1(new_n302));
  inv040aa1n08x5               g207(.a(new_n300), .o1(new_n303));
  inv000aa1n02x5               g208(.a(new_n295), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n303), .b(new_n304), .c(new_n302), .d(new_n290), .o1(new_n305));
  aoi022aa1n02x7               g210(.a(new_n305), .b(new_n299), .c(new_n296), .d(new_n301), .o1(\s[28] ));
  and002aa1n02x5               g211(.a(new_n299), .b(new_n295), .o(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n294), .c(new_n193), .d(new_n289), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n307), .o1(new_n309));
  oao003aa1n09x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n303), .carry(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n309), .c(new_n302), .d(new_n290), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n308), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g220(.a(new_n304), .b(new_n299), .c(new_n312), .out0(new_n316));
  aoai13aa1n02x5               g221(.a(new_n316), .b(new_n294), .c(new_n193), .d(new_n289), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n316), .o1(new_n318));
  tech160nm_fioaoi03aa1n03p5x5 g223(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n319), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n318), .c(new_n302), .d(new_n290), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  and002aa1n02x5               g227(.a(\b[28] ), .b(\a[29] ), .o(new_n323));
  oabi12aa1n02x5               g228(.a(new_n322), .b(\a[29] ), .c(\b[28] ), .out0(new_n324));
  oab012aa1n02x4               g229(.a(new_n324), .b(new_n310), .c(new_n323), .out0(new_n325));
  aoi022aa1n03x5               g230(.a(new_n321), .b(new_n322), .c(new_n317), .d(new_n325), .o1(\s[30] ));
  nano32aa1n03x7               g231(.a(new_n304), .b(new_n322), .c(new_n299), .d(new_n312), .out0(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n294), .c(new_n193), .d(new_n289), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  inv000aa1d42x5               g234(.a(\a[30] ), .o1(new_n330));
  inv000aa1d42x5               g235(.a(\b[29] ), .o1(new_n331));
  oabi12aa1n02x5               g236(.a(new_n329), .b(\a[30] ), .c(\b[29] ), .out0(new_n332));
  oaoi13aa1n02x5               g237(.a(new_n332), .b(new_n319), .c(new_n330), .d(new_n331), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n327), .o1(new_n334));
  oaoi03aa1n02x5               g239(.a(new_n330), .b(new_n331), .c(new_n319), .o1(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n334), .c(new_n302), .d(new_n290), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n336), .b(new_n329), .c(new_n328), .d(new_n333), .o1(\s[31] ));
  nanp03aa1n02x5               g242(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n338));
  xnbna2aa1n03x5               g243(.a(new_n106), .b(new_n338), .c(new_n101), .out0(\s[3] ));
  nanp02aa1n02x5               g244(.a(new_n104), .b(new_n106), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n105), .b(new_n340), .c(new_n109), .out0(\s[4] ));
  xnbna2aa1n03x5               g246(.a(new_n116), .b(new_n107), .c(new_n110), .out0(\s[5] ));
  aoai13aa1n02x5               g247(.a(new_n114), .b(new_n122), .c(new_n111), .d(new_n116), .o1(new_n343));
  aoi112aa1n02x5               g248(.a(new_n122), .b(new_n114), .c(new_n111), .d(new_n116), .o1(new_n344));
  norb02aa1n02x5               g249(.a(new_n343), .b(new_n344), .out0(\s[6] ));
  xnbna2aa1n03x5               g250(.a(new_n118), .b(new_n343), .c(new_n121), .out0(\s[7] ));
  aob012aa1n02x5               g251(.a(new_n118), .b(new_n343), .c(new_n121), .out0(new_n347));
  aoai13aa1n02x5               g252(.a(new_n124), .b(new_n132), .c(new_n343), .d(new_n121), .o1(new_n348));
  norb02aa1n02x5               g253(.a(new_n124), .b(new_n117), .out0(new_n349));
  aoi022aa1n02x5               g254(.a(new_n348), .b(new_n117), .c(new_n347), .d(new_n349), .o1(\s[8] ));
  nanp02aa1n02x5               g255(.a(new_n111), .b(new_n120), .o1(new_n351));
  aoi113aa1n02x5               g256(.a(new_n128), .b(new_n125), .c(new_n123), .d(new_n118), .e(new_n117), .o1(new_n352));
  aoi022aa1n02x5               g257(.a(new_n134), .b(new_n128), .c(new_n351), .d(new_n352), .o1(\s[9] ));
endmodule


