// Benchmark "adder" written by ABC on Wed Jul 17 19:27:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n367, new_n368, new_n370, new_n371, new_n372, new_n373, new_n375,
    new_n376, new_n378, new_n380, new_n381, new_n382, new_n384, new_n385,
    new_n386;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n09x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  nanb02aa1n12x5               g004(.a(\b[1] ), .b(new_n99), .out0(new_n100));
  nand42aa1n08x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n12x5               g006(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(new_n102));
  nor042aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  tech160nm_finand02aa1n03p5x5 g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  norb02aa1n06x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  inv000aa1n04x5               g010(.a(new_n105), .o1(new_n106));
  nor002aa1n03x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  norb03aa1n03x5               g013(.a(new_n108), .b(new_n103), .c(new_n107), .out0(new_n109));
  aoai13aa1n06x5               g014(.a(new_n109), .b(new_n106), .c(new_n100), .d(new_n102), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand02aa1d08x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand23aa1n02x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .o1(new_n114));
  tech160nm_fioai012aa1n04x5   g019(.a(new_n108), .b(\b[6] ), .c(\a[7] ), .o1(new_n115));
  nor002aa1n12x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  orn002aa1n24x5               g021(.a(\a[6] ), .b(\b[5] ), .o(new_n117));
  nor002aa1n06x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nand42aa1n06x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nona23aa1n03x5               g024(.a(new_n119), .b(new_n117), .c(new_n116), .d(new_n118), .out0(new_n120));
  nor043aa1n02x5               g025(.a(new_n120), .b(new_n115), .c(new_n114), .o1(new_n121));
  nor042aa1n02x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  oai012aa1n02x5               g027(.a(new_n113), .b(new_n118), .c(new_n122), .o1(new_n123));
  oai112aa1n06x5               g028(.a(new_n117), .b(new_n119), .c(\b[4] ), .d(\a[5] ), .o1(new_n124));
  aoi022aa1n12x5               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  nona23aa1n09x5               g030(.a(new_n125), .b(new_n113), .c(new_n122), .d(new_n118), .out0(new_n126));
  oaib12aa1n09x5               g031(.a(new_n123), .b(new_n126), .c(new_n124), .out0(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n03x5               g033(.a(new_n128), .b(new_n127), .c(new_n110), .d(new_n121), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[10] ), .b(\b[9] ), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  nand02aa1n03x5               g036(.a(new_n102), .b(new_n100), .o1(new_n132));
  nona22aa1n03x5               g037(.a(new_n108), .b(new_n107), .c(new_n103), .out0(new_n133));
  aoi012aa1n12x5               g038(.a(new_n133), .b(new_n132), .c(new_n105), .o1(new_n134));
  oai022aa1n03x5               g039(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n135));
  aoi112aa1n03x5               g040(.a(new_n135), .b(new_n118), .c(\a[6] ), .d(\b[5] ), .o1(new_n136));
  nona22aa1n09x5               g041(.a(new_n136), .b(new_n114), .c(new_n115), .out0(new_n137));
  oai022aa1n02x5               g042(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n138));
  aoai13aa1n12x5               g043(.a(new_n113), .b(new_n138), .c(new_n124), .d(new_n125), .o1(new_n139));
  oai012aa1d24x5               g044(.a(new_n139), .b(new_n134), .c(new_n137), .o1(new_n140));
  aoai13aa1n06x5               g045(.a(new_n130), .b(new_n97), .c(new_n140), .d(new_n128), .o1(new_n141));
  tech160nm_fioaoi03aa1n02p5x5 g046(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n142));
  inv000aa1d42x5               g047(.a(new_n142), .o1(new_n143));
  nor002aa1n04x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nand42aa1n16x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  norb02aa1n02x7               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n141), .c(new_n143), .out0(\s[11] ));
  nanp02aa1n03x5               g052(.a(new_n129), .b(new_n98), .o1(new_n148));
  aoai13aa1n03x5               g053(.a(new_n146), .b(new_n142), .c(new_n148), .d(new_n130), .o1(new_n149));
  inv040aa1d32x5               g054(.a(\a[11] ), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\b[10] ), .o1(new_n151));
  nanp02aa1n04x5               g056(.a(new_n151), .b(new_n150), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n146), .o1(new_n153));
  aoai13aa1n02x5               g058(.a(new_n152), .b(new_n153), .c(new_n141), .d(new_n143), .o1(new_n154));
  nor002aa1n20x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand42aa1n10x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  aboi22aa1n03x5               g062(.a(new_n155), .b(new_n156), .c(new_n150), .d(new_n151), .out0(new_n158));
  aoi022aa1n03x5               g063(.a(new_n154), .b(new_n157), .c(new_n149), .d(new_n158), .o1(\s[12] ));
  nano23aa1d15x5               g064(.a(new_n144), .b(new_n155), .c(new_n156), .d(new_n145), .out0(new_n160));
  nand23aa1d12x5               g065(.a(new_n160), .b(new_n128), .c(new_n130), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n127), .c(new_n110), .d(new_n121), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(\b[9] ), .b(\a[10] ), .o1(new_n164));
  oai022aa1n02x5               g069(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n165));
  nanb03aa1n02x5               g070(.a(new_n155), .b(new_n156), .c(new_n145), .out0(new_n166));
  nano32aa1n03x7               g071(.a(new_n166), .b(new_n165), .c(new_n152), .d(new_n164), .out0(new_n167));
  oaoi03aa1n12x5               g072(.a(\a[12] ), .b(\b[11] ), .c(new_n152), .o1(new_n168));
  norp02aa1n02x5               g073(.a(new_n167), .b(new_n168), .o1(new_n169));
  nanp02aa1n03x5               g074(.a(new_n163), .b(new_n169), .o1(new_n170));
  nor002aa1d32x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nand42aa1n06x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  norb02aa1n03x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  norp03aa1n02x5               g078(.a(new_n167), .b(new_n168), .c(new_n173), .o1(new_n174));
  aoi022aa1n02x5               g079(.a(new_n170), .b(new_n173), .c(new_n163), .d(new_n174), .o1(\s[13] ));
  orn002aa1n02x5               g080(.a(\a[13] ), .b(\b[12] ), .o(new_n176));
  inv000aa1n02x5               g081(.a(new_n169), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n173), .b(new_n177), .c(new_n140), .d(new_n162), .o1(new_n178));
  nor002aa1d32x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nand42aa1n06x5               g084(.a(\b[13] ), .b(\a[14] ), .o1(new_n180));
  norb02aa1n06x4               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n178), .c(new_n176), .out0(\s[14] ));
  nona23aa1d24x5               g087(.a(new_n180), .b(new_n172), .c(new_n171), .d(new_n179), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  aoai13aa1n06x5               g089(.a(new_n184), .b(new_n177), .c(new_n140), .d(new_n162), .o1(new_n185));
  oaoi03aa1n12x5               g090(.a(\a[14] ), .b(\b[13] ), .c(new_n176), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  nor002aa1n16x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  nand42aa1n04x5               g093(.a(\b[14] ), .b(\a[15] ), .o1(new_n189));
  norb02aa1n15x5               g094(.a(new_n189), .b(new_n188), .out0(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n190), .b(new_n185), .c(new_n187), .out0(\s[15] ));
  aoai13aa1n03x5               g096(.a(new_n190), .b(new_n186), .c(new_n170), .d(new_n184), .o1(new_n192));
  inv040aa1n02x5               g097(.a(new_n188), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n190), .o1(new_n194));
  aoai13aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n185), .d(new_n187), .o1(new_n195));
  nor042aa1d18x5               g100(.a(\b[15] ), .b(\a[16] ), .o1(new_n196));
  nand02aa1n06x5               g101(.a(\b[15] ), .b(\a[16] ), .o1(new_n197));
  norb02aa1n06x5               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n196), .o1(new_n199));
  aoi012aa1n02x5               g104(.a(new_n188), .b(new_n199), .c(new_n197), .o1(new_n200));
  aoi022aa1n03x5               g105(.a(new_n195), .b(new_n198), .c(new_n192), .d(new_n200), .o1(\s[16] ));
  nano23aa1n06x5               g106(.a(new_n188), .b(new_n196), .c(new_n197), .d(new_n189), .out0(new_n202));
  nano32aa1d12x5               g107(.a(new_n161), .b(new_n202), .c(new_n173), .d(new_n181), .out0(new_n203));
  nanp02aa1n02x5               g108(.a(new_n140), .b(new_n203), .o1(new_n204));
  aoi012aa1n09x5               g109(.a(new_n127), .b(new_n110), .c(new_n121), .o1(new_n205));
  nano22aa1n12x5               g110(.a(new_n183), .b(new_n190), .c(new_n198), .out0(new_n206));
  nanb02aa1n03x5               g111(.a(new_n161), .b(new_n206), .out0(new_n207));
  oai012aa1n12x5               g112(.a(new_n206), .b(new_n167), .c(new_n168), .o1(new_n208));
  aoi022aa1d24x5               g113(.a(\b[14] ), .b(\a[15] ), .c(\a[14] ), .d(\b[13] ), .o1(new_n209));
  oai012aa1n06x5               g114(.a(new_n209), .b(new_n179), .c(new_n171), .o1(new_n210));
  nand02aa1n04x5               g115(.a(new_n210), .b(new_n193), .o1(new_n211));
  aoi012aa1d18x5               g116(.a(new_n196), .b(new_n211), .c(new_n197), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  norb02aa1n06x5               g118(.a(new_n208), .b(new_n213), .out0(new_n214));
  oai012aa1n12x5               g119(.a(new_n214), .b(new_n205), .c(new_n207), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[17] ), .b(\b[16] ), .out0(new_n216));
  nanp02aa1n02x5               g121(.a(new_n211), .b(new_n197), .o1(new_n217));
  nano32aa1n02x4               g122(.a(new_n216), .b(new_n208), .c(new_n217), .d(new_n199), .out0(new_n218));
  aoi022aa1n02x5               g123(.a(new_n215), .b(new_n216), .c(new_n218), .d(new_n204), .o1(\s[17] ));
  nor042aa1d18x5               g124(.a(\b[16] ), .b(\a[17] ), .o1(new_n220));
  inv000aa1n02x5               g125(.a(new_n220), .o1(new_n221));
  nand22aa1n12x5               g126(.a(new_n208), .b(new_n212), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n216), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n223));
  nor042aa1d18x5               g128(.a(\b[17] ), .b(\a[18] ), .o1(new_n224));
  nand42aa1n06x5               g129(.a(\b[17] ), .b(\a[18] ), .o1(new_n225));
  norb02aa1n02x5               g130(.a(new_n225), .b(new_n224), .out0(new_n226));
  xnbna2aa1n03x5               g131(.a(new_n226), .b(new_n223), .c(new_n221), .out0(\s[18] ));
  nand42aa1n02x5               g132(.a(\b[16] ), .b(\a[17] ), .o1(new_n228));
  nano23aa1n06x5               g133(.a(new_n220), .b(new_n224), .c(new_n225), .d(new_n228), .out0(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n230));
  oaoi03aa1n02x5               g135(.a(\a[18] ), .b(\b[17] ), .c(new_n221), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  xorc02aa1n12x5               g137(.a(\a[19] ), .b(\b[18] ), .out0(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n230), .c(new_n232), .out0(\s[19] ));
  xnrc02aa1n02x5               g139(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g140(.a(new_n233), .b(new_n231), .c(new_n215), .d(new_n229), .o1(new_n236));
  nor002aa1d32x5               g141(.a(\b[18] ), .b(\a[19] ), .o1(new_n237));
  inv030aa1n06x5               g142(.a(new_n237), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n233), .o1(new_n239));
  aoai13aa1n02x5               g144(.a(new_n238), .b(new_n239), .c(new_n230), .d(new_n232), .o1(new_n240));
  norp02aa1n24x5               g145(.a(\b[19] ), .b(\a[20] ), .o1(new_n241));
  nand42aa1n10x5               g146(.a(\b[19] ), .b(\a[20] ), .o1(new_n242));
  norb02aa1n06x5               g147(.a(new_n242), .b(new_n241), .out0(new_n243));
  inv000aa1d42x5               g148(.a(\a[19] ), .o1(new_n244));
  inv000aa1d42x5               g149(.a(\b[18] ), .o1(new_n245));
  aboi22aa1n03x5               g150(.a(new_n241), .b(new_n242), .c(new_n244), .d(new_n245), .out0(new_n246));
  aoi022aa1n03x5               g151(.a(new_n240), .b(new_n243), .c(new_n236), .d(new_n246), .o1(\s[20] ));
  nand23aa1d12x5               g152(.a(new_n229), .b(new_n233), .c(new_n243), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n12x5               g154(.a(new_n249), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n250));
  tech160nm_finand02aa1n03p5x5 g155(.a(\b[18] ), .b(\a[19] ), .o1(new_n251));
  nanb03aa1n12x5               g156(.a(new_n241), .b(new_n242), .c(new_n251), .out0(new_n252));
  oai112aa1n06x5               g157(.a(new_n238), .b(new_n225), .c(new_n224), .d(new_n220), .o1(new_n253));
  aoi012aa1d24x5               g158(.a(new_n241), .b(new_n237), .c(new_n242), .o1(new_n254));
  oai012aa1d24x5               g159(.a(new_n254), .b(new_n253), .c(new_n252), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  nand42aa1n06x5               g161(.a(new_n250), .b(new_n256), .o1(new_n257));
  nor002aa1d32x5               g162(.a(\b[20] ), .b(\a[21] ), .o1(new_n258));
  nanp02aa1n04x5               g163(.a(\b[20] ), .b(\a[21] ), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n259), .b(new_n258), .out0(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  oai112aa1n02x5               g166(.a(new_n254), .b(new_n261), .c(new_n253), .d(new_n252), .o1(new_n262));
  aboi22aa1n03x5               g167(.a(new_n262), .b(new_n250), .c(new_n257), .d(new_n260), .out0(\s[21] ));
  nand02aa1n02x5               g168(.a(new_n257), .b(new_n260), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n258), .o1(new_n265));
  aoai13aa1n04x5               g170(.a(new_n265), .b(new_n261), .c(new_n250), .d(new_n256), .o1(new_n266));
  nor022aa1n12x5               g171(.a(\b[21] ), .b(\a[22] ), .o1(new_n267));
  nand22aa1n12x5               g172(.a(\b[21] ), .b(\a[22] ), .o1(new_n268));
  norb02aa1n02x5               g173(.a(new_n268), .b(new_n267), .out0(new_n269));
  aoib12aa1n02x5               g174(.a(new_n258), .b(new_n268), .c(new_n267), .out0(new_n270));
  aoi022aa1n03x5               g175(.a(new_n266), .b(new_n269), .c(new_n264), .d(new_n270), .o1(\s[22] ));
  nona23aa1d16x5               g176(.a(new_n268), .b(new_n259), .c(new_n258), .d(new_n267), .out0(new_n272));
  nano32aa1n02x4               g177(.a(new_n272), .b(new_n229), .c(new_n233), .d(new_n243), .out0(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n272), .o1(new_n275));
  aoi012aa1n02x5               g180(.a(new_n267), .b(new_n258), .c(new_n268), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n276), .o1(new_n277));
  aoi012aa1n02x5               g182(.a(new_n277), .b(new_n255), .c(new_n275), .o1(new_n278));
  nand42aa1n02x5               g183(.a(new_n274), .b(new_n278), .o1(new_n279));
  nor042aa1n12x5               g184(.a(\b[22] ), .b(\a[23] ), .o1(new_n280));
  nand02aa1n03x5               g185(.a(\b[22] ), .b(\a[23] ), .o1(new_n281));
  norb02aa1d21x5               g186(.a(new_n281), .b(new_n280), .out0(new_n282));
  aoi112aa1n02x5               g187(.a(new_n282), .b(new_n277), .c(new_n255), .d(new_n275), .o1(new_n283));
  aoi022aa1n02x5               g188(.a(new_n279), .b(new_n282), .c(new_n274), .d(new_n283), .o1(\s[23] ));
  nanp02aa1n03x5               g189(.a(new_n279), .b(new_n282), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n280), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n282), .o1(new_n287));
  aoai13aa1n02x7               g192(.a(new_n286), .b(new_n287), .c(new_n274), .d(new_n278), .o1(new_n288));
  norp02aa1n06x5               g193(.a(\b[23] ), .b(\a[24] ), .o1(new_n289));
  nand42aa1n03x5               g194(.a(\b[23] ), .b(\a[24] ), .o1(new_n290));
  norb02aa1n06x4               g195(.a(new_n290), .b(new_n289), .out0(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n280), .o1(new_n292));
  aoi022aa1n03x5               g197(.a(new_n288), .b(new_n291), .c(new_n285), .d(new_n292), .o1(\s[24] ));
  nano22aa1d15x5               g198(.a(new_n272), .b(new_n282), .c(new_n291), .out0(new_n294));
  norb02aa1n06x4               g199(.a(new_n294), .b(new_n248), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n296));
  aoai13aa1n02x7               g201(.a(new_n281), .b(new_n267), .c(new_n258), .d(new_n268), .o1(new_n297));
  aoi022aa1n06x5               g202(.a(new_n297), .b(new_n286), .c(\a[24] ), .d(\b[23] ), .o1(new_n298));
  aoi112aa1n09x5               g203(.a(new_n289), .b(new_n298), .c(new_n255), .d(new_n294), .o1(new_n299));
  nand42aa1n04x5               g204(.a(new_n296), .b(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[25] ), .b(\b[24] ), .out0(new_n301));
  nand02aa1d04x5               g206(.a(new_n255), .b(new_n294), .o1(new_n302));
  nona32aa1n02x4               g207(.a(new_n302), .b(new_n298), .c(new_n301), .d(new_n289), .out0(new_n303));
  aboi22aa1n03x5               g208(.a(new_n303), .b(new_n296), .c(new_n300), .d(new_n301), .out0(\s[25] ));
  nand02aa1n02x5               g209(.a(new_n300), .b(new_n301), .o1(new_n305));
  nor042aa1n03x5               g210(.a(\b[24] ), .b(\a[25] ), .o1(new_n306));
  inv040aa1n03x5               g211(.a(new_n306), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n301), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n307), .b(new_n308), .c(new_n296), .d(new_n299), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[26] ), .b(\b[25] ), .out0(new_n310));
  norp02aa1n02x5               g215(.a(new_n310), .b(new_n306), .o1(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n305), .d(new_n311), .o1(\s[26] ));
  and002aa1n12x5               g217(.a(new_n310), .b(new_n301), .o(new_n313));
  nano22aa1d15x5               g218(.a(new_n248), .b(new_n313), .c(new_n294), .out0(new_n314));
  aoai13aa1n12x5               g219(.a(new_n314), .b(new_n222), .c(new_n140), .d(new_n203), .o1(new_n315));
  nona22aa1n03x5               g220(.a(new_n302), .b(new_n298), .c(new_n289), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[26] ), .b(\b[25] ), .c(new_n307), .carry(new_n317));
  inv000aa1n02x5               g222(.a(new_n317), .o1(new_n318));
  tech160nm_fiaoi012aa1n05x5   g223(.a(new_n318), .b(new_n316), .c(new_n313), .o1(new_n319));
  nanp02aa1n02x5               g224(.a(new_n319), .b(new_n315), .o1(new_n320));
  xorc02aa1n12x5               g225(.a(\a[27] ), .b(\b[26] ), .out0(new_n321));
  aoi112aa1n02x5               g226(.a(new_n321), .b(new_n318), .c(new_n316), .d(new_n313), .o1(new_n322));
  aoi022aa1n02x5               g227(.a(new_n320), .b(new_n321), .c(new_n315), .d(new_n322), .o1(\s[27] ));
  oaib12aa1n12x5               g228(.a(new_n317), .b(new_n299), .c(new_n313), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n321), .b(new_n324), .c(new_n215), .d(new_n314), .o1(new_n325));
  norp02aa1n02x5               g230(.a(\b[26] ), .b(\a[27] ), .o1(new_n326));
  inv000aa1n03x5               g231(.a(new_n326), .o1(new_n327));
  inv000aa1d42x5               g232(.a(new_n321), .o1(new_n328));
  aoai13aa1n02x7               g233(.a(new_n327), .b(new_n328), .c(new_n319), .d(new_n315), .o1(new_n329));
  tech160nm_fixorc02aa1n03p5x5 g234(.a(\a[28] ), .b(\b[27] ), .out0(new_n330));
  norp02aa1n02x5               g235(.a(new_n330), .b(new_n326), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n329), .b(new_n330), .c(new_n325), .d(new_n331), .o1(\s[28] ));
  and002aa1n06x5               g237(.a(new_n330), .b(new_n321), .o(new_n333));
  aoai13aa1n03x5               g238(.a(new_n333), .b(new_n324), .c(new_n215), .d(new_n314), .o1(new_n334));
  inv000aa1d42x5               g239(.a(new_n333), .o1(new_n335));
  oao003aa1n02x5               g240(.a(\a[28] ), .b(\b[27] ), .c(new_n327), .carry(new_n336));
  aoai13aa1n02x7               g241(.a(new_n336), .b(new_n335), .c(new_n319), .d(new_n315), .o1(new_n337));
  tech160nm_fixorc02aa1n03p5x5 g242(.a(\a[29] ), .b(\b[28] ), .out0(new_n338));
  norb02aa1n02x5               g243(.a(new_n336), .b(new_n338), .out0(new_n339));
  aoi022aa1n03x5               g244(.a(new_n337), .b(new_n338), .c(new_n334), .d(new_n339), .o1(\s[29] ));
  xorb03aa1n02x5               g245(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d33x5               g246(.a(new_n328), .b(new_n330), .c(new_n338), .out0(new_n342));
  aoai13aa1n03x5               g247(.a(new_n342), .b(new_n324), .c(new_n215), .d(new_n314), .o1(new_n343));
  inv000aa1d42x5               g248(.a(new_n342), .o1(new_n344));
  inv000aa1d42x5               g249(.a(\b[28] ), .o1(new_n345));
  inv000aa1d42x5               g250(.a(\a[29] ), .o1(new_n346));
  oaib12aa1n02x5               g251(.a(new_n336), .b(\b[28] ), .c(new_n346), .out0(new_n347));
  oaib12aa1n02x5               g252(.a(new_n347), .b(new_n345), .c(\a[29] ), .out0(new_n348));
  aoai13aa1n02x7               g253(.a(new_n348), .b(new_n344), .c(new_n319), .d(new_n315), .o1(new_n349));
  xorc02aa1n02x5               g254(.a(\a[30] ), .b(\b[29] ), .out0(new_n350));
  oaoi13aa1n02x5               g255(.a(new_n350), .b(new_n347), .c(new_n346), .d(new_n345), .o1(new_n351));
  aoi022aa1n03x5               g256(.a(new_n349), .b(new_n350), .c(new_n343), .d(new_n351), .o1(\s[30] ));
  nanb02aa1n02x5               g257(.a(\b[30] ), .b(\a[31] ), .out0(new_n353));
  nanb02aa1n02x5               g258(.a(\a[31] ), .b(\b[30] ), .out0(new_n354));
  nanp02aa1n02x5               g259(.a(new_n354), .b(new_n353), .o1(new_n355));
  nano32aa1n03x7               g260(.a(new_n328), .b(new_n350), .c(new_n330), .d(new_n338), .out0(new_n356));
  aoai13aa1n03x5               g261(.a(new_n356), .b(new_n324), .c(new_n215), .d(new_n314), .o1(new_n357));
  inv000aa1d42x5               g262(.a(new_n356), .o1(new_n358));
  norp02aa1n02x5               g263(.a(\b[29] ), .b(\a[30] ), .o1(new_n359));
  aoi022aa1n02x5               g264(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n360));
  aoi012aa1n02x5               g265(.a(new_n359), .b(new_n347), .c(new_n360), .o1(new_n361));
  aoai13aa1n02x7               g266(.a(new_n361), .b(new_n358), .c(new_n319), .d(new_n315), .o1(new_n362));
  oai112aa1n02x5               g267(.a(new_n353), .b(new_n354), .c(\b[29] ), .d(\a[30] ), .o1(new_n363));
  aoi012aa1n02x5               g268(.a(new_n363), .b(new_n347), .c(new_n360), .o1(new_n364));
  aoi022aa1n03x5               g269(.a(new_n362), .b(new_n355), .c(new_n357), .d(new_n364), .o1(\s[31] ));
  xnbna2aa1n03x5               g270(.a(new_n105), .b(new_n102), .c(new_n100), .out0(\s[3] ));
  norb02aa1n02x5               g271(.a(new_n108), .b(new_n107), .out0(new_n367));
  aoi012aa1n02x5               g272(.a(new_n103), .b(new_n132), .c(new_n105), .o1(new_n368));
  oai012aa1n02x5               g273(.a(new_n110), .b(new_n368), .c(new_n367), .o1(\s[4] ));
  inv000aa1d42x5               g274(.a(new_n116), .o1(new_n370));
  aoi022aa1n02x5               g275(.a(new_n110), .b(new_n108), .c(new_n370), .d(new_n111), .o1(new_n371));
  nano22aa1n02x4               g276(.a(new_n116), .b(new_n108), .c(new_n111), .out0(new_n372));
  aoai13aa1n02x5               g277(.a(new_n372), .b(new_n133), .c(new_n132), .d(new_n105), .o1(new_n373));
  norb02aa1n02x5               g278(.a(new_n373), .b(new_n371), .out0(\s[5] ));
  xorc02aa1n02x5               g279(.a(\a[6] ), .b(\b[5] ), .out0(new_n375));
  nanb02aa1n02x5               g280(.a(new_n124), .b(new_n373), .out0(new_n376));
  aoai13aa1n02x5               g281(.a(new_n376), .b(new_n375), .c(new_n370), .d(new_n373), .o1(\s[6] ));
  norb02aa1n02x5               g282(.a(new_n112), .b(new_n122), .out0(new_n378));
  xobna2aa1n03x5               g283(.a(new_n378), .b(new_n376), .c(new_n119), .out0(\s[7] ));
  aoi013aa1n02x4               g284(.a(new_n122), .b(new_n376), .c(new_n378), .d(new_n119), .o1(new_n380));
  norb02aa1n02x5               g285(.a(new_n113), .b(new_n118), .out0(new_n381));
  aoi113aa1n02x5               g286(.a(new_n381), .b(new_n122), .c(new_n376), .d(new_n378), .e(new_n119), .o1(new_n382));
  aoib12aa1n02x5               g287(.a(new_n382), .b(new_n381), .c(new_n380), .out0(\s[8] ));
  nanp02aa1n02x5               g288(.a(new_n121), .b(new_n110), .o1(new_n384));
  nanb02aa1n02x5               g289(.a(new_n128), .b(new_n123), .out0(new_n385));
  aoib12aa1n02x5               g290(.a(new_n385), .b(new_n124), .c(new_n126), .out0(new_n386));
  aoi022aa1n02x5               g291(.a(new_n140), .b(new_n128), .c(new_n384), .d(new_n386), .o1(\s[9] ));
endmodule


