// Benchmark "adder" written by ABC on Wed Jul 17 18:11:21 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n311, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n331, new_n333, new_n334, new_n336, new_n337, new_n339, new_n341,
    new_n343;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nor042aa1n06x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nand02aa1d28x5               g005(.a(\b[7] ), .b(\a[8] ), .o1(new_n101));
  nor042aa1n06x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nand02aa1d20x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nano23aa1n06x5               g008(.a(new_n100), .b(new_n102), .c(new_n103), .d(new_n101), .out0(new_n104));
  nona23aa1d18x5               g009(.a(new_n103), .b(new_n101), .c(new_n100), .d(new_n102), .out0(new_n105));
  oai022aa1d24x5               g010(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n106));
  aob012aa1d15x5               g011(.a(new_n106), .b(\b[5] ), .c(\a[6] ), .out0(new_n107));
  oa0012aa1n03x5               g012(.a(new_n101), .b(new_n102), .c(new_n100), .o(new_n108));
  oabi12aa1n06x5               g013(.a(new_n108), .b(new_n105), .c(new_n107), .out0(new_n109));
  oai022aa1d18x5               g014(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n110));
  nor002aa1n06x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nand42aa1d28x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  norb02aa1n06x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nor022aa1n06x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  aoi022aa1d24x5               g019(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n115));
  tech160nm_fioai012aa1n05x5   g020(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n116));
  tech160nm_fixorc02aa1n04x5   g021(.a(\a[6] ), .b(\b[5] ), .out0(new_n117));
  and002aa1n02x5               g022(.a(\b[4] ), .b(\a[5] ), .o(new_n118));
  nanp02aa1n09x5               g023(.a(\b[3] ), .b(\a[4] ), .o1(new_n119));
  oai012aa1n06x5               g024(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .o1(new_n120));
  nor042aa1n03x5               g025(.a(new_n120), .b(new_n118), .o1(new_n121));
  nanp02aa1n09x5               g026(.a(new_n121), .b(new_n117), .o1(new_n122));
  aoib12aa1n06x5               g027(.a(new_n122), .b(new_n116), .c(new_n110), .out0(new_n123));
  xnrc02aa1n12x5               g028(.a(\b[8] ), .b(\a[9] ), .out0(new_n124));
  inv000aa1d42x5               g029(.a(new_n124), .o1(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n109), .c(new_n123), .d(new_n104), .o1(new_n126));
  nor002aa1d32x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n16x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n15x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  aob012aa1n03x5               g035(.a(new_n129), .b(new_n126), .c(new_n99), .out0(new_n131));
  aoai13aa1n12x5               g036(.a(new_n128), .b(new_n127), .c(new_n97), .d(new_n98), .o1(new_n132));
  xorc02aa1n12x5               g037(.a(\a[11] ), .b(\b[10] ), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n133), .b(new_n131), .c(new_n132), .out0(\s[11] ));
  inv000aa1d42x5               g039(.a(new_n129), .o1(new_n135));
  aoai13aa1n04x5               g040(.a(new_n132), .b(new_n135), .c(new_n126), .d(new_n99), .o1(new_n136));
  inv040aa1d28x5               g041(.a(\a[11] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(\b[10] ), .o1(new_n138));
  nand02aa1n08x5               g043(.a(new_n138), .b(new_n137), .o1(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  orn002aa1n24x5               g045(.a(\a[12] ), .b(\b[11] ), .o(new_n141));
  nand02aa1n08x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nanp02aa1n06x5               g047(.a(new_n141), .b(new_n142), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n140), .c(new_n136), .d(new_n133), .o1(new_n144));
  aoi112aa1n02x7               g049(.a(new_n140), .b(new_n143), .c(new_n136), .d(new_n133), .o1(new_n145));
  nanb02aa1n03x5               g050(.a(new_n145), .b(new_n144), .out0(\s[12] ));
  nona23aa1d18x5               g051(.a(new_n129), .b(new_n133), .c(new_n124), .d(new_n143), .out0(new_n147));
  inv040aa1n03x5               g052(.a(new_n147), .o1(new_n148));
  aoai13aa1n06x5               g053(.a(new_n148), .b(new_n109), .c(new_n123), .d(new_n104), .o1(new_n149));
  and002aa1n02x5               g054(.a(\b[10] ), .b(\a[11] ), .o(new_n150));
  aoai13aa1n12x5               g055(.a(new_n141), .b(new_n150), .c(new_n132), .d(new_n139), .o1(new_n151));
  nand42aa1n03x5               g056(.a(new_n151), .b(new_n142), .o1(new_n152));
  nor002aa1n12x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanp02aa1n04x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  xnbna2aa1n03x5               g060(.a(new_n155), .b(new_n149), .c(new_n152), .out0(\s[13] ));
  inv000aa1d42x5               g061(.a(\a[13] ), .o1(new_n157));
  inv000aa1d42x5               g062(.a(\b[12] ), .o1(new_n158));
  aoib12aa1n06x5               g063(.a(new_n108), .b(new_n104), .c(new_n107), .out0(new_n159));
  oaoi13aa1n12x5               g064(.a(new_n110), .b(new_n113), .c(new_n115), .d(new_n114), .o1(new_n160));
  inv000aa1n02x5               g065(.a(new_n160), .o1(new_n161));
  nona22aa1n03x5               g066(.a(new_n161), .b(new_n122), .c(new_n105), .out0(new_n162));
  aoai13aa1n02x5               g067(.a(new_n152), .b(new_n147), .c(new_n162), .d(new_n159), .o1(new_n163));
  oaoi03aa1n03x5               g068(.a(new_n157), .b(new_n158), .c(new_n163), .o1(new_n164));
  xnrb03aa1n03x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n24x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nand22aa1n09x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nona23aa1d18x5               g072(.a(new_n167), .b(new_n154), .c(new_n153), .d(new_n166), .out0(new_n168));
  aoai13aa1n06x5               g073(.a(new_n167), .b(new_n166), .c(new_n157), .d(new_n158), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n168), .c(new_n149), .d(new_n152), .o1(new_n170));
  nor042aa1n06x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nand22aa1n09x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  oai022aa1d18x5               g078(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n174));
  aboi22aa1n03x5               g079(.a(new_n171), .b(new_n172), .c(new_n174), .d(new_n167), .out0(new_n175));
  aoai13aa1n02x5               g080(.a(new_n175), .b(new_n168), .c(new_n149), .d(new_n152), .o1(new_n176));
  aobi12aa1n02x5               g081(.a(new_n176), .b(new_n173), .c(new_n170), .out0(\s[15] ));
  nor042aa1n04x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nand02aa1n03x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  aoai13aa1n03x5               g085(.a(new_n180), .b(new_n171), .c(new_n170), .d(new_n172), .o1(new_n181));
  aoi112aa1n03x5               g086(.a(new_n171), .b(new_n180), .c(new_n170), .d(new_n172), .o1(new_n182));
  nanb02aa1n03x5               g087(.a(new_n182), .b(new_n181), .out0(\s[16] ));
  oai013aa1d12x5               g088(.a(new_n159), .b(new_n160), .c(new_n122), .d(new_n105), .o1(new_n184));
  nona23aa1n09x5               g089(.a(new_n179), .b(new_n172), .c(new_n171), .d(new_n178), .out0(new_n185));
  nor042aa1n09x5               g090(.a(new_n185), .b(new_n168), .o1(new_n186));
  norb02aa1d21x5               g091(.a(new_n186), .b(new_n147), .out0(new_n187));
  nand22aa1n12x5               g092(.a(new_n184), .b(new_n187), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n172), .b(new_n171), .c(new_n174), .d(new_n167), .o1(new_n189));
  oaoi03aa1n03x5               g094(.a(\a[16] ), .b(\b[15] ), .c(new_n189), .o1(new_n190));
  aoi013aa1n09x5               g095(.a(new_n190), .b(new_n151), .c(new_n186), .d(new_n142), .o1(new_n191));
  nand02aa1d10x5               g096(.a(new_n188), .b(new_n191), .o1(new_n192));
  xorc02aa1n12x5               g097(.a(\a[17] ), .b(\b[16] ), .out0(new_n193));
  aoi113aa1n02x5               g098(.a(new_n193), .b(new_n190), .c(new_n151), .d(new_n186), .e(new_n142), .o1(new_n194));
  aoi022aa1n02x5               g099(.a(new_n192), .b(new_n193), .c(new_n188), .d(new_n194), .o1(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[17] ), .o1(new_n196));
  inv000aa1d42x5               g101(.a(\b[16] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  nanp03aa1n03x5               g103(.a(new_n151), .b(new_n186), .c(new_n142), .o1(new_n199));
  oaoi03aa1n02x5               g104(.a(\a[15] ), .b(\b[14] ), .c(new_n169), .o1(new_n200));
  oai012aa1n02x7               g105(.a(new_n179), .b(new_n200), .c(new_n178), .o1(new_n201));
  nand02aa1d04x5               g106(.a(new_n199), .b(new_n201), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n193), .b(new_n202), .c(new_n184), .d(new_n187), .o1(new_n203));
  nor002aa1n03x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  nand42aa1n06x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  nanb02aa1n18x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  xobna2aa1n03x5               g111(.a(new_n206), .b(new_n203), .c(new_n198), .out0(\s[18] ));
  norb02aa1n02x5               g112(.a(new_n193), .b(new_n206), .out0(new_n208));
  aoai13aa1n06x5               g113(.a(new_n208), .b(new_n202), .c(new_n184), .d(new_n187), .o1(new_n209));
  aoai13aa1n12x5               g114(.a(new_n205), .b(new_n204), .c(new_n196), .d(new_n197), .o1(new_n210));
  nor002aa1n10x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand22aa1n04x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n03x5               g120(.a(new_n209), .b(new_n210), .o1(new_n216));
  nor022aa1n08x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1d28x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  aoai13aa1n02x5               g124(.a(new_n219), .b(new_n211), .c(new_n216), .d(new_n213), .o1(new_n220));
  oaoi03aa1n03x5               g125(.a(\a[18] ), .b(\b[17] ), .c(new_n198), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n213), .b(new_n221), .c(new_n192), .d(new_n208), .o1(new_n222));
  nona22aa1n03x5               g127(.a(new_n222), .b(new_n219), .c(new_n211), .out0(new_n223));
  nanp02aa1n03x5               g128(.a(new_n220), .b(new_n223), .o1(\s[20] ));
  nona23aa1d18x5               g129(.a(new_n218), .b(new_n212), .c(new_n211), .d(new_n217), .out0(new_n225));
  ao0012aa1n12x5               g130(.a(new_n217), .b(new_n211), .c(new_n218), .o(new_n226));
  oabi12aa1n18x5               g131(.a(new_n226), .b(new_n225), .c(new_n210), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  norb03aa1n12x5               g133(.a(new_n193), .b(new_n225), .c(new_n206), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n12x5               g135(.a(new_n228), .b(new_n230), .c(new_n188), .d(new_n191), .o1(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoi012aa1n03x5               g138(.a(new_n233), .b(new_n192), .c(new_n229), .o1(new_n234));
  aoi022aa1n02x5               g139(.a(new_n234), .b(new_n228), .c(new_n231), .d(new_n233), .o1(\s[21] ));
  nor042aa1n03x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[21] ), .b(\a[22] ), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n236), .c(new_n231), .d(new_n233), .o1(new_n238));
  nand02aa1n02x5               g143(.a(new_n231), .b(new_n233), .o1(new_n239));
  nona22aa1n03x5               g144(.a(new_n239), .b(new_n237), .c(new_n236), .out0(new_n240));
  nanp02aa1n03x5               g145(.a(new_n240), .b(new_n238), .o1(\s[22] ));
  nor042aa1n06x5               g146(.a(new_n237), .b(new_n232), .o1(new_n242));
  nona23aa1n09x5               g147(.a(new_n242), .b(new_n193), .c(new_n225), .d(new_n206), .out0(new_n243));
  nano23aa1n06x5               g148(.a(new_n211), .b(new_n217), .c(new_n218), .d(new_n212), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n242), .b(new_n226), .c(new_n244), .d(new_n221), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oaoi03aa1n12x5               g152(.a(new_n246), .b(new_n247), .c(new_n236), .o1(new_n248));
  nanp02aa1n02x5               g153(.a(new_n245), .b(new_n248), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n250), .b(new_n243), .c(new_n188), .d(new_n191), .o1(new_n251));
  xorc02aa1n12x5               g156(.a(\a[23] ), .b(\b[22] ), .out0(new_n252));
  nanp02aa1n03x5               g157(.a(new_n251), .b(new_n252), .o1(new_n253));
  aoi113aa1n03x5               g158(.a(new_n249), .b(new_n252), .c(new_n192), .d(new_n229), .e(new_n242), .o1(new_n254));
  norb02aa1n02x7               g159(.a(new_n253), .b(new_n254), .out0(\s[23] ));
  norp02aa1n02x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  tech160nm_fixnrc02aa1n05x5   g161(.a(\b[23] ), .b(\a[24] ), .out0(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n256), .c(new_n251), .d(new_n252), .o1(new_n258));
  nona22aa1n03x5               g163(.a(new_n253), .b(new_n257), .c(new_n256), .out0(new_n259));
  nanp02aa1n03x5               g164(.a(new_n259), .b(new_n258), .o1(\s[24] ));
  norb02aa1n03x5               g165(.a(new_n252), .b(new_n257), .out0(new_n261));
  nand23aa1n03x5               g166(.a(new_n229), .b(new_n242), .c(new_n261), .o1(new_n262));
  inv000aa1n03x5               g167(.a(new_n261), .o1(new_n263));
  orn002aa1n02x5               g168(.a(\a[23] ), .b(\b[22] ), .o(new_n264));
  oao003aa1n02x5               g169(.a(\a[24] ), .b(\b[23] ), .c(new_n264), .carry(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n263), .c(new_n245), .d(new_n248), .o1(new_n266));
  inv040aa1n06x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n12x5               g172(.a(new_n267), .b(new_n262), .c(new_n188), .d(new_n191), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  xorc02aa1n12x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  tech160nm_fixnrc02aa1n05x5   g176(.a(\b[25] ), .b(\a[26] ), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n270), .c(new_n268), .d(new_n271), .o1(new_n273));
  nand42aa1n02x5               g178(.a(new_n268), .b(new_n271), .o1(new_n274));
  nona22aa1n03x5               g179(.a(new_n274), .b(new_n272), .c(new_n270), .out0(new_n275));
  nanp02aa1n03x5               g180(.a(new_n275), .b(new_n273), .o1(\s[26] ));
  norb02aa1n12x5               g181(.a(new_n271), .b(new_n272), .out0(new_n277));
  nano22aa1n03x7               g182(.a(new_n243), .b(new_n261), .c(new_n277), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n202), .c(new_n184), .d(new_n187), .o1(new_n279));
  tech160nm_finand02aa1n05x5   g184(.a(new_n266), .b(new_n277), .o1(new_n280));
  aoi112aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n281));
  oab012aa1n02x4               g186(.a(new_n281), .b(\a[26] ), .c(\b[25] ), .out0(new_n282));
  nanp03aa1n06x5               g187(.a(new_n279), .b(new_n280), .c(new_n282), .o1(new_n283));
  xorc02aa1n12x5               g188(.a(\a[27] ), .b(\b[26] ), .out0(new_n284));
  nano22aa1n02x4               g189(.a(new_n284), .b(new_n280), .c(new_n282), .out0(new_n285));
  aoi022aa1n02x5               g190(.a(new_n285), .b(new_n279), .c(new_n283), .d(new_n284), .o1(\s[27] ));
  nor042aa1n03x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  xnrc02aa1n12x5               g192(.a(\b[27] ), .b(\a[28] ), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n287), .c(new_n283), .d(new_n284), .o1(new_n289));
  aobi12aa1n09x5               g194(.a(new_n278), .b(new_n188), .c(new_n191), .out0(new_n290));
  inv040aa1d30x5               g195(.a(new_n248), .o1(new_n291));
  aoai13aa1n06x5               g196(.a(new_n261), .b(new_n291), .c(new_n227), .d(new_n242), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n277), .o1(new_n293));
  aoai13aa1n04x5               g198(.a(new_n282), .b(new_n293), .c(new_n292), .d(new_n265), .o1(new_n294));
  oaih12aa1n02x5               g199(.a(new_n284), .b(new_n294), .c(new_n290), .o1(new_n295));
  nona22aa1n03x5               g200(.a(new_n295), .b(new_n288), .c(new_n287), .out0(new_n296));
  nanp02aa1n03x5               g201(.a(new_n289), .b(new_n296), .o1(\s[28] ));
  norb02aa1n03x5               g202(.a(new_n284), .b(new_n288), .out0(new_n298));
  oaih12aa1n02x5               g203(.a(new_n298), .b(new_n294), .c(new_n290), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[29] ), .b(\b[28] ), .out0(new_n300));
  inv000aa1d42x5               g205(.a(\a[28] ), .o1(new_n301));
  inv000aa1d42x5               g206(.a(\b[27] ), .o1(new_n302));
  aoi112aa1n02x5               g207(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n303));
  aoi112aa1n02x5               g208(.a(new_n300), .b(new_n303), .c(new_n301), .d(new_n302), .o1(new_n304));
  aobi12aa1n06x5               g209(.a(new_n282), .b(new_n266), .c(new_n277), .out0(new_n305));
  inv000aa1d42x5               g210(.a(new_n298), .o1(new_n306));
  oao003aa1n09x5               g211(.a(new_n301), .b(new_n302), .c(new_n287), .carry(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n306), .c(new_n305), .d(new_n279), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n309), .b(new_n300), .c(new_n299), .d(new_n304), .o1(\s[29] ));
  nanp02aa1n02x5               g215(.a(\b[0] ), .b(\a[1] ), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n311), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g217(.a(new_n288), .b(new_n284), .c(new_n300), .out0(new_n313));
  oaih12aa1n02x5               g218(.a(new_n313), .b(new_n294), .c(new_n290), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[30] ), .b(\b[29] ), .out0(new_n315));
  inv000aa1d42x5               g220(.a(\a[29] ), .o1(new_n316));
  inv000aa1d42x5               g221(.a(\b[28] ), .o1(new_n317));
  oabi12aa1n02x5               g222(.a(new_n315), .b(\a[29] ), .c(\b[28] ), .out0(new_n318));
  oaoi13aa1n02x5               g223(.a(new_n318), .b(new_n307), .c(new_n316), .d(new_n317), .o1(new_n319));
  inv000aa1n02x5               g224(.a(new_n313), .o1(new_n320));
  oaoi03aa1n03x5               g225(.a(new_n316), .b(new_n317), .c(new_n307), .o1(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n320), .c(new_n305), .d(new_n279), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n322), .b(new_n315), .c(new_n314), .d(new_n319), .o1(\s[30] ));
  nand03aa1n02x5               g228(.a(new_n298), .b(new_n300), .c(new_n315), .o1(new_n324));
  oabi12aa1n03x5               g229(.a(new_n324), .b(new_n294), .c(new_n290), .out0(new_n325));
  xorc02aa1n02x5               g230(.a(\a[31] ), .b(\b[30] ), .out0(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n327));
  norb02aa1n02x5               g232(.a(new_n327), .b(new_n326), .out0(new_n328));
  aoai13aa1n02x7               g233(.a(new_n327), .b(new_n324), .c(new_n305), .d(new_n279), .o1(new_n329));
  aoi022aa1n03x5               g234(.a(new_n329), .b(new_n326), .c(new_n325), .d(new_n328), .o1(\s[31] ));
  norp03aa1n02x5               g235(.a(new_n113), .b(new_n114), .c(new_n115), .o1(new_n331));
  norb02aa1n02x5               g236(.a(new_n116), .b(new_n331), .out0(\s[3] ));
  xorc02aa1n02x5               g237(.a(\a[4] ), .b(\b[3] ), .out0(new_n333));
  norp02aa1n02x5               g238(.a(new_n333), .b(new_n111), .o1(new_n334));
  aboi22aa1n03x5               g239(.a(new_n160), .b(new_n333), .c(new_n334), .d(new_n116), .out0(\s[4] ));
  xnrc02aa1n02x5               g240(.a(\b[4] ), .b(\a[5] ), .out0(new_n336));
  oaib12aa1n02x5               g241(.a(new_n119), .b(new_n110), .c(new_n116), .out0(new_n337));
  aoi022aa1n02x5               g242(.a(new_n337), .b(new_n336), .c(new_n161), .d(new_n121), .o1(\s[5] ));
  obai22aa1n02x7               g243(.a(new_n121), .b(new_n160), .c(\a[5] ), .d(\b[4] ), .out0(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oai012aa1n02x5               g245(.a(new_n107), .b(new_n160), .c(new_n122), .o1(new_n341));
  xorb03aa1n02x5               g246(.a(new_n341), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g247(.a(new_n102), .b(new_n341), .c(new_n103), .o1(new_n343));
  xnrb03aa1n02x5               g248(.a(new_n343), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g249(.a(new_n125), .b(new_n162), .c(new_n159), .out0(\s[9] ));
endmodule


