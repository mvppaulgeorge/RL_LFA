// Benchmark "adder" written by ABC on Thu Jul 18 07:13:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n328, new_n331, new_n332, new_n333,
    new_n334, new_n336, new_n337, new_n338, new_n340;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[2] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[1] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  oaoi03aa1n09x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  nand02aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nor022aa1n16x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1n06x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nor022aa1n06x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nona23aa1n09x5               g012(.a(new_n106), .b(new_n104), .c(new_n107), .d(new_n105), .out0(new_n108));
  tech160nm_fiaoi012aa1n03p5x5 g013(.a(new_n107), .b(new_n105), .c(new_n106), .o1(new_n109));
  oai012aa1n09x5               g014(.a(new_n109), .b(new_n108), .c(new_n103), .o1(new_n110));
  tech160nm_fixnrc02aa1n02p5x5 g015(.a(\b[6] ), .b(\a[7] ), .out0(new_n111));
  nor022aa1n16x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand42aa1n03x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  norp02aa1n06x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand02aa1n03x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nona23aa1n02x4               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nor043aa1n02x5               g022(.a(new_n116), .b(new_n117), .c(new_n111), .o1(new_n118));
  and002aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o(new_n119));
  inv000aa1d42x5               g024(.a(new_n112), .o1(new_n120));
  nor002aa1n12x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  oai022aa1n06x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  aoai13aa1n02x5               g027(.a(new_n113), .b(new_n121), .c(new_n122), .d(new_n115), .o1(new_n123));
  tech160nm_fioai012aa1n05x5   g028(.a(new_n120), .b(new_n123), .c(new_n119), .o1(new_n124));
  xorc02aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n03x5               g030(.a(new_n125), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n126));
  nor002aa1n06x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n03x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  nanp02aa1n03x5               g035(.a(new_n126), .b(new_n99), .o1(new_n131));
  aoai13aa1n12x5               g036(.a(new_n128), .b(new_n127), .c(new_n97), .d(new_n98), .o1(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  aoi012aa1n02x5               g038(.a(new_n133), .b(new_n131), .c(new_n129), .o1(new_n134));
  nor002aa1n12x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nand42aa1n10x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  xnbna2aa1n03x5               g042(.a(new_n134), .b(new_n137), .c(new_n136), .out0(\s[11] ));
  nanb02aa1d24x5               g043(.a(new_n135), .b(new_n137), .out0(new_n139));
  inv000aa1d42x5               g044(.a(new_n139), .o1(new_n140));
  aoai13aa1n03x5               g045(.a(new_n140), .b(new_n133), .c(new_n131), .d(new_n129), .o1(new_n141));
  nor002aa1n16x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  nand42aa1n03x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n142), .b(new_n143), .out0(new_n144));
  tech160nm_fiaoi012aa1n04x5   g049(.a(new_n144), .b(new_n141), .c(new_n136), .o1(new_n145));
  nanp03aa1n03x5               g050(.a(new_n141), .b(new_n136), .c(new_n144), .o1(new_n146));
  norb02aa1n03x4               g051(.a(new_n146), .b(new_n145), .out0(\s[12] ));
  nona23aa1n03x5               g052(.a(new_n143), .b(new_n137), .c(new_n135), .d(new_n142), .out0(new_n148));
  nano22aa1n02x5               g053(.a(new_n148), .b(new_n125), .c(new_n129), .out0(new_n149));
  aoai13aa1n03x5               g054(.a(new_n149), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n142), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n135), .b(new_n143), .o1(new_n152));
  nor043aa1n03x5               g057(.a(new_n132), .b(new_n139), .c(new_n144), .o1(new_n153));
  nano22aa1n03x7               g058(.a(new_n153), .b(new_n151), .c(new_n152), .out0(new_n154));
  nor042aa1n06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand42aa1n06x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n150), .c(new_n154), .out0(\s[13] ));
  inv000aa1n06x5               g063(.a(new_n155), .o1(new_n159));
  oao003aa1n02x5               g064(.a(new_n100), .b(new_n101), .c(new_n102), .carry(new_n160));
  nano23aa1n02x4               g065(.a(new_n107), .b(new_n105), .c(new_n104), .d(new_n106), .out0(new_n161));
  aobi12aa1n02x5               g066(.a(new_n109), .b(new_n161), .c(new_n160), .out0(new_n162));
  norb02aa1n02x5               g067(.a(new_n113), .b(new_n112), .out0(new_n163));
  norb02aa1n09x5               g068(.a(new_n115), .b(new_n114), .out0(new_n164));
  nona23aa1n02x4               g069(.a(new_n164), .b(new_n163), .c(new_n117), .d(new_n111), .out0(new_n165));
  oab012aa1n02x4               g070(.a(new_n112), .b(new_n123), .c(new_n119), .out0(new_n166));
  tech160nm_fioai012aa1n03p5x5 g071(.a(new_n166), .b(new_n165), .c(new_n162), .o1(new_n167));
  oai112aa1n06x5               g072(.a(new_n152), .b(new_n151), .c(new_n148), .d(new_n132), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n157), .b(new_n168), .c(new_n167), .d(new_n149), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand42aa1n03x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n169), .c(new_n159), .out0(\s[14] ));
  nona23aa1n02x4               g078(.a(new_n171), .b(new_n156), .c(new_n155), .d(new_n170), .out0(new_n174));
  oaoi03aa1n12x5               g079(.a(\a[14] ), .b(\b[13] ), .c(new_n159), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  aoai13aa1n04x5               g081(.a(new_n176), .b(new_n174), .c(new_n150), .d(new_n154), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n04x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nand42aa1n10x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  norp02aa1n04x5               g085(.a(\b[15] ), .b(\a[16] ), .o1(new_n181));
  nand42aa1n06x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  norb02aa1n02x5               g087(.a(new_n182), .b(new_n181), .out0(new_n183));
  aoai13aa1n02x5               g088(.a(new_n183), .b(new_n179), .c(new_n177), .d(new_n180), .o1(new_n184));
  aoi112aa1n02x5               g089(.a(new_n179), .b(new_n183), .c(new_n177), .d(new_n180), .o1(new_n185));
  norb02aa1n03x4               g090(.a(new_n184), .b(new_n185), .out0(\s[16] ));
  nano23aa1n03x5               g091(.a(new_n135), .b(new_n142), .c(new_n143), .d(new_n137), .out0(new_n187));
  nano23aa1n06x5               g092(.a(new_n155), .b(new_n170), .c(new_n171), .d(new_n156), .out0(new_n188));
  nano23aa1n06x5               g093(.a(new_n179), .b(new_n181), .c(new_n182), .d(new_n180), .out0(new_n189));
  nand42aa1n02x5               g094(.a(new_n189), .b(new_n188), .o1(new_n190));
  nano32aa1n03x7               g095(.a(new_n190), .b(new_n187), .c(new_n129), .d(new_n125), .out0(new_n191));
  aoai13aa1n09x5               g096(.a(new_n191), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n192));
  inv000aa1n02x5               g097(.a(new_n190), .o1(new_n193));
  aoi112aa1n02x5               g098(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n194));
  nanp02aa1n06x5               g099(.a(new_n189), .b(new_n175), .o1(new_n195));
  nona22aa1n03x5               g100(.a(new_n195), .b(new_n194), .c(new_n181), .out0(new_n196));
  aoi012aa1d18x5               g101(.a(new_n196), .b(new_n168), .c(new_n193), .o1(new_n197));
  xorc02aa1n02x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  xnbna2aa1n03x5               g103(.a(new_n198), .b(new_n192), .c(new_n197), .out0(\s[17] ));
  inv040aa1d32x5               g104(.a(\a[18] ), .o1(new_n200));
  nanp02aa1n03x5               g105(.a(new_n192), .b(new_n197), .o1(new_n201));
  norp02aa1n02x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  aoi012aa1n03x5               g107(.a(new_n202), .b(new_n201), .c(new_n198), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[17] ), .c(new_n200), .out0(\s[18] ));
  inv000aa1d42x5               g109(.a(\a[17] ), .o1(new_n205));
  xroi22aa1d06x4               g110(.a(new_n205), .b(\b[16] ), .c(new_n200), .d(\b[17] ), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  nand42aa1n02x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  oai022aa1d24x5               g113(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n209));
  and002aa1n02x5               g114(.a(new_n209), .b(new_n208), .o(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n207), .c(new_n192), .d(new_n197), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n03x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand42aa1n03x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norp02aa1n04x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand42aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n215), .c(new_n212), .d(new_n216), .o1(new_n220));
  aoi112aa1n02x5               g125(.a(new_n215), .b(new_n219), .c(new_n212), .d(new_n216), .o1(new_n221));
  norb02aa1n02x7               g126(.a(new_n220), .b(new_n221), .out0(\s[20] ));
  nanb03aa1n06x5               g127(.a(new_n217), .b(new_n218), .c(new_n216), .out0(new_n223));
  nona22aa1n03x5               g128(.a(new_n206), .b(new_n215), .c(new_n223), .out0(new_n224));
  oai112aa1n06x5               g129(.a(new_n209), .b(new_n208), .c(\b[18] ), .d(\a[19] ), .o1(new_n225));
  tech160nm_fiaoi012aa1n03p5x5 g130(.a(new_n217), .b(new_n215), .c(new_n218), .o1(new_n226));
  oai012aa1n12x5               g131(.a(new_n226), .b(new_n225), .c(new_n223), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n224), .c(new_n192), .d(new_n197), .o1(new_n229));
  xorb03aa1n02x5               g134(.a(new_n229), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[21] ), .b(\a[22] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n231), .c(new_n229), .d(new_n233), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(new_n231), .b(new_n235), .c(new_n229), .d(new_n233), .o1(new_n237));
  norb02aa1n02x7               g142(.a(new_n236), .b(new_n237), .out0(\s[22] ));
  nor042aa1n06x5               g143(.a(new_n234), .b(new_n232), .o1(new_n239));
  nona23aa1n08x5               g144(.a(new_n206), .b(new_n239), .c(new_n223), .d(new_n215), .out0(new_n240));
  nano22aa1n02x4               g145(.a(new_n217), .b(new_n216), .c(new_n218), .out0(new_n241));
  oai012aa1n02x5               g146(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n209), .b(new_n242), .out0(new_n243));
  inv040aa1n03x5               g148(.a(new_n226), .o1(new_n244));
  aoai13aa1n06x5               g149(.a(new_n239), .b(new_n244), .c(new_n243), .d(new_n241), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oao003aa1n12x5               g152(.a(new_n246), .b(new_n247), .c(new_n231), .carry(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  nand02aa1n03x5               g154(.a(new_n245), .b(new_n249), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n240), .c(new_n192), .d(new_n197), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  xorc02aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  aoai13aa1n03x5               g161(.a(new_n256), .b(new_n254), .c(new_n252), .d(new_n255), .o1(new_n257));
  aoi112aa1n02x5               g162(.a(new_n254), .b(new_n256), .c(new_n252), .d(new_n255), .o1(new_n258));
  norb02aa1n03x4               g163(.a(new_n257), .b(new_n258), .out0(\s[24] ));
  nano32aa1n03x7               g164(.a(new_n224), .b(new_n256), .c(new_n239), .d(new_n255), .out0(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  and002aa1n02x5               g166(.a(new_n256), .b(new_n255), .o(new_n262));
  inv000aa1d42x5               g167(.a(\a[24] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(\b[23] ), .o1(new_n264));
  oao003aa1n02x5               g169(.a(new_n263), .b(new_n264), .c(new_n254), .carry(new_n265));
  aoi012aa1n06x5               g170(.a(new_n265), .b(new_n250), .c(new_n262), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n261), .c(new_n192), .d(new_n197), .o1(new_n267));
  xorb03aa1n02x5               g172(.a(new_n267), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  tech160nm_fixorc02aa1n02p5x5 g174(.a(\a[25] ), .b(\b[24] ), .out0(new_n270));
  xorc02aa1n02x5               g175(.a(\a[26] ), .b(\b[25] ), .out0(new_n271));
  aoai13aa1n03x5               g176(.a(new_n271), .b(new_n269), .c(new_n267), .d(new_n270), .o1(new_n272));
  aoi112aa1n02x5               g177(.a(new_n269), .b(new_n271), .c(new_n267), .d(new_n270), .o1(new_n273));
  norb02aa1n03x4               g178(.a(new_n272), .b(new_n273), .out0(\s[26] ));
  oabi12aa1n03x5               g179(.a(new_n196), .b(new_n154), .c(new_n190), .out0(new_n275));
  and002aa1n06x5               g180(.a(new_n271), .b(new_n270), .o(new_n276));
  nano22aa1n03x7               g181(.a(new_n240), .b(new_n262), .c(new_n276), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n275), .c(new_n167), .d(new_n191), .o1(new_n278));
  inv000aa1n02x5               g183(.a(new_n262), .o1(new_n279));
  inv030aa1n02x5               g184(.a(new_n265), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n279), .c(new_n245), .d(new_n249), .o1(new_n281));
  oai022aa1n02x5               g186(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n282));
  aob012aa1n02x5               g187(.a(new_n282), .b(\b[25] ), .c(\a[26] ), .out0(new_n283));
  aobi12aa1n06x5               g188(.a(new_n283), .b(new_n281), .c(new_n276), .out0(new_n284));
  xorc02aa1n02x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n284), .c(new_n278), .out0(\s[27] ));
  norp02aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  inv040aa1n03x5               g192(.a(new_n287), .o1(new_n288));
  nand02aa1n02x5               g193(.a(new_n260), .b(new_n276), .o1(new_n289));
  aoi012aa1n06x5               g194(.a(new_n289), .b(new_n192), .c(new_n197), .o1(new_n290));
  aoai13aa1n02x7               g195(.a(new_n262), .b(new_n248), .c(new_n227), .d(new_n239), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n276), .o1(new_n292));
  aoai13aa1n04x5               g197(.a(new_n283), .b(new_n292), .c(new_n291), .d(new_n280), .o1(new_n293));
  oaih12aa1n02x5               g198(.a(new_n285), .b(new_n293), .c(new_n290), .o1(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  tech160nm_fiaoi012aa1n02p5x5 g200(.a(new_n295), .b(new_n294), .c(new_n288), .o1(new_n296));
  aobi12aa1n02x7               g201(.a(new_n285), .b(new_n284), .c(new_n278), .out0(new_n297));
  nano22aa1n03x5               g202(.a(new_n297), .b(new_n288), .c(new_n295), .out0(new_n298));
  norp02aa1n03x5               g203(.a(new_n296), .b(new_n298), .o1(\s[28] ));
  norb02aa1n02x5               g204(.a(new_n285), .b(new_n295), .out0(new_n300));
  oaih12aa1n02x5               g205(.a(new_n300), .b(new_n293), .c(new_n290), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[28] ), .b(\b[27] ), .c(new_n288), .carry(new_n302));
  xnrc02aa1n02x5               g207(.a(\b[28] ), .b(\a[29] ), .out0(new_n303));
  tech160nm_fiaoi012aa1n02p5x5 g208(.a(new_n303), .b(new_n301), .c(new_n302), .o1(new_n304));
  aobi12aa1n02x7               g209(.a(new_n300), .b(new_n284), .c(new_n278), .out0(new_n305));
  nano22aa1n03x5               g210(.a(new_n305), .b(new_n302), .c(new_n303), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n304), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g213(.a(new_n285), .b(new_n303), .c(new_n295), .out0(new_n309));
  oaih12aa1n02x5               g214(.a(new_n309), .b(new_n293), .c(new_n290), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n302), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .out0(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n312), .b(new_n310), .c(new_n311), .o1(new_n313));
  aobi12aa1n02x7               g218(.a(new_n309), .b(new_n284), .c(new_n278), .out0(new_n314));
  nano22aa1n03x5               g219(.a(new_n314), .b(new_n311), .c(new_n312), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n313), .b(new_n315), .o1(\s[30] ));
  norb02aa1n02x5               g221(.a(new_n309), .b(new_n312), .out0(new_n317));
  aobi12aa1n02x7               g222(.a(new_n317), .b(new_n284), .c(new_n278), .out0(new_n318));
  oao003aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n319));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n320), .out0(new_n321));
  oaih12aa1n02x5               g226(.a(new_n317), .b(new_n293), .c(new_n290), .o1(new_n322));
  tech160nm_fiaoi012aa1n02p5x5 g227(.a(new_n320), .b(new_n322), .c(new_n319), .o1(new_n323));
  norp02aa1n03x5               g228(.a(new_n323), .b(new_n321), .o1(\s[31] ));
  xnrb03aa1n02x5               g229(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanb02aa1n02x5               g230(.a(new_n107), .b(new_n106), .out0(new_n326));
  oai112aa1n02x5               g231(.a(new_n326), .b(new_n104), .c(new_n160), .d(new_n105), .o1(new_n327));
  oabi12aa1n02x5               g232(.a(new_n105), .b(new_n108), .c(new_n103), .out0(new_n328));
  oai012aa1n02x5               g233(.a(new_n327), .b(new_n328), .c(new_n326), .o1(\s[4] ));
  xorb03aa1n02x5               g234(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g235(.a(new_n164), .o1(new_n331));
  nanb02aa1n06x5               g236(.a(new_n117), .b(new_n110), .out0(new_n332));
  oaoi13aa1n06x5               g237(.a(new_n331), .b(new_n332), .c(\a[5] ), .d(\b[4] ), .o1(new_n333));
  oai112aa1n02x5               g238(.a(new_n332), .b(new_n331), .c(\b[4] ), .d(\a[5] ), .o1(new_n334));
  norb02aa1n02x5               g239(.a(new_n334), .b(new_n333), .out0(\s[6] ));
  and002aa1n02x5               g240(.a(new_n122), .b(new_n115), .o(new_n336));
  oabi12aa1n06x5               g241(.a(new_n111), .b(new_n333), .c(new_n336), .out0(new_n337));
  norb03aa1n02x5               g242(.a(new_n111), .b(new_n333), .c(new_n336), .out0(new_n338));
  norb02aa1n02x5               g243(.a(new_n337), .b(new_n338), .out0(\s[7] ));
  inv000aa1d42x5               g244(.a(new_n121), .o1(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n163), .b(new_n337), .c(new_n340), .out0(\s[8] ));
  xorb03aa1n02x5               g246(.a(new_n167), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


