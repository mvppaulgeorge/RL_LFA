// Benchmark "adder" written by ABC on Wed Jul 17 19:46:04 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n310, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n331,
    new_n332, new_n334, new_n335, new_n336, new_n338, new_n339, new_n341,
    new_n342, new_n343;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  nor002aa1n16x5               g002(.a(\b[2] ), .b(\a[3] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  nanb02aa1n12x5               g004(.a(new_n98), .b(new_n99), .out0(new_n100));
  nanp02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai112aa1n06x5               g006(.a(\a[1] ), .b(\b[0] ), .c(\b[1] ), .d(\a[2] ), .o1(new_n102));
  nand02aa1d08x5               g007(.a(new_n102), .b(new_n101), .o1(new_n103));
  and002aa1n02x7               g008(.a(\b[3] ), .b(\a[4] ), .o(new_n104));
  nor002aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor043aa1n06x5               g010(.a(new_n104), .b(new_n105), .c(new_n98), .o1(new_n106));
  oai012aa1d24x5               g011(.a(new_n106), .b(new_n103), .c(new_n100), .o1(new_n107));
  nand42aa1n20x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nor022aa1n12x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n12x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb03aa1n03x5               g015(.a(new_n109), .b(new_n110), .c(new_n108), .out0(new_n111));
  tech160nm_fixnrc02aa1n02p5x5 g016(.a(\b[7] ), .b(\a[8] ), .out0(new_n112));
  aoi022aa1d24x5               g017(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  oai122aa1n06x5               g018(.a(new_n113), .b(\a[6] ), .c(\b[5] ), .d(\a[5] ), .e(\b[4] ), .o1(new_n114));
  nor043aa1n06x5               g019(.a(new_n114), .b(new_n111), .c(new_n112), .o1(new_n115));
  nano22aa1n03x7               g020(.a(new_n109), .b(new_n108), .c(new_n110), .out0(new_n116));
  xorc02aa1n12x5               g021(.a(\a[8] ), .b(\b[7] ), .out0(new_n117));
  nor022aa1n04x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  orn002aa1n24x5               g023(.a(\a[5] ), .b(\b[4] ), .o(new_n119));
  nanb03aa1d18x5               g024(.a(new_n118), .b(new_n119), .c(new_n108), .out0(new_n120));
  nanp03aa1n03x5               g025(.a(new_n120), .b(new_n116), .c(new_n117), .o1(new_n121));
  orn002aa1n03x5               g026(.a(\a[7] ), .b(\b[6] ), .o(new_n122));
  oaoi03aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  nanb02aa1n06x5               g028(.a(new_n123), .b(new_n121), .out0(new_n124));
  xorc02aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n107), .d(new_n115), .o1(new_n126));
  xorc02aa1n02x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  and002aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  oai022aa1d24x5               g033(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n129));
  nor042aa1n09x5               g034(.a(new_n129), .b(new_n128), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(new_n126), .b(new_n130), .o1(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n127), .c(new_n97), .d(new_n126), .o1(\s[10] ));
  inv000aa1d42x5               g037(.a(new_n129), .o1(new_n133));
  aoi022aa1n09x5               g038(.a(new_n126), .b(new_n133), .c(\b[9] ), .d(\a[10] ), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  xorc02aa1n02x5               g041(.a(\a[11] ), .b(\b[10] ), .out0(new_n137));
  nor002aa1d32x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1d28x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n15x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n136), .c(new_n134), .d(new_n137), .o1(new_n142));
  aoi112aa1n03x5               g047(.a(new_n141), .b(new_n136), .c(new_n134), .d(new_n137), .o1(new_n143));
  nanb02aa1n03x5               g048(.a(new_n143), .b(new_n142), .out0(\s[12] ));
  nand22aa1n12x5               g049(.a(new_n115), .b(new_n107), .o1(new_n145));
  aoi013aa1n09x5               g050(.a(new_n123), .b(new_n120), .c(new_n116), .d(new_n117), .o1(new_n146));
  aoi022aa1d24x5               g051(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n147));
  norb02aa1n03x5               g052(.a(new_n147), .b(new_n136), .out0(new_n148));
  tech160nm_fiaoi012aa1n05x5   g053(.a(new_n129), .b(\a[9] ), .c(\b[8] ), .o1(new_n149));
  nand23aa1n03x5               g054(.a(new_n148), .b(new_n140), .c(new_n149), .o1(new_n150));
  nona23aa1d18x5               g055(.a(new_n147), .b(new_n139), .c(new_n136), .d(new_n138), .out0(new_n151));
  aoi012aa1d24x5               g056(.a(new_n138), .b(new_n136), .c(new_n139), .o1(new_n152));
  oai012aa1d24x5               g057(.a(new_n152), .b(new_n151), .c(new_n130), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n150), .c(new_n145), .d(new_n146), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nand02aa1n04x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  aoi012aa1n03x5               g063(.a(new_n157), .b(new_n155), .c(new_n158), .o1(new_n159));
  xnrb03aa1n03x5               g064(.a(new_n159), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand02aa1d06x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nano23aa1n06x5               g067(.a(new_n157), .b(new_n161), .c(new_n162), .d(new_n158), .out0(new_n163));
  nanp02aa1n02x5               g068(.a(new_n155), .b(new_n163), .o1(new_n164));
  aoi012aa1n06x5               g069(.a(new_n161), .b(new_n157), .c(new_n162), .o1(new_n165));
  nor002aa1d32x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nand02aa1n04x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n164), .c(new_n165), .out0(\s[15] ));
  nanp02aa1n02x5               g075(.a(new_n164), .b(new_n165), .o1(new_n171));
  nor002aa1d32x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand02aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  aoai13aa1n03x5               g079(.a(new_n174), .b(new_n166), .c(new_n171), .d(new_n169), .o1(new_n175));
  inv020aa1n03x5               g080(.a(new_n165), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n169), .b(new_n176), .c(new_n155), .d(new_n163), .o1(new_n177));
  nona22aa1n02x4               g082(.a(new_n177), .b(new_n174), .c(new_n166), .out0(new_n178));
  nanp02aa1n02x5               g083(.a(new_n175), .b(new_n178), .o1(\s[16] ));
  nona23aa1n09x5               g084(.a(new_n173), .b(new_n167), .c(new_n166), .d(new_n172), .out0(new_n180));
  nona23aa1n09x5               g085(.a(new_n163), .b(new_n149), .c(new_n180), .d(new_n151), .out0(new_n181));
  norb02aa1n02x5               g086(.a(new_n158), .b(new_n157), .out0(new_n182));
  orn002aa1n02x5               g087(.a(\a[14] ), .b(\b[13] ), .o(new_n183));
  nano32aa1n03x7               g088(.a(new_n180), .b(new_n182), .c(new_n183), .d(new_n162), .out0(new_n184));
  oai012aa1n02x7               g089(.a(new_n173), .b(new_n172), .c(new_n166), .o1(new_n185));
  oai012aa1n12x5               g090(.a(new_n185), .b(new_n180), .c(new_n165), .o1(new_n186));
  aoi012aa1d24x5               g091(.a(new_n186), .b(new_n153), .c(new_n184), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n181), .c(new_n145), .d(new_n146), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1d18x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nand42aa1d28x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  tech160nm_fiaoi012aa1n05x5   g096(.a(new_n190), .b(new_n188), .c(new_n191), .o1(new_n192));
  xnrb03aa1n03x5               g097(.a(new_n192), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nand02aa1d08x5               g098(.a(new_n145), .b(new_n146), .o1(new_n194));
  nano23aa1n06x5               g099(.a(new_n166), .b(new_n172), .c(new_n173), .d(new_n167), .out0(new_n195));
  nand02aa1n03x5               g100(.a(new_n195), .b(new_n163), .o1(new_n196));
  nor042aa1n06x5               g101(.a(new_n150), .b(new_n196), .o1(new_n197));
  oai112aa1n02x5               g102(.a(new_n148), .b(new_n140), .c(new_n129), .d(new_n128), .o1(new_n198));
  aobi12aa1n06x5               g103(.a(new_n185), .b(new_n195), .c(new_n176), .out0(new_n199));
  aoai13aa1n06x5               g104(.a(new_n199), .b(new_n196), .c(new_n198), .d(new_n152), .o1(new_n200));
  nor002aa1n16x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand42aa1d28x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nano23aa1d15x5               g107(.a(new_n190), .b(new_n201), .c(new_n202), .d(new_n191), .out0(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n200), .c(new_n194), .d(new_n197), .o1(new_n204));
  aoi012aa1d24x5               g109(.a(new_n201), .b(new_n190), .c(new_n202), .o1(new_n205));
  xorc02aa1n12x5               g110(.a(\a[19] ), .b(\b[18] ), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n204), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g113(.a(new_n204), .b(new_n205), .o1(new_n209));
  norp02aa1n02x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  xnrc02aa1n12x5               g115(.a(\b[19] ), .b(\a[20] ), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n210), .c(new_n209), .d(new_n206), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n205), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n206), .b(new_n213), .c(new_n188), .d(new_n203), .o1(new_n214));
  nona22aa1n03x5               g119(.a(new_n214), .b(new_n211), .c(new_n210), .out0(new_n215));
  nanp02aa1n03x5               g120(.a(new_n212), .b(new_n215), .o1(\s[20] ));
  aoai13aa1n06x5               g121(.a(new_n197), .b(new_n124), .c(new_n107), .d(new_n115), .o1(new_n217));
  xorc02aa1n03x5               g122(.a(\a[20] ), .b(\b[19] ), .out0(new_n218));
  nand23aa1n06x5               g123(.a(new_n203), .b(new_n206), .c(new_n218), .o1(new_n219));
  xnrc02aa1n12x5               g124(.a(\b[18] ), .b(\a[19] ), .out0(new_n220));
  orn002aa1n03x5               g125(.a(\a[19] ), .b(\b[18] ), .o(new_n221));
  oao003aa1n03x5               g126(.a(\a[20] ), .b(\b[19] ), .c(new_n221), .carry(new_n222));
  oai013aa1d12x5               g127(.a(new_n222), .b(new_n220), .c(new_n211), .d(new_n205), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n219), .c(new_n217), .d(new_n187), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  nand42aa1d28x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  norb02aa1n06x5               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  nor002aa1n16x5               g134(.a(\b[21] ), .b(\a[22] ), .o1(new_n230));
  nand42aa1d28x5               g135(.a(\b[21] ), .b(\a[22] ), .o1(new_n231));
  norb02aa1n12x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n03x5               g138(.a(new_n233), .b(new_n227), .c(new_n225), .d(new_n229), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n219), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n229), .b(new_n223), .c(new_n188), .d(new_n235), .o1(new_n236));
  nona22aa1n03x5               g141(.a(new_n236), .b(new_n233), .c(new_n227), .out0(new_n237));
  nanp02aa1n03x5               g142(.a(new_n234), .b(new_n237), .o1(\s[22] ));
  nano23aa1d12x5               g143(.a(new_n227), .b(new_n230), .c(new_n231), .d(new_n228), .out0(new_n239));
  nona23aa1d18x5               g144(.a(new_n203), .b(new_n239), .c(new_n211), .d(new_n220), .out0(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n200), .c(new_n194), .d(new_n197), .o1(new_n242));
  aoi012aa1n06x5               g147(.a(new_n230), .b(new_n227), .c(new_n231), .o1(new_n243));
  aobi12aa1n02x7               g148(.a(new_n243), .b(new_n223), .c(new_n239), .out0(new_n244));
  xorc02aa1n12x5               g149(.a(\a[23] ), .b(\b[22] ), .out0(new_n245));
  xnbna2aa1n03x5               g150(.a(new_n245), .b(new_n242), .c(new_n244), .out0(\s[23] ));
  aoai13aa1n04x5               g151(.a(new_n244), .b(new_n240), .c(new_n217), .d(new_n187), .o1(new_n247));
  nor002aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  xnrc02aa1n12x5               g153(.a(\b[23] ), .b(\a[24] ), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n248), .c(new_n247), .d(new_n245), .o1(new_n250));
  nanp02aa1n02x5               g155(.a(new_n247), .b(new_n245), .o1(new_n251));
  nona22aa1n02x4               g156(.a(new_n251), .b(new_n249), .c(new_n248), .out0(new_n252));
  nanp02aa1n03x5               g157(.a(new_n252), .b(new_n250), .o1(\s[24] ));
  xorc02aa1n12x5               g158(.a(\a[24] ), .b(\b[23] ), .out0(new_n254));
  nano32aa1n03x7               g159(.a(new_n219), .b(new_n254), .c(new_n239), .d(new_n245), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n200), .c(new_n194), .d(new_n197), .o1(new_n256));
  tech160nm_fixnrc02aa1n03p5x5 g161(.a(\b[22] ), .b(\a[23] ), .out0(new_n257));
  nano23aa1n09x5               g162(.a(new_n249), .b(new_n257), .c(new_n232), .d(new_n229), .out0(new_n258));
  nor002aa1n02x5               g163(.a(\b[23] ), .b(\a[24] ), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  aob012aa1n02x5               g165(.a(new_n248), .b(\b[23] ), .c(\a[24] ), .out0(new_n261));
  nanb03aa1n03x5               g166(.a(new_n243), .b(new_n254), .c(new_n245), .out0(new_n262));
  nand23aa1n06x5               g167(.a(new_n262), .b(new_n260), .c(new_n261), .o1(new_n263));
  aoi012aa1d24x5               g168(.a(new_n263), .b(new_n223), .c(new_n258), .o1(new_n264));
  nand42aa1n04x5               g169(.a(new_n256), .b(new_n264), .o1(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  aoi112aa1n02x5               g171(.a(new_n263), .b(new_n266), .c(new_n223), .d(new_n258), .o1(new_n267));
  aoi022aa1n02x5               g172(.a(new_n265), .b(new_n266), .c(new_n256), .d(new_n267), .o1(\s[25] ));
  nor002aa1n02x5               g173(.a(\b[24] ), .b(\a[25] ), .o1(new_n269));
  xnrc02aa1n12x5               g174(.a(\b[25] ), .b(\a[26] ), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n265), .d(new_n266), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n264), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n266), .b(new_n272), .c(new_n188), .d(new_n255), .o1(new_n273));
  nona22aa1n03x5               g178(.a(new_n273), .b(new_n270), .c(new_n269), .out0(new_n274));
  nanp02aa1n02x5               g179(.a(new_n271), .b(new_n274), .o1(\s[26] ));
  norb02aa1n15x5               g180(.a(new_n266), .b(new_n270), .out0(new_n276));
  nano32aa1d12x5               g181(.a(new_n240), .b(new_n276), .c(new_n245), .d(new_n254), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n200), .c(new_n194), .d(new_n197), .o1(new_n278));
  nanb03aa1n03x5               g183(.a(new_n205), .b(new_n218), .c(new_n206), .out0(new_n279));
  nanp03aa1n02x5               g184(.a(new_n239), .b(new_n245), .c(new_n254), .o1(new_n280));
  tech160nm_fiaoi012aa1n04x5   g185(.a(new_n280), .b(new_n279), .c(new_n222), .o1(new_n281));
  inv000aa1d42x5               g186(.a(\a[26] ), .o1(new_n282));
  inv000aa1d42x5               g187(.a(\b[25] ), .o1(new_n283));
  oao003aa1n02x5               g188(.a(new_n282), .b(new_n283), .c(new_n269), .carry(new_n284));
  oaoi13aa1n09x5               g189(.a(new_n284), .b(new_n276), .c(new_n281), .d(new_n263), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n278), .c(new_n285), .out0(\s[27] ));
  nand02aa1n03x5               g192(.a(new_n278), .b(new_n285), .o1(new_n288));
  norp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  xorc02aa1n12x5               g194(.a(\a[28] ), .b(\b[27] ), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n289), .c(new_n288), .d(new_n286), .o1(new_n292));
  nand02aa1d04x5               g197(.a(new_n223), .b(new_n258), .o1(new_n293));
  norp03aa1n02x5               g198(.a(new_n249), .b(new_n257), .c(new_n243), .o1(new_n294));
  nano22aa1n02x4               g199(.a(new_n294), .b(new_n260), .c(new_n261), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n276), .o1(new_n296));
  inv000aa1n02x5               g201(.a(new_n284), .o1(new_n297));
  aoai13aa1n12x5               g202(.a(new_n297), .b(new_n296), .c(new_n293), .d(new_n295), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n286), .b(new_n298), .c(new_n188), .d(new_n277), .o1(new_n299));
  nona22aa1n03x5               g204(.a(new_n299), .b(new_n291), .c(new_n289), .out0(new_n300));
  nanp02aa1n03x5               g205(.a(new_n292), .b(new_n300), .o1(\s[28] ));
  and002aa1n02x5               g206(.a(new_n290), .b(new_n286), .o(new_n302));
  aoai13aa1n06x5               g207(.a(new_n302), .b(new_n298), .c(new_n188), .d(new_n277), .o1(new_n303));
  orn002aa1n03x5               g208(.a(\a[27] ), .b(\b[26] ), .o(new_n304));
  oao003aa1n03x5               g209(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n305));
  nanp02aa1n03x5               g210(.a(new_n303), .b(new_n305), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n306), .b(new_n307), .c(new_n303), .d(new_n308), .o1(\s[29] ));
  nanp02aa1n02x5               g214(.a(\b[0] ), .b(\a[1] ), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n310), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g216(.a(new_n290), .b(new_n286), .c(new_n307), .o1(new_n312));
  nanb02aa1n03x5               g217(.a(new_n312), .b(new_n288), .out0(new_n313));
  oaoi03aa1n09x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n305), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n312), .c(new_n278), .d(new_n285), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .out0(new_n317));
  aoi012aa1n02x5               g222(.a(new_n305), .b(\a[29] ), .c(\b[28] ), .o1(new_n318));
  oabi12aa1n02x5               g223(.a(new_n317), .b(\a[29] ), .c(\b[28] ), .out0(new_n319));
  norp02aa1n02x5               g224(.a(new_n318), .b(new_n319), .o1(new_n320));
  aoi022aa1n03x5               g225(.a(new_n320), .b(new_n313), .c(new_n316), .d(new_n317), .o1(\s[30] ));
  norb02aa1n02x5               g226(.a(new_n317), .b(new_n312), .out0(new_n322));
  aoai13aa1n06x5               g227(.a(new_n322), .b(new_n298), .c(new_n188), .d(new_n277), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n315), .carry(new_n324));
  xnrc02aa1n02x5               g229(.a(\b[30] ), .b(\a[31] ), .out0(new_n325));
  aoi012aa1n02x7               g230(.a(new_n325), .b(new_n323), .c(new_n324), .o1(new_n326));
  aobi12aa1n02x7               g231(.a(new_n322), .b(new_n278), .c(new_n285), .out0(new_n327));
  nano22aa1n02x4               g232(.a(new_n327), .b(new_n324), .c(new_n325), .out0(new_n328));
  nor002aa1n02x5               g233(.a(new_n326), .b(new_n328), .o1(\s[31] ));
  xnbna2aa1n03x5               g234(.a(new_n100), .b(new_n102), .c(new_n101), .out0(\s[3] ));
  xnrc02aa1n02x5               g235(.a(\b[3] ), .b(\a[4] ), .out0(new_n331));
  aoi013aa1n02x4               g236(.a(new_n98), .b(new_n102), .c(new_n101), .d(new_n99), .o1(new_n332));
  oaib12aa1n02x5               g237(.a(new_n107), .b(new_n332), .c(new_n331), .out0(\s[4] ));
  and002aa1n02x5               g238(.a(new_n113), .b(new_n119), .o(new_n334));
  nanb02aa1n02x5               g239(.a(new_n104), .b(new_n107), .out0(new_n335));
  xnrc02aa1n02x5               g240(.a(\b[4] ), .b(\a[5] ), .out0(new_n336));
  aoi022aa1n02x5               g241(.a(new_n335), .b(new_n336), .c(new_n334), .d(new_n107), .o1(\s[5] ));
  norb02aa1n02x5               g242(.a(new_n108), .b(new_n118), .out0(new_n338));
  nanp02aa1n02x5               g243(.a(new_n107), .b(new_n334), .o1(new_n339));
  xnbna2aa1n03x5               g244(.a(new_n338), .b(new_n339), .c(new_n119), .out0(\s[6] ));
  norb02aa1n02x5               g245(.a(new_n110), .b(new_n109), .out0(new_n341));
  aoai13aa1n02x5               g246(.a(new_n116), .b(new_n120), .c(new_n107), .d(new_n334), .o1(new_n342));
  aboi22aa1n03x5               g247(.a(new_n120), .b(new_n339), .c(\a[6] ), .d(\b[5] ), .out0(new_n343));
  oa0012aa1n02x5               g248(.a(new_n342), .b(new_n343), .c(new_n341), .o(\s[7] ));
  xnbna2aa1n03x5               g249(.a(new_n117), .b(new_n342), .c(new_n122), .out0(\s[8] ));
  xnbna2aa1n03x5               g250(.a(new_n125), .b(new_n145), .c(new_n146), .out0(\s[9] ));
endmodule


