// Benchmark "adder" written by ABC on Thu Jul 18 15:21:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n312, new_n315, new_n316, new_n318, new_n319, new_n320,
    new_n321, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  tech160nm_fioai012aa1n03p5x5 g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  nor022aa1n04x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n06x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  aoi012aa1n02x5               g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  oai012aa1n06x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  norp02aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n03x5               g016(.a(new_n108), .b(new_n111), .c(new_n110), .d(new_n109), .out0(new_n112));
  tech160nm_fixorc02aa1n02p5x5 g017(.a(\a[6] ), .b(\b[5] ), .out0(new_n113));
  xorc02aa1n02x5               g018(.a(\a[5] ), .b(\b[4] ), .out0(new_n114));
  nano22aa1n03x7               g019(.a(new_n112), .b(new_n113), .c(new_n114), .out0(new_n115));
  and002aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o(new_n116));
  oai022aa1n02x5               g021(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  nanb02aa1n02x5               g022(.a(new_n116), .b(new_n117), .out0(new_n118));
  inv000aa1d42x5               g023(.a(new_n110), .o1(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .o1(new_n120));
  oabi12aa1n06x5               g025(.a(new_n120), .b(new_n112), .c(new_n118), .out0(new_n121));
  aoi012aa1n03x5               g026(.a(new_n121), .b(new_n115), .c(new_n107), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[9] ), .b(\b[8] ), .c(new_n122), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n16x5               g029(.a(\b[10] ), .b(\a[11] ), .o1(new_n125));
  nand42aa1n04x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  nor042aa1n06x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  nor022aa1n08x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand22aa1n04x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  nano23aa1n06x5               g036(.a(new_n128), .b(new_n130), .c(new_n131), .d(new_n129), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n121), .c(new_n115), .d(new_n107), .o1(new_n133));
  aoi012aa1n06x5               g038(.a(new_n130), .b(new_n128), .c(new_n131), .o1(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n127), .b(new_n133), .c(new_n134), .out0(\s[11] ));
  inv040aa1n06x5               g040(.a(new_n125), .o1(new_n136));
  inv000aa1n03x5               g041(.a(new_n122), .o1(new_n137));
  inv040aa1n03x5               g042(.a(new_n134), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n127), .b(new_n138), .c(new_n137), .d(new_n132), .o1(new_n139));
  nor022aa1n16x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanp02aa1n04x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n139), .c(new_n136), .out0(\s[12] ));
  nona23aa1n09x5               g048(.a(new_n141), .b(new_n126), .c(new_n125), .d(new_n140), .out0(new_n144));
  norb02aa1n02x5               g049(.a(new_n132), .b(new_n144), .out0(new_n145));
  aoai13aa1n03x5               g050(.a(new_n145), .b(new_n121), .c(new_n115), .d(new_n107), .o1(new_n146));
  oaoi03aa1n12x5               g051(.a(\a[12] ), .b(\b[11] ), .c(new_n136), .o1(new_n147));
  oabi12aa1n18x5               g052(.a(new_n147), .b(new_n144), .c(new_n134), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n146), .b(new_n149), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1d28x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n152), .b(new_n150), .c(new_n153), .o1(new_n154));
  xnrb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n04x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nand42aa1n20x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nano23aa1d15x5               g062(.a(new_n152), .b(new_n156), .c(new_n157), .d(new_n153), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoi012aa1n09x5               g064(.a(new_n156), .b(new_n152), .c(new_n157), .o1(new_n160));
  aoai13aa1n03x5               g065(.a(new_n160), .b(new_n159), .c(new_n146), .d(new_n149), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  and002aa1n02x5               g068(.a(\b[14] ), .b(\a[15] ), .o(new_n164));
  nona22aa1n03x5               g069(.a(new_n161), .b(new_n164), .c(new_n163), .out0(new_n165));
  nor042aa1n03x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand42aa1n16x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  oai112aa1n02x5               g073(.a(new_n165), .b(new_n168), .c(\b[14] ), .d(\a[15] ), .o1(new_n169));
  oaoi13aa1n02x5               g074(.a(new_n168), .b(new_n165), .c(\a[15] ), .d(\b[14] ), .o1(new_n170));
  norb02aa1n03x4               g075(.a(new_n169), .b(new_n170), .out0(\s[16] ));
  nano23aa1n03x7               g076(.a(new_n125), .b(new_n140), .c(new_n141), .d(new_n126), .out0(new_n172));
  nand42aa1d28x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nano23aa1n03x7               g078(.a(new_n163), .b(new_n166), .c(new_n167), .d(new_n173), .out0(new_n174));
  inv000aa1n02x5               g079(.a(new_n174), .o1(new_n175));
  nano32aa1n03x7               g080(.a(new_n175), .b(new_n158), .c(new_n172), .d(new_n132), .out0(new_n176));
  aoai13aa1n06x5               g081(.a(new_n176), .b(new_n121), .c(new_n107), .d(new_n115), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n160), .o1(new_n178));
  aoai13aa1n04x5               g083(.a(new_n174), .b(new_n178), .c(new_n148), .d(new_n158), .o1(new_n179));
  oai012aa1n02x5               g084(.a(new_n167), .b(new_n166), .c(new_n163), .o1(new_n180));
  nand23aa1n06x5               g085(.a(new_n177), .b(new_n179), .c(new_n180), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1n12x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  nand42aa1n16x5               g088(.a(\b[16] ), .b(\a[17] ), .o1(new_n184));
  tech160nm_fiaoi012aa1n05x5   g089(.a(new_n183), .b(new_n181), .c(new_n184), .o1(new_n185));
  xnrb03aa1n03x5               g090(.a(new_n185), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  aoai13aa1n03x5               g091(.a(new_n158), .b(new_n147), .c(new_n172), .d(new_n138), .o1(new_n187));
  nand02aa1n02x5               g092(.a(new_n187), .b(new_n160), .o1(new_n188));
  aobi12aa1n06x5               g093(.a(new_n180), .b(new_n188), .c(new_n174), .out0(new_n189));
  nor042aa1n06x5               g094(.a(\b[17] ), .b(\a[18] ), .o1(new_n190));
  nand02aa1n12x5               g095(.a(\b[17] ), .b(\a[18] ), .o1(new_n191));
  nano23aa1d15x5               g096(.a(new_n183), .b(new_n190), .c(new_n191), .d(new_n184), .out0(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  aoi012aa1n12x5               g098(.a(new_n190), .b(new_n183), .c(new_n191), .o1(new_n194));
  aoai13aa1n02x7               g099(.a(new_n194), .b(new_n193), .c(new_n189), .d(new_n177), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g101(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand22aa1n06x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  nor022aa1n06x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand22aa1n04x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n02x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  aoi112aa1n02x5               g108(.a(new_n198), .b(new_n203), .c(new_n195), .d(new_n200), .o1(new_n204));
  inv000aa1n06x5               g109(.a(new_n198), .o1(new_n205));
  inv020aa1n03x5               g110(.a(new_n194), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n200), .b(new_n206), .c(new_n181), .d(new_n192), .o1(new_n207));
  aobi12aa1n02x7               g112(.a(new_n203), .b(new_n207), .c(new_n205), .out0(new_n208));
  nor002aa1n02x5               g113(.a(new_n208), .b(new_n204), .o1(\s[20] ));
  nano23aa1n06x5               g114(.a(new_n198), .b(new_n201), .c(new_n202), .d(new_n199), .out0(new_n210));
  nand22aa1n06x5               g115(.a(new_n210), .b(new_n192), .o1(new_n211));
  nona23aa1d18x5               g116(.a(new_n202), .b(new_n199), .c(new_n198), .d(new_n201), .out0(new_n212));
  oaoi03aa1n12x5               g117(.a(\a[20] ), .b(\b[19] ), .c(new_n205), .o1(new_n213));
  inv040aa1n06x5               g118(.a(new_n213), .o1(new_n214));
  oai012aa1d24x5               g119(.a(new_n214), .b(new_n212), .c(new_n194), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n02x7               g121(.a(new_n216), .b(new_n211), .c(new_n189), .d(new_n177), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[21] ), .b(\b[20] ), .out0(new_n220));
  xorc02aa1n02x5               g125(.a(\a[22] ), .b(\b[21] ), .out0(new_n221));
  aoi112aa1n02x5               g126(.a(new_n219), .b(new_n221), .c(new_n217), .d(new_n220), .o1(new_n222));
  inv040aa1n03x5               g127(.a(new_n219), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n211), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n220), .b(new_n215), .c(new_n181), .d(new_n224), .o1(new_n225));
  aobi12aa1n02x7               g130(.a(new_n221), .b(new_n225), .c(new_n223), .out0(new_n226));
  nor002aa1n02x5               g131(.a(new_n226), .b(new_n222), .o1(\s[22] ));
  nano22aa1n03x7               g132(.a(new_n211), .b(new_n220), .c(new_n221), .out0(new_n228));
  inv000aa1n02x5               g133(.a(new_n228), .o1(new_n229));
  inv030aa1d32x5               g134(.a(\a[21] ), .o1(new_n230));
  inv000aa1n06x5               g135(.a(\a[22] ), .o1(new_n231));
  xroi22aa1d06x4               g136(.a(new_n230), .b(\b[20] ), .c(new_n231), .d(\b[21] ), .out0(new_n232));
  oaoi03aa1n09x5               g137(.a(\a[22] ), .b(\b[21] ), .c(new_n223), .o1(new_n233));
  aoi012aa1d18x5               g138(.a(new_n233), .b(new_n215), .c(new_n232), .o1(new_n234));
  aoai13aa1n04x5               g139(.a(new_n234), .b(new_n229), .c(new_n189), .d(new_n177), .o1(new_n235));
  xorb03aa1n02x5               g140(.a(new_n235), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g141(.a(\b[22] ), .b(\a[23] ), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  tech160nm_fixorc02aa1n05x5   g143(.a(\a[24] ), .b(\b[23] ), .out0(new_n239));
  aoi112aa1n02x5               g144(.a(new_n237), .b(new_n239), .c(new_n235), .d(new_n238), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n237), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n234), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n238), .b(new_n242), .c(new_n181), .d(new_n228), .o1(new_n243));
  aobi12aa1n03x5               g148(.a(new_n239), .b(new_n243), .c(new_n241), .out0(new_n244));
  nor002aa1n02x5               g149(.a(new_n244), .b(new_n240), .o1(\s[24] ));
  and002aa1n02x5               g150(.a(new_n239), .b(new_n238), .o(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  nano32aa1n02x4               g152(.a(new_n247), .b(new_n232), .c(new_n210), .d(new_n192), .out0(new_n248));
  inv000aa1n02x5               g153(.a(new_n248), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n232), .b(new_n213), .c(new_n210), .d(new_n206), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n233), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  oai022aa1n02x5               g157(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(new_n253), .b(new_n252), .o1(new_n254));
  aoai13aa1n12x5               g159(.a(new_n254), .b(new_n247), .c(new_n250), .d(new_n251), .o1(new_n255));
  inv000aa1n02x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n02x7               g161(.a(new_n256), .b(new_n249), .c(new_n189), .d(new_n177), .o1(new_n257));
  xorb03aa1n02x5               g162(.a(new_n257), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  tech160nm_fixorc02aa1n02p5x5 g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  xorc02aa1n02x5               g165(.a(\a[26] ), .b(\b[25] ), .out0(new_n261));
  aoi112aa1n02x5               g166(.a(new_n259), .b(new_n261), .c(new_n257), .d(new_n260), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n259), .o1(new_n263));
  aoai13aa1n03x5               g168(.a(new_n260), .b(new_n255), .c(new_n181), .d(new_n248), .o1(new_n264));
  aobi12aa1n02x7               g169(.a(new_n261), .b(new_n264), .c(new_n263), .out0(new_n265));
  nor002aa1n02x5               g170(.a(new_n265), .b(new_n262), .o1(\s[26] ));
  aoai13aa1n02x5               g171(.a(new_n180), .b(new_n175), .c(new_n187), .d(new_n160), .o1(new_n267));
  and002aa1n06x5               g172(.a(new_n261), .b(new_n260), .o(new_n268));
  inv000aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  nano23aa1n06x5               g174(.a(new_n211), .b(new_n269), .c(new_n246), .d(new_n232), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n267), .c(new_n137), .d(new_n176), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n272));
  aobi12aa1n12x5               g177(.a(new_n272), .b(new_n255), .c(new_n268), .out0(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n271), .c(new_n273), .out0(\s[27] ));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  inv040aa1n03x5               g181(.a(new_n276), .o1(new_n277));
  aobi12aa1n02x7               g182(.a(new_n274), .b(new_n271), .c(new_n273), .out0(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[27] ), .b(\a[28] ), .out0(new_n279));
  nano22aa1n03x5               g184(.a(new_n278), .b(new_n277), .c(new_n279), .out0(new_n280));
  aoai13aa1n02x7               g185(.a(new_n246), .b(new_n233), .c(new_n215), .d(new_n232), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n272), .b(new_n269), .c(new_n281), .d(new_n254), .o1(new_n282));
  aoai13aa1n03x5               g187(.a(new_n274), .b(new_n282), .c(new_n181), .d(new_n270), .o1(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n279), .b(new_n283), .c(new_n277), .o1(new_n284));
  nor002aa1n02x5               g189(.a(new_n284), .b(new_n280), .o1(\s[28] ));
  norb02aa1n02x5               g190(.a(new_n274), .b(new_n279), .out0(new_n286));
  aobi12aa1n02x7               g191(.a(new_n286), .b(new_n271), .c(new_n273), .out0(new_n287));
  oao003aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .c(new_n277), .carry(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[28] ), .b(\a[29] ), .out0(new_n289));
  nano22aa1n03x5               g194(.a(new_n287), .b(new_n288), .c(new_n289), .out0(new_n290));
  aoai13aa1n03x5               g195(.a(new_n286), .b(new_n282), .c(new_n181), .d(new_n270), .o1(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n289), .b(new_n291), .c(new_n288), .o1(new_n292));
  norp02aa1n03x5               g197(.a(new_n292), .b(new_n290), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g199(.a(new_n274), .b(new_n289), .c(new_n279), .out0(new_n295));
  aobi12aa1n02x7               g200(.a(new_n295), .b(new_n271), .c(new_n273), .out0(new_n296));
  oao003aa1n02x5               g201(.a(\a[29] ), .b(\b[28] ), .c(new_n288), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[29] ), .b(\a[30] ), .out0(new_n298));
  nano22aa1n02x4               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  aoai13aa1n03x5               g204(.a(new_n295), .b(new_n282), .c(new_n181), .d(new_n270), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  norp02aa1n03x5               g206(.a(new_n301), .b(new_n299), .o1(\s[30] ));
  norb02aa1n02x5               g207(.a(new_n295), .b(new_n298), .out0(new_n303));
  aobi12aa1n02x7               g208(.a(new_n303), .b(new_n271), .c(new_n273), .out0(new_n304));
  oao003aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .c(new_n297), .carry(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  nano22aa1n02x4               g211(.a(new_n304), .b(new_n305), .c(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n303), .b(new_n282), .c(new_n181), .d(new_n270), .o1(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n306), .b(new_n308), .c(new_n305), .o1(new_n309));
  norp02aa1n03x5               g214(.a(new_n309), .b(new_n307), .o1(\s[31] ));
  xnrb03aa1n02x5               g215(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g216(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g218(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai112aa1n02x5               g219(.a(new_n106), .b(new_n114), .c(new_n105), .d(new_n100), .o1(new_n315));
  aob012aa1n02x5               g220(.a(new_n315), .b(\b[4] ), .c(\a[5] ), .out0(new_n316));
  xnrc02aa1n02x5               g221(.a(new_n316), .b(new_n113), .out0(\s[6] ));
  nanb02aa1n02x5               g222(.a(new_n110), .b(new_n111), .out0(new_n318));
  nanp02aa1n02x5               g223(.a(new_n316), .b(new_n113), .o1(new_n319));
  nona22aa1n02x4               g224(.a(new_n319), .b(new_n116), .c(new_n318), .out0(new_n320));
  aoai13aa1n02x5               g225(.a(new_n318), .b(new_n116), .c(new_n316), .d(new_n113), .o1(new_n321));
  and002aa1n02x5               g226(.a(new_n320), .b(new_n321), .o(\s[7] ));
  norb02aa1n02x5               g227(.a(new_n108), .b(new_n109), .out0(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n323), .b(new_n320), .c(new_n119), .out0(\s[8] ));
  xnrb03aa1n02x5               g229(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


