// Benchmark "adder" written by ABC on Wed Jul 17 21:28:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n343, new_n346, new_n348,
    new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n09x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  inv040aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(new_n101), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1d04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n20x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanp02aa1n02x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n03x5               g011(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n107));
  inv000aa1d42x5               g012(.a(\a[2] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[1] ), .o1(new_n109));
  nand22aa1n04x5               g014(.a(\b[0] ), .b(\a[1] ), .o1(new_n110));
  tech160nm_fioaoi03aa1n03p5x5 g015(.a(new_n108), .b(new_n109), .c(new_n110), .o1(new_n111));
  tech160nm_fiaoi012aa1n03p5x5 g016(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n112));
  oai012aa1n04x7               g017(.a(new_n112), .b(new_n107), .c(new_n111), .o1(new_n113));
  nor022aa1n06x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nand42aa1n03x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nona23aa1n03x5               g022(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n118));
  tech160nm_fixnrc02aa1n05x5   g023(.a(\b[5] ), .b(\a[6] ), .out0(new_n119));
  nor042aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nanb02aa1n02x5               g026(.a(new_n120), .b(new_n121), .out0(new_n122));
  nor043aa1n02x5               g027(.a(new_n118), .b(new_n119), .c(new_n122), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\a[6] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[5] ), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(new_n124), .b(new_n125), .c(new_n120), .o1(new_n126));
  oai012aa1n02x5               g031(.a(new_n115), .b(new_n116), .c(new_n114), .o1(new_n127));
  tech160nm_fioai012aa1n04x5   g032(.a(new_n127), .b(new_n118), .c(new_n126), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  nanb02aa1n03x5               g034(.a(new_n101), .b(new_n129), .out0(new_n130));
  inv040aa1n02x5               g035(.a(new_n130), .o1(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n128), .c(new_n113), .d(new_n123), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n100), .b(new_n132), .c(new_n102), .out0(\s[10] ));
  nano23aa1n02x4               g038(.a(new_n103), .b(new_n105), .c(new_n106), .d(new_n104), .out0(new_n134));
  oao003aa1n02x5               g039(.a(new_n108), .b(new_n109), .c(new_n110), .carry(new_n135));
  aobi12aa1n02x5               g040(.a(new_n112), .b(new_n134), .c(new_n135), .out0(new_n136));
  nano23aa1n02x4               g041(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n137));
  nona22aa1n02x4               g042(.a(new_n137), .b(new_n119), .c(new_n122), .out0(new_n138));
  oabi12aa1n06x5               g043(.a(new_n128), .b(new_n136), .c(new_n138), .out0(new_n139));
  aoi012aa1d24x5               g044(.a(new_n97), .b(new_n101), .c(new_n98), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  aoi013aa1n02x4               g046(.a(new_n141), .b(new_n139), .c(new_n131), .d(new_n100), .o1(new_n142));
  nor002aa1d32x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  inv040aa1n08x5               g048(.a(new_n143), .o1(new_n144));
  nand02aa1d28x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n142), .b(new_n145), .c(new_n144), .out0(\s[11] ));
  oaoi03aa1n02x5               g051(.a(\a[11] ), .b(\b[10] ), .c(new_n142), .o1(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1n20x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nand02aa1d28x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nona23aa1n12x5               g055(.a(new_n150), .b(new_n145), .c(new_n143), .d(new_n149), .out0(new_n151));
  oaoi03aa1n12x5               g056(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n152));
  inv020aa1n08x5               g057(.a(new_n152), .o1(new_n153));
  oai012aa1n12x5               g058(.a(new_n153), .b(new_n151), .c(new_n140), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  oai013aa1n02x4               g060(.a(new_n155), .b(new_n132), .c(new_n99), .d(new_n151), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nano23aa1n03x7               g062(.a(new_n143), .b(new_n149), .c(new_n150), .d(new_n145), .out0(new_n158));
  nano22aa1n03x7               g063(.a(new_n132), .b(new_n100), .c(new_n158), .out0(new_n159));
  nor042aa1n12x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nanp02aa1n12x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nanb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  tech160nm_fioai012aa1n05x5   g068(.a(new_n163), .b(new_n159), .c(new_n154), .o1(new_n164));
  nor002aa1d32x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand02aa1d16x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nanb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(new_n167));
  oai112aa1n02x5               g072(.a(new_n164), .b(new_n167), .c(\b[12] ), .d(\a[13] ), .o1(new_n168));
  oaoi13aa1n06x5               g073(.a(new_n167), .b(new_n164), .c(\a[13] ), .d(\b[12] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(\s[14] ));
  aoi112aa1n09x5               g075(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n171));
  norb02aa1n06x4               g076(.a(new_n145), .b(new_n143), .out0(new_n172));
  norb02aa1n12x5               g077(.a(new_n150), .b(new_n149), .out0(new_n173));
  oai112aa1n06x5               g078(.a(new_n172), .b(new_n173), .c(new_n171), .d(new_n97), .o1(new_n174));
  nano23aa1n09x5               g079(.a(new_n160), .b(new_n165), .c(new_n166), .d(new_n161), .out0(new_n175));
  inv020aa1n04x5               g080(.a(new_n175), .o1(new_n176));
  aoi012aa1d24x5               g081(.a(new_n165), .b(new_n160), .c(new_n166), .o1(new_n177));
  aoai13aa1n12x5               g082(.a(new_n177), .b(new_n176), .c(new_n174), .d(new_n153), .o1(new_n178));
  inv000aa1d42x5               g083(.a(new_n178), .o1(new_n179));
  nanp02aa1n03x5               g084(.a(new_n175), .b(new_n158), .o1(new_n180));
  nona23aa1n02x4               g085(.a(new_n139), .b(new_n131), .c(new_n180), .d(new_n99), .out0(new_n181));
  nor042aa1d18x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nand42aa1d28x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n181), .c(new_n179), .out0(\s[15] ));
  inv000aa1d42x5               g090(.a(new_n182), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n184), .o1(new_n187));
  aoai13aa1n02x5               g092(.a(new_n186), .b(new_n187), .c(new_n181), .d(new_n179), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nor042aa1n04x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nand42aa1n16x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nano23aa1d15x5               g096(.a(new_n182), .b(new_n190), .c(new_n191), .d(new_n183), .out0(new_n192));
  oai012aa1n02x5               g097(.a(new_n191), .b(new_n190), .c(new_n182), .o1(new_n193));
  aobi12aa1n12x5               g098(.a(new_n193), .b(new_n178), .c(new_n192), .out0(new_n194));
  nano32aa1n03x7               g099(.a(new_n180), .b(new_n192), .c(new_n100), .d(new_n131), .out0(new_n195));
  aoai13aa1n12x5               g100(.a(new_n195), .b(new_n128), .c(new_n113), .d(new_n123), .o1(new_n196));
  nor042aa1n03x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nanp02aa1n02x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  nanb02aa1n06x5               g103(.a(new_n197), .b(new_n198), .out0(new_n199));
  xobna2aa1n03x5               g104(.a(new_n199), .b(new_n194), .c(new_n196), .out0(\s[17] ));
  xorc02aa1n12x5               g105(.a(\a[18] ), .b(\b[17] ), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  oai112aa1n02x5               g107(.a(new_n194), .b(new_n196), .c(\b[16] ), .d(\a[17] ), .o1(new_n203));
  xnbna2aa1n03x5               g108(.a(new_n202), .b(new_n203), .c(new_n198), .out0(\s[18] ));
  norb02aa1n02x5               g109(.a(new_n201), .b(new_n199), .out0(new_n205));
  inv000aa1n02x5               g110(.a(new_n205), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\a[18] ), .o1(new_n207));
  inv000aa1d42x5               g112(.a(\b[17] ), .o1(new_n208));
  tech160nm_fioaoi03aa1n04x5   g113(.a(new_n207), .b(new_n208), .c(new_n197), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n206), .c(new_n194), .d(new_n196), .o1(new_n210));
  xorb03aa1n02x5               g115(.a(new_n210), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g116(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n03x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  xorc02aa1n02x5               g118(.a(\a[19] ), .b(\b[18] ), .out0(new_n214));
  xorc02aa1n06x5               g119(.a(\a[20] ), .b(\b[19] ), .out0(new_n215));
  aoi112aa1n02x5               g120(.a(new_n213), .b(new_n215), .c(new_n210), .d(new_n214), .o1(new_n216));
  inv040aa1n03x5               g121(.a(new_n213), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n177), .o1(new_n218));
  aoai13aa1n04x5               g123(.a(new_n192), .b(new_n218), .c(new_n154), .d(new_n175), .o1(new_n219));
  nand43aa1n08x5               g124(.a(new_n196), .b(new_n219), .c(new_n193), .o1(new_n220));
  oao003aa1n02x5               g125(.a(new_n207), .b(new_n208), .c(new_n197), .carry(new_n221));
  aoai13aa1n03x5               g126(.a(new_n214), .b(new_n221), .c(new_n220), .d(new_n205), .o1(new_n222));
  xnrc02aa1n12x5               g127(.a(\b[19] ), .b(\a[20] ), .out0(new_n223));
  tech160nm_fiaoi012aa1n03p5x5 g128(.a(new_n223), .b(new_n222), .c(new_n217), .o1(new_n224));
  nor002aa1n02x5               g129(.a(new_n224), .b(new_n216), .o1(\s[20] ));
  tech160nm_fixnrc02aa1n04x5   g130(.a(\b[18] ), .b(\a[19] ), .out0(new_n226));
  nona23aa1d18x5               g131(.a(new_n201), .b(new_n215), .c(new_n226), .d(new_n199), .out0(new_n227));
  oaoi03aa1n09x5               g132(.a(\a[20] ), .b(\b[19] ), .c(new_n217), .o1(new_n228));
  aoi013aa1n02x4               g133(.a(new_n228), .b(new_n221), .c(new_n214), .d(new_n215), .o1(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n227), .c(new_n194), .d(new_n196), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n06x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  nanp02aa1n02x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n233), .b(new_n232), .out0(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[21] ), .b(\a[22] ), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(new_n232), .b(new_n236), .c(new_n230), .d(new_n234), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n232), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n227), .o1(new_n239));
  inv000aa1n02x5               g144(.a(new_n228), .o1(new_n240));
  oai013aa1n06x5               g145(.a(new_n240), .b(new_n209), .c(new_n226), .d(new_n223), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n234), .b(new_n241), .c(new_n220), .d(new_n239), .o1(new_n242));
  tech160nm_fiaoi012aa1n03p5x5 g147(.a(new_n235), .b(new_n242), .c(new_n238), .o1(new_n243));
  nor002aa1n02x5               g148(.a(new_n243), .b(new_n237), .o1(\s[22] ));
  nano22aa1d15x5               g149(.a(new_n235), .b(new_n238), .c(new_n233), .out0(new_n245));
  oaoi03aa1n12x5               g150(.a(\a[22] ), .b(\b[21] ), .c(new_n238), .o1(new_n246));
  aoi012aa1d24x5               g151(.a(new_n246), .b(new_n241), .c(new_n245), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n245), .o1(new_n248));
  norp02aa1n02x5               g153(.a(new_n227), .b(new_n248), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  aoai13aa1n04x5               g155(.a(new_n247), .b(new_n250), .c(new_n194), .d(new_n196), .o1(new_n251));
  xorb03aa1n02x5               g156(.a(new_n251), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n09x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  nanp02aa1n02x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  xorc02aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  aoi112aa1n02x5               g161(.a(new_n253), .b(new_n256), .c(new_n251), .d(new_n255), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n253), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n247), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n255), .b(new_n259), .c(new_n220), .d(new_n249), .o1(new_n260));
  xnrc02aa1n02x5               g165(.a(\b[23] ), .b(\a[24] ), .out0(new_n261));
  tech160nm_fiaoi012aa1n03p5x5 g166(.a(new_n261), .b(new_n260), .c(new_n258), .o1(new_n262));
  nor002aa1n02x5               g167(.a(new_n262), .b(new_n257), .o1(\s[24] ));
  nano22aa1n02x5               g168(.a(new_n261), .b(new_n258), .c(new_n254), .out0(new_n264));
  nano22aa1n02x4               g169(.a(new_n227), .b(new_n245), .c(new_n264), .out0(new_n265));
  inv000aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  nand02aa1d08x5               g171(.a(new_n264), .b(new_n245), .o1(new_n267));
  norp02aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .o1(new_n268));
  aoi112aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n269));
  nanp03aa1n02x5               g174(.a(new_n246), .b(new_n255), .c(new_n256), .o1(new_n270));
  nona22aa1n02x4               g175(.a(new_n270), .b(new_n269), .c(new_n268), .out0(new_n271));
  aoib12aa1n12x5               g176(.a(new_n271), .b(new_n241), .c(new_n267), .out0(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n266), .c(new_n194), .d(new_n196), .o1(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  xorc02aa1n02x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  aoi112aa1n03x4               g182(.a(new_n275), .b(new_n277), .c(new_n273), .d(new_n276), .o1(new_n278));
  inv000aa1n02x5               g183(.a(new_n275), .o1(new_n279));
  inv020aa1n02x5               g184(.a(new_n272), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n276), .b(new_n280), .c(new_n220), .d(new_n265), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n277), .o1(new_n282));
  tech160nm_fiaoi012aa1n03p5x5 g187(.a(new_n282), .b(new_n281), .c(new_n279), .o1(new_n283));
  nor002aa1n02x5               g188(.a(new_n283), .b(new_n278), .o1(\s[26] ));
  and002aa1n02x5               g189(.a(new_n277), .b(new_n276), .o(new_n285));
  inv040aa1n02x5               g190(.a(new_n285), .o1(new_n286));
  nano23aa1n06x5               g191(.a(new_n227), .b(new_n286), .c(new_n245), .d(new_n264), .out0(new_n287));
  inv000aa1n02x5               g192(.a(new_n287), .o1(new_n288));
  nanp03aa1n02x5               g193(.a(new_n221), .b(new_n214), .c(new_n215), .o1(new_n289));
  tech160nm_fiaoi012aa1n04x5   g194(.a(new_n267), .b(new_n289), .c(new_n240), .o1(new_n290));
  oaoi03aa1n12x5               g195(.a(\a[26] ), .b(\b[25] ), .c(new_n279), .o1(new_n291));
  oaoi13aa1n09x5               g196(.a(new_n291), .b(new_n285), .c(new_n290), .d(new_n271), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n288), .c(new_n194), .d(new_n196), .o1(new_n293));
  xorb03aa1n02x5               g198(.a(new_n293), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nanp02aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .out0(new_n296));
  nanb02aa1n06x5               g201(.a(new_n267), .b(new_n241), .out0(new_n297));
  aoi113aa1n02x5               g202(.a(new_n269), .b(new_n268), .c(new_n246), .d(new_n256), .e(new_n255), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n291), .o1(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n286), .c(new_n297), .d(new_n298), .o1(new_n300));
  nor042aa1d18x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  aoi112aa1n03x4               g206(.a(new_n300), .b(new_n301), .c(new_n220), .d(new_n287), .o1(new_n302));
  nano22aa1n03x7               g207(.a(new_n302), .b(new_n295), .c(new_n296), .out0(new_n303));
  aoai13aa1n02x5               g208(.a(new_n175), .b(new_n152), .c(new_n158), .d(new_n141), .o1(new_n304));
  inv000aa1d42x5               g209(.a(new_n192), .o1(new_n305));
  aoai13aa1n02x5               g210(.a(new_n193), .b(new_n305), .c(new_n304), .d(new_n177), .o1(new_n306));
  aoai13aa1n02x5               g211(.a(new_n287), .b(new_n306), .c(new_n139), .d(new_n195), .o1(new_n307));
  oaoi13aa1n02x5               g212(.a(new_n286), .b(new_n298), .c(new_n229), .d(new_n267), .o1(new_n308));
  nona32aa1n02x4               g213(.a(new_n307), .b(new_n301), .c(new_n291), .d(new_n308), .out0(new_n309));
  aoi012aa1n02x5               g214(.a(new_n296), .b(new_n309), .c(new_n295), .o1(new_n310));
  norp02aa1n03x5               g215(.a(new_n310), .b(new_n303), .o1(\s[28] ));
  nano22aa1n02x4               g216(.a(new_n301), .b(new_n296), .c(new_n295), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n300), .c(new_n220), .d(new_n287), .o1(new_n313));
  inv000aa1d42x5               g218(.a(\a[28] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(\b[27] ), .o1(new_n315));
  oaoi03aa1n12x5               g220(.a(new_n314), .b(new_n315), .c(new_n301), .o1(new_n316));
  xorc02aa1n12x5               g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  inv000aa1d42x5               g222(.a(new_n317), .o1(new_n318));
  tech160nm_fiaoi012aa1n02p5x5 g223(.a(new_n318), .b(new_n313), .c(new_n316), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n316), .o1(new_n320));
  aoi112aa1n03x4               g225(.a(new_n317), .b(new_n320), .c(new_n293), .d(new_n312), .o1(new_n321));
  norp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[29] ));
  xorb03aa1n02x5               g227(.a(new_n110), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano23aa1n02x4               g228(.a(new_n318), .b(new_n301), .c(new_n296), .d(new_n295), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n300), .c(new_n220), .d(new_n287), .o1(new_n325));
  tech160nm_fioaoi03aa1n03p5x5 g230(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .o1(new_n326));
  inv040aa1n03x5               g231(.a(new_n326), .o1(new_n327));
  xorc02aa1n12x5               g232(.a(\a[30] ), .b(\b[29] ), .out0(new_n328));
  inv000aa1d42x5               g233(.a(new_n328), .o1(new_n329));
  tech160nm_fiaoi012aa1n03p5x5 g234(.a(new_n329), .b(new_n325), .c(new_n327), .o1(new_n330));
  aoi112aa1n03x4               g235(.a(new_n328), .b(new_n326), .c(new_n293), .d(new_n324), .o1(new_n331));
  nor002aa1n02x5               g236(.a(new_n330), .b(new_n331), .o1(\s[30] ));
  and003aa1n02x5               g237(.a(new_n312), .b(new_n328), .c(new_n317), .o(new_n333));
  tech160nm_fioaoi03aa1n02p5x5 g238(.a(\a[30] ), .b(\b[29] ), .c(new_n327), .o1(new_n334));
  xorc02aa1n02x5               g239(.a(\a[31] ), .b(\b[30] ), .out0(new_n335));
  aoi112aa1n03x4               g240(.a(new_n335), .b(new_n334), .c(new_n293), .d(new_n333), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n333), .b(new_n300), .c(new_n220), .d(new_n287), .o1(new_n337));
  inv000aa1n02x5               g242(.a(new_n334), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n335), .o1(new_n339));
  tech160nm_fiaoi012aa1n03p5x5 g244(.a(new_n339), .b(new_n337), .c(new_n338), .o1(new_n340));
  nor042aa1n03x5               g245(.a(new_n340), .b(new_n336), .o1(\s[31] ));
  xnrb03aa1n02x5               g246(.a(new_n111), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g247(.a(\a[3] ), .b(\b[2] ), .c(new_n111), .o1(new_n343));
  xorb03aa1n02x5               g248(.a(new_n343), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g249(.a(new_n113), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n02x5               g250(.a(new_n121), .b(new_n113), .c(new_n120), .o1(new_n346));
  xorb03aa1n02x5               g251(.a(new_n346), .b(\b[5] ), .c(new_n124), .out0(\s[6] ));
  oaoi03aa1n02x5               g252(.a(\a[6] ), .b(\b[5] ), .c(new_n346), .o1(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g254(.a(new_n116), .b(new_n348), .c(new_n117), .o1(new_n350));
  xnrb03aa1n02x5               g255(.a(new_n350), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g256(.a(new_n139), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


