// Benchmark "adder" written by ABC on Wed Jul 17 13:01:14 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n317, new_n319, new_n320,
    new_n321, new_n322, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n12x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor042aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  norp02aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nor002aa1n03x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nano23aa1n03x7               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\a[6] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[5] ), .o1(new_n108));
  nor002aa1n02x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  oao003aa1n02x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .carry(new_n110));
  inv000aa1d42x5               g015(.a(new_n104), .o1(new_n111));
  oaoi03aa1n02x5               g016(.a(\a[8] ), .b(\b[7] ), .c(new_n111), .o1(new_n112));
  tech160nm_fiaoi012aa1n03p5x5 g017(.a(new_n112), .b(new_n106), .c(new_n110), .o1(new_n113));
  norp02aa1n02x5               g018(.a(\b[3] ), .b(\a[4] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[3] ), .b(\a[4] ), .o1(new_n115));
  nor022aa1n04x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  nano23aa1n02x4               g022(.a(new_n114), .b(new_n116), .c(new_n117), .d(new_n115), .out0(new_n118));
  and002aa1n02x5               g023(.a(\b[1] ), .b(\a[2] ), .o(new_n119));
  nanp02aa1n02x5               g024(.a(\b[0] ), .b(\a[1] ), .o1(new_n120));
  nor002aa1n02x5               g025(.a(\b[1] ), .b(\a[2] ), .o1(new_n121));
  oab012aa1n02x4               g026(.a(new_n119), .b(new_n121), .c(new_n120), .out0(new_n122));
  nanp02aa1n02x5               g027(.a(new_n118), .b(new_n122), .o1(new_n123));
  aoi012aa1n02x7               g028(.a(new_n114), .b(new_n116), .c(new_n115), .o1(new_n124));
  xorc02aa1n02x5               g029(.a(\a[6] ), .b(\b[5] ), .out0(new_n125));
  xorc02aa1n02x5               g030(.a(\a[5] ), .b(\b[4] ), .out0(new_n126));
  nanp03aa1n02x5               g031(.a(new_n106), .b(new_n125), .c(new_n126), .o1(new_n127));
  aoai13aa1n06x5               g032(.a(new_n113), .b(new_n127), .c(new_n123), .d(new_n124), .o1(new_n128));
  aob012aa1n03x5               g033(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n99), .b(new_n129), .c(new_n101), .out0(\s[10] ));
  aoi013aa1n03x5               g035(.a(new_n98), .b(new_n129), .c(new_n101), .d(new_n99), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n02x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanp02aa1n02x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n06x4               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  nor002aa1n04x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1n10x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n09x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  aoai13aa1n03x5               g044(.a(new_n139), .b(new_n133), .c(new_n131), .d(new_n135), .o1(new_n140));
  nona32aa1n02x4               g045(.a(new_n129), .b(new_n100), .c(new_n98), .d(new_n97), .out0(new_n141));
  nanb03aa1n02x5               g046(.a(new_n98), .b(new_n141), .c(new_n135), .out0(new_n142));
  nona22aa1n02x4               g047(.a(new_n142), .b(new_n139), .c(new_n133), .out0(new_n143));
  nanp02aa1n02x5               g048(.a(new_n140), .b(new_n143), .o1(\s[12] ));
  aoi112aa1n02x5               g049(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n145));
  oai112aa1n03x5               g050(.a(new_n138), .b(new_n135), .c(new_n145), .d(new_n97), .o1(new_n146));
  aoi012aa1n02x5               g051(.a(new_n136), .b(new_n133), .c(new_n137), .o1(new_n147));
  and002aa1n02x5               g052(.a(new_n146), .b(new_n147), .o(new_n148));
  nona23aa1n06x5               g053(.a(new_n105), .b(new_n103), .c(new_n102), .d(new_n104), .out0(new_n149));
  oaoi03aa1n02x5               g054(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n150));
  oabi12aa1n02x5               g055(.a(new_n112), .b(new_n149), .c(new_n150), .out0(new_n151));
  nona23aa1n03x5               g056(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n152));
  oabi12aa1n02x5               g057(.a(new_n119), .b(new_n120), .c(new_n121), .out0(new_n153));
  tech160nm_fioai012aa1n04x5   g058(.a(new_n124), .b(new_n152), .c(new_n153), .o1(new_n154));
  nano22aa1n02x5               g059(.a(new_n149), .b(new_n125), .c(new_n126), .out0(new_n155));
  xorc02aa1n02x5               g060(.a(\a[9] ), .b(\b[8] ), .out0(new_n156));
  nano32aa1n02x4               g061(.a(new_n139), .b(new_n156), .c(new_n99), .d(new_n135), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n151), .c(new_n155), .d(new_n154), .o1(new_n158));
  tech160nm_fixorc02aa1n02p5x5 g063(.a(\a[13] ), .b(\b[12] ), .out0(new_n159));
  xnbna2aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n148), .out0(\s[13] ));
  inv000aa1d42x5               g065(.a(\a[14] ), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(new_n158), .b(new_n148), .o1(new_n162));
  nor042aa1n03x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n163), .b(new_n162), .c(new_n159), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[13] ), .c(new_n161), .out0(\s[14] ));
  xorc02aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  and002aa1n02x5               g071(.a(new_n166), .b(new_n159), .o(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  inv000aa1d42x5               g073(.a(\b[13] ), .o1(new_n169));
  oao003aa1n09x5               g074(.a(new_n161), .b(new_n169), .c(new_n163), .carry(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  aoai13aa1n06x5               g076(.a(new_n171), .b(new_n168), .c(new_n158), .d(new_n148), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nanp02aa1n04x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nor022aa1n04x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nand42aa1n03x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n174), .c(new_n172), .d(new_n175), .o1(new_n179));
  aoi112aa1n03x5               g084(.a(new_n178), .b(new_n174), .c(new_n172), .d(new_n175), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(\s[16] ));
  nano23aa1n09x5               g086(.a(new_n174), .b(new_n176), .c(new_n177), .d(new_n175), .out0(new_n182));
  tech160nm_fiao0012aa1n02p5x5 g087(.a(new_n176), .b(new_n174), .c(new_n177), .o(new_n183));
  aoi012aa1n06x5               g088(.a(new_n183), .b(new_n182), .c(new_n170), .o1(new_n184));
  nand23aa1n03x5               g089(.a(new_n182), .b(new_n159), .c(new_n166), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n184), .b(new_n185), .c(new_n147), .d(new_n146), .o1(new_n186));
  inv040aa1n03x5               g091(.a(new_n186), .o1(new_n187));
  nano23aa1n02x4               g092(.a(new_n133), .b(new_n136), .c(new_n137), .d(new_n134), .out0(new_n188));
  nano32aa1n03x7               g093(.a(new_n185), .b(new_n156), .c(new_n188), .d(new_n99), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n151), .c(new_n155), .d(new_n154), .o1(new_n190));
  nanp02aa1n06x5               g095(.a(new_n190), .b(new_n187), .o1(new_n191));
  xorb03aa1n02x5               g096(.a(new_n191), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g097(.a(\a[18] ), .o1(new_n193));
  inv040aa1d30x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  oaoi03aa1n02x5               g100(.a(new_n194), .b(new_n195), .c(new_n191), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  xroi22aa1d06x4               g102(.a(new_n194), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  nor002aa1n02x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  aoi112aa1n03x5               g105(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n201));
  norp02aa1n06x5               g106(.a(new_n201), .b(new_n200), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n187), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand02aa1n04x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nor042aa1n06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1d12x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n12x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n206), .c(new_n203), .d(new_n207), .o1(new_n212));
  norb02aa1n03x4               g117(.a(new_n207), .b(new_n206), .out0(new_n213));
  nanp02aa1n02x5               g118(.a(new_n203), .b(new_n213), .o1(new_n214));
  nona22aa1n02x4               g119(.a(new_n214), .b(new_n211), .c(new_n206), .out0(new_n215));
  nanp02aa1n02x5               g120(.a(new_n215), .b(new_n212), .o1(\s[20] ));
  nona23aa1n12x5               g121(.a(new_n209), .b(new_n207), .c(new_n206), .d(new_n208), .out0(new_n217));
  aoi012aa1n06x5               g122(.a(new_n208), .b(new_n206), .c(new_n209), .o1(new_n218));
  oai012aa1n12x5               g123(.a(new_n218), .b(new_n217), .c(new_n202), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  nanb02aa1n06x5               g125(.a(new_n217), .b(new_n198), .out0(new_n221));
  aoai13aa1n06x5               g126(.a(new_n220), .b(new_n221), .c(new_n190), .d(new_n187), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor022aa1n03x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  tech160nm_fixorc02aa1n05x5   g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  tech160nm_fixnrc02aa1n04x5   g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  aoai13aa1n03x5               g131(.a(new_n226), .b(new_n224), .c(new_n222), .d(new_n225), .o1(new_n227));
  nanp02aa1n02x5               g132(.a(new_n222), .b(new_n225), .o1(new_n228));
  nona22aa1n02x4               g133(.a(new_n228), .b(new_n226), .c(new_n224), .out0(new_n229));
  nanp02aa1n02x5               g134(.a(new_n229), .b(new_n227), .o1(\s[22] ));
  oai112aa1n06x5               g135(.a(new_n213), .b(new_n210), .c(new_n201), .d(new_n200), .o1(new_n231));
  nanb02aa1n03x5               g136(.a(new_n226), .b(new_n225), .out0(new_n232));
  inv000aa1d42x5               g137(.a(\a[22] ), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\b[21] ), .o1(new_n234));
  oaoi03aa1n12x5               g139(.a(new_n233), .b(new_n234), .c(new_n224), .o1(new_n235));
  aoai13aa1n12x5               g140(.a(new_n235), .b(new_n232), .c(new_n231), .d(new_n218), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nona23aa1n08x5               g142(.a(new_n198), .b(new_n225), .c(new_n226), .d(new_n217), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n237), .b(new_n238), .c(new_n190), .d(new_n187), .o1(new_n239));
  xorb03aa1n02x5               g144(.a(new_n239), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  xorc02aa1n02x5               g146(.a(\a[23] ), .b(\b[22] ), .out0(new_n242));
  xorc02aa1n12x5               g147(.a(\a[24] ), .b(\b[23] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n241), .c(new_n239), .d(new_n242), .o1(new_n245));
  nanp02aa1n02x5               g150(.a(new_n239), .b(new_n242), .o1(new_n246));
  nona22aa1n02x4               g151(.a(new_n246), .b(new_n244), .c(new_n241), .out0(new_n247));
  nanp02aa1n02x5               g152(.a(new_n247), .b(new_n245), .o1(\s[24] ));
  norb02aa1n02x5               g153(.a(new_n225), .b(new_n226), .out0(new_n249));
  and002aa1n02x5               g154(.a(new_n243), .b(new_n242), .o(new_n250));
  nano22aa1n06x5               g155(.a(new_n221), .b(new_n250), .c(new_n249), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n186), .c(new_n128), .d(new_n189), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n235), .o1(new_n253));
  aoai13aa1n04x5               g158(.a(new_n250), .b(new_n253), .c(new_n219), .d(new_n249), .o1(new_n254));
  inv000aa1d42x5               g159(.a(\a[24] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(\b[23] ), .o1(new_n256));
  oaoi03aa1n12x5               g161(.a(new_n255), .b(new_n256), .c(new_n241), .o1(new_n257));
  nanp02aa1n03x5               g162(.a(new_n254), .b(new_n257), .o1(new_n258));
  nanb02aa1n03x5               g163(.a(new_n258), .b(new_n252), .out0(new_n259));
  xorb03aa1n02x5               g164(.a(new_n259), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xorc02aa1n12x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n261), .c(new_n259), .d(new_n262), .o1(new_n265));
  aoai13aa1n02x5               g170(.a(new_n262), .b(new_n258), .c(new_n191), .d(new_n251), .o1(new_n266));
  nona22aa1n02x4               g171(.a(new_n266), .b(new_n264), .c(new_n261), .out0(new_n267));
  nanp02aa1n03x5               g172(.a(new_n265), .b(new_n267), .o1(\s[26] ));
  inv000aa1d42x5               g173(.a(new_n257), .o1(new_n269));
  and002aa1n06x5               g174(.a(new_n263), .b(new_n262), .o(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n269), .c(new_n236), .d(new_n250), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n272));
  oab012aa1n02x4               g177(.a(new_n272), .b(\a[26] ), .c(\b[25] ), .out0(new_n273));
  nano22aa1n03x7               g178(.a(new_n238), .b(new_n250), .c(new_n270), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n186), .c(new_n128), .d(new_n189), .o1(new_n275));
  nand43aa1n04x5               g180(.a(new_n275), .b(new_n271), .c(new_n273), .o1(new_n276));
  xorb03aa1n02x5               g181(.a(new_n276), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  xorc02aa1n02x5               g183(.a(\a[27] ), .b(\b[26] ), .out0(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[27] ), .b(\a[28] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n278), .c(new_n276), .d(new_n279), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n270), .o1(new_n282));
  aoai13aa1n06x5               g187(.a(new_n273), .b(new_n282), .c(new_n254), .d(new_n257), .o1(new_n283));
  aobi12aa1n12x5               g188(.a(new_n274), .b(new_n190), .c(new_n187), .out0(new_n284));
  oaih12aa1n02x5               g189(.a(new_n279), .b(new_n283), .c(new_n284), .o1(new_n285));
  nona22aa1n02x5               g190(.a(new_n285), .b(new_n280), .c(new_n278), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n281), .b(new_n286), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n279), .b(new_n280), .out0(new_n288));
  oaih12aa1n02x5               g193(.a(new_n288), .b(new_n283), .c(new_n284), .o1(new_n289));
  aob012aa1n02x5               g194(.a(new_n278), .b(\b[27] ), .c(\a[28] ), .out0(new_n290));
  oa0012aa1n12x5               g195(.a(new_n290), .b(\b[27] ), .c(\a[28] ), .o(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  nona22aa1n02x5               g198(.a(new_n289), .b(new_n292), .c(new_n293), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n293), .b(new_n292), .c(new_n276), .d(new_n288), .o1(new_n295));
  nanp02aa1n03x5               g200(.a(new_n295), .b(new_n294), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n120), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g202(.a(new_n279), .b(new_n293), .c(new_n280), .out0(new_n298));
  oaoi03aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .o1(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[29] ), .b(\a[30] ), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n299), .c(new_n276), .d(new_n298), .o1(new_n301));
  oaih12aa1n02x5               g206(.a(new_n298), .b(new_n283), .c(new_n284), .o1(new_n302));
  nona22aa1n02x5               g207(.a(new_n302), .b(new_n299), .c(new_n300), .out0(new_n303));
  nanp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[30] ));
  nanb02aa1n02x5               g209(.a(new_n300), .b(new_n299), .out0(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(\b[29] ), .c(\a[30] ), .o1(new_n306));
  norb02aa1n02x5               g211(.a(new_n298), .b(new_n300), .out0(new_n307));
  oaih12aa1n02x5               g212(.a(new_n307), .b(new_n283), .c(new_n284), .o1(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[30] ), .b(\a[31] ), .out0(new_n309));
  nona22aa1n02x5               g214(.a(new_n308), .b(new_n309), .c(new_n306), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n309), .b(new_n306), .c(new_n276), .d(new_n307), .o1(new_n311));
  nanp02aa1n03x5               g216(.a(new_n311), .b(new_n310), .o1(\s[31] ));
  xorb03aa1n02x5               g217(.a(new_n122), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi012aa1n02x5               g218(.a(new_n116), .b(new_n122), .c(new_n117), .o1(new_n314));
  xnrb03aa1n02x5               g219(.a(new_n314), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g220(.a(new_n154), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g221(.a(new_n109), .b(new_n154), .c(new_n126), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[5] ), .c(new_n107), .out0(\s[6] ));
  and002aa1n02x5               g223(.a(\b[5] ), .b(\a[6] ), .o(new_n319));
  nanp02aa1n02x5               g224(.a(new_n317), .b(new_n125), .o1(new_n320));
  nona23aa1n02x4               g225(.a(new_n320), .b(new_n105), .c(new_n104), .d(new_n319), .out0(new_n321));
  aboi22aa1n03x5               g226(.a(new_n319), .b(new_n320), .c(new_n111), .d(new_n105), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n321), .b(new_n322), .out0(\s[7] ));
  norb02aa1n02x5               g228(.a(new_n103), .b(new_n102), .out0(new_n324));
  xnbna2aa1n03x5               g229(.a(new_n324), .b(new_n321), .c(new_n111), .out0(\s[8] ));
  xorb03aa1n02x5               g230(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


