// Benchmark "adder" written by ABC on Wed Jul 17 18:13:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n340, new_n341, new_n342, new_n344, new_n345, new_n346,
    new_n348, new_n350, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n09x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nor042aa1n09x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nand42aa1n16x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nano23aa1d15x5               g005(.a(new_n97), .b(new_n99), .c(new_n100), .d(new_n98), .out0(new_n101));
  nona23aa1n02x4               g006(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n102));
  nor002aa1n06x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nand22aa1n04x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nor042aa1n04x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  aoi012aa1n06x5               g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  ao0012aa1n03x7               g011(.a(new_n97), .b(new_n99), .c(new_n98), .o(new_n107));
  oabi12aa1n06x5               g012(.a(new_n107), .b(new_n102), .c(new_n106), .out0(new_n108));
  oa0022aa1n06x5               g013(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n109));
  inv040aa1d32x5               g014(.a(\a[3] ), .o1(new_n110));
  inv040aa1d28x5               g015(.a(\b[2] ), .o1(new_n111));
  nanp02aa1n06x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nand22aa1n04x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nand02aa1n08x5               g018(.a(new_n112), .b(new_n113), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nor042aa1n06x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand22aa1n12x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  oaih12aa1n12x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  oai012aa1d24x5               g023(.a(new_n109), .b(new_n118), .c(new_n114), .o1(new_n119));
  nand02aa1n06x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nanp02aa1n12x5               g025(.a(\b[3] ), .b(\a[4] ), .o1(new_n121));
  oai012aa1n12x5               g026(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .o1(new_n122));
  nano23aa1d15x5               g027(.a(new_n122), .b(new_n103), .c(new_n104), .d(new_n120), .out0(new_n123));
  aoi013aa1n09x5               g028(.a(new_n108), .b(new_n119), .c(new_n101), .d(new_n123), .o1(new_n124));
  oaoi03aa1n09x5               g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  nor002aa1d32x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand02aa1d08x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1n15x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  norp02aa1n24x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  aoib12aa1n12x5               g034(.a(new_n107), .b(new_n101), .c(new_n106), .out0(new_n130));
  nand23aa1n06x5               g035(.a(new_n119), .b(new_n101), .c(new_n123), .o1(new_n131));
  nand02aa1d10x5               g036(.a(new_n131), .b(new_n130), .o1(new_n132));
  xnrc02aa1n12x5               g037(.a(\b[8] ), .b(\a[9] ), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  aoi112aa1n02x5               g039(.a(new_n128), .b(new_n129), .c(new_n132), .d(new_n134), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n135), .b(new_n125), .c(new_n128), .o1(\s[10] ));
  aoai13aa1n02x5               g041(.a(new_n128), .b(new_n129), .c(new_n132), .d(new_n134), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n126), .b(new_n129), .c(new_n127), .o1(new_n138));
  nor002aa1d32x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand02aa1d28x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n06x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n137), .c(new_n138), .out0(\s[11] ));
  norp02aa1n09x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n08x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  inv000aa1n02x5               g050(.a(new_n138), .o1(new_n146));
  aoi112aa1n06x5               g051(.a(new_n139), .b(new_n146), .c(new_n125), .d(new_n128), .o1(new_n147));
  nano22aa1n03x7               g052(.a(new_n147), .b(new_n140), .c(new_n145), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n140), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n144), .b(new_n143), .out0(new_n150));
  oai012aa1n03x5               g055(.a(new_n150), .b(new_n147), .c(new_n149), .o1(new_n151));
  nanb02aa1n03x5               g056(.a(new_n148), .b(new_n151), .out0(\s[12] ));
  nona23aa1d18x5               g057(.a(new_n128), .b(new_n141), .c(new_n133), .d(new_n145), .out0(new_n153));
  nanp02aa1n03x5               g058(.a(new_n129), .b(new_n127), .o1(new_n154));
  nona22aa1n03x5               g059(.a(new_n154), .b(new_n139), .c(new_n126), .out0(new_n155));
  aoai13aa1n04x5               g060(.a(new_n144), .b(new_n143), .c(new_n155), .d(new_n140), .o1(new_n156));
  aoai13aa1n06x5               g061(.a(new_n156), .b(new_n153), .c(new_n131), .d(new_n130), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n20x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  aoi012aa1n02x5               g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n02x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n12x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand22aa1n12x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1d15x5               g069(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n165));
  nanp02aa1n03x5               g070(.a(new_n157), .b(new_n165), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n163), .b(new_n159), .c(new_n164), .o1(new_n167));
  orn002aa1n24x5               g072(.a(\a[15] ), .b(\b[14] ), .o(new_n168));
  nand02aa1n16x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand02aa1d28x5               g074(.a(new_n168), .b(new_n169), .o1(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n166), .c(new_n167), .out0(\s[15] ));
  nand22aa1n02x5               g077(.a(new_n166), .b(new_n167), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n168), .o1(new_n174));
  xnrc02aa1n12x5               g079(.a(\b[15] ), .b(\a[16] ), .out0(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n174), .c(new_n173), .d(new_n169), .o1(new_n176));
  nand42aa1n03x5               g081(.a(new_n173), .b(new_n171), .o1(new_n177));
  nona22aa1n02x4               g082(.a(new_n177), .b(new_n175), .c(new_n174), .out0(new_n178));
  nanp02aa1n03x5               g083(.a(new_n178), .b(new_n176), .o1(\s[16] ));
  nona22aa1d24x5               g084(.a(new_n165), .b(new_n175), .c(new_n170), .out0(new_n180));
  nor042aa1n09x5               g085(.a(new_n153), .b(new_n180), .o1(new_n181));
  nand02aa1d06x5               g086(.a(new_n132), .b(new_n181), .o1(new_n182));
  aoi112aa1n03x5               g087(.a(new_n126), .b(new_n139), .c(new_n129), .d(new_n127), .o1(new_n183));
  oai022aa1n06x5               g088(.a(new_n183), .b(new_n149), .c(\b[11] ), .d(\a[12] ), .o1(new_n184));
  nona23aa1n09x5               g089(.a(new_n164), .b(new_n160), .c(new_n159), .d(new_n163), .out0(new_n185));
  nor043aa1n06x5               g090(.a(new_n185), .b(new_n170), .c(new_n175), .o1(new_n186));
  orn002aa1n02x5               g091(.a(\a[16] ), .b(\b[15] ), .o(new_n187));
  and002aa1n02x5               g092(.a(\b[15] ), .b(\a[16] ), .o(new_n188));
  aoai13aa1n06x5               g093(.a(new_n169), .b(new_n163), .c(new_n159), .d(new_n164), .o1(new_n189));
  aoai13aa1n06x5               g094(.a(new_n187), .b(new_n188), .c(new_n189), .d(new_n168), .o1(new_n190));
  aoi013aa1n09x5               g095(.a(new_n190), .b(new_n186), .c(new_n184), .d(new_n144), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[17] ), .b(\b[16] ), .out0(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n192), .b(new_n182), .c(new_n191), .out0(\s[17] ));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[16] ), .o1(new_n195));
  nanp02aa1n02x5               g100(.a(new_n195), .b(new_n194), .o1(new_n196));
  oabi12aa1n18x5               g101(.a(new_n190), .b(new_n156), .c(new_n180), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n192), .b(new_n197), .c(new_n132), .d(new_n181), .o1(new_n198));
  nor002aa1n10x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nand22aa1n12x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nanb02aa1n12x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  xobna2aa1n03x5               g106(.a(new_n201), .b(new_n198), .c(new_n196), .out0(\s[18] ));
  nanp02aa1n02x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  nano22aa1n12x5               g108(.a(new_n201), .b(new_n196), .c(new_n203), .out0(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n197), .c(new_n132), .d(new_n181), .o1(new_n205));
  aoi013aa1n09x5               g110(.a(new_n199), .b(new_n200), .c(new_n194), .d(new_n195), .o1(new_n206));
  nor002aa1d32x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand02aa1d08x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n12x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n205), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g116(.a(new_n205), .b(new_n206), .o1(new_n212));
  nor002aa1d32x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d28x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1n15x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n207), .c(new_n212), .d(new_n208), .o1(new_n217));
  nano32aa1n03x5               g122(.a(new_n133), .b(new_n150), .c(new_n128), .d(new_n141), .out0(new_n218));
  nand22aa1n03x5               g123(.a(new_n218), .b(new_n186), .o1(new_n219));
  oai012aa1n09x5               g124(.a(new_n191), .b(new_n124), .c(new_n219), .o1(new_n220));
  oaoi03aa1n02x5               g125(.a(\a[18] ), .b(\b[17] ), .c(new_n196), .o1(new_n221));
  aoai13aa1n03x5               g126(.a(new_n209), .b(new_n221), .c(new_n220), .d(new_n204), .o1(new_n222));
  nona22aa1n03x5               g127(.a(new_n222), .b(new_n216), .c(new_n207), .out0(new_n223));
  nanp02aa1n03x5               g128(.a(new_n217), .b(new_n223), .o1(\s[20] ));
  nano23aa1n09x5               g129(.a(new_n207), .b(new_n213), .c(new_n214), .d(new_n208), .out0(new_n225));
  nand22aa1n09x5               g130(.a(new_n204), .b(new_n225), .o1(new_n226));
  nona23aa1n09x5               g131(.a(new_n214), .b(new_n208), .c(new_n207), .d(new_n213), .out0(new_n227));
  oaih12aa1n06x5               g132(.a(new_n214), .b(new_n213), .c(new_n207), .o1(new_n228));
  oai012aa1n18x5               g133(.a(new_n228), .b(new_n227), .c(new_n206), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n226), .c(new_n182), .d(new_n191), .o1(new_n231));
  xnrc02aa1n12x5               g136(.a(\b[20] ), .b(\a[21] ), .out0(new_n232));
  inv040aa1n03x5               g137(.a(new_n232), .o1(new_n233));
  inv040aa1n06x5               g138(.a(new_n226), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n233), .b(new_n229), .c(new_n220), .d(new_n234), .o1(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(new_n231), .c(new_n233), .o1(\s[21] ));
  nor042aa1n09x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  tech160nm_fixnrc02aa1n05x5   g142(.a(\b[21] ), .b(\a[22] ), .out0(new_n238));
  aoai13aa1n02x5               g143(.a(new_n238), .b(new_n237), .c(new_n231), .d(new_n233), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n233), .b(new_n229), .c(new_n220), .d(new_n234), .o1(new_n240));
  nona22aa1n02x4               g145(.a(new_n240), .b(new_n238), .c(new_n237), .out0(new_n241));
  nanp02aa1n02x5               g146(.a(new_n239), .b(new_n241), .o1(\s[22] ));
  nanb02aa1n06x5               g147(.a(new_n238), .b(new_n233), .out0(new_n243));
  nano22aa1n02x4               g148(.a(new_n243), .b(new_n204), .c(new_n225), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n197), .c(new_n132), .d(new_n181), .o1(new_n245));
  aoi112aa1n09x5               g150(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n246));
  oai112aa1n06x5               g151(.a(new_n209), .b(new_n215), .c(new_n246), .d(new_n199), .o1(new_n247));
  inv000aa1d42x5               g152(.a(\a[22] ), .o1(new_n248));
  inv040aa1d32x5               g153(.a(\b[21] ), .o1(new_n249));
  oao003aa1n03x5               g154(.a(new_n248), .b(new_n249), .c(new_n237), .carry(new_n250));
  inv040aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  aoai13aa1n12x5               g156(.a(new_n251), .b(new_n243), .c(new_n247), .d(new_n228), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  xorc02aa1n12x5               g158(.a(\a[23] ), .b(\b[22] ), .out0(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n245), .c(new_n253), .out0(\s[23] ));
  nand02aa1n03x5               g160(.a(new_n245), .b(new_n253), .o1(new_n256));
  norp02aa1n02x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  tech160nm_fixnrc02aa1n04x5   g162(.a(\b[23] ), .b(\a[24] ), .out0(new_n258));
  aoai13aa1n02x5               g163(.a(new_n258), .b(new_n257), .c(new_n256), .d(new_n254), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n254), .b(new_n252), .c(new_n220), .d(new_n244), .o1(new_n260));
  nona22aa1n03x5               g165(.a(new_n260), .b(new_n258), .c(new_n257), .out0(new_n261));
  nanp02aa1n03x5               g166(.a(new_n259), .b(new_n261), .o1(\s[24] ));
  nor042aa1n02x5               g167(.a(new_n238), .b(new_n232), .o1(new_n263));
  norb02aa1n03x5               g168(.a(new_n254), .b(new_n258), .out0(new_n264));
  nanb03aa1n02x5               g169(.a(new_n226), .b(new_n264), .c(new_n263), .out0(new_n265));
  inv000aa1n02x5               g170(.a(new_n228), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n263), .b(new_n266), .c(new_n225), .d(new_n221), .o1(new_n267));
  nanb02aa1n06x5               g172(.a(new_n258), .b(new_n254), .out0(new_n268));
  inv000aa1d42x5               g173(.a(\a[24] ), .o1(new_n269));
  inv000aa1d42x5               g174(.a(\b[23] ), .o1(new_n270));
  oao003aa1n02x5               g175(.a(new_n269), .b(new_n270), .c(new_n257), .carry(new_n271));
  inv040aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n268), .c(new_n267), .d(new_n251), .o1(new_n273));
  inv000aa1n02x5               g178(.a(new_n273), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n265), .c(new_n182), .d(new_n191), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  xnrc02aa1n12x5               g183(.a(\b[25] ), .b(\a[26] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  nand42aa1n02x5               g185(.a(new_n275), .b(new_n278), .o1(new_n281));
  nona22aa1n03x5               g186(.a(new_n281), .b(new_n279), .c(new_n277), .out0(new_n282));
  nanp02aa1n03x5               g187(.a(new_n282), .b(new_n280), .o1(\s[26] ));
  norb02aa1n12x5               g188(.a(new_n278), .b(new_n279), .out0(new_n284));
  nano23aa1n06x5               g189(.a(new_n226), .b(new_n268), .c(new_n284), .d(new_n263), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n197), .c(new_n132), .d(new_n181), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n284), .b(new_n271), .c(new_n252), .d(new_n264), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\a[26] ), .o1(new_n288));
  inv000aa1d42x5               g193(.a(\b[25] ), .o1(new_n289));
  oao003aa1n02x5               g194(.a(new_n288), .b(new_n289), .c(new_n277), .carry(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  nanp03aa1n03x5               g196(.a(new_n286), .b(new_n287), .c(new_n291), .o1(new_n292));
  xorc02aa1n12x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  aoi112aa1n02x5               g198(.a(new_n293), .b(new_n290), .c(new_n273), .d(new_n284), .o1(new_n294));
  aoi022aa1n02x5               g199(.a(new_n292), .b(new_n293), .c(new_n294), .d(new_n286), .o1(\s[27] ));
  nor042aa1n03x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  xnrc02aa1n12x5               g201(.a(\b[27] ), .b(\a[28] ), .out0(new_n297));
  aoai13aa1n03x5               g202(.a(new_n297), .b(new_n296), .c(new_n292), .d(new_n293), .o1(new_n298));
  nona23aa1n09x5               g203(.a(new_n234), .b(new_n284), .c(new_n243), .d(new_n268), .out0(new_n299));
  oaoi13aa1n09x5               g204(.a(new_n299), .b(new_n191), .c(new_n124), .d(new_n219), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n264), .b(new_n250), .c(new_n229), .d(new_n263), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n284), .o1(new_n302));
  aoai13aa1n06x5               g207(.a(new_n291), .b(new_n302), .c(new_n301), .d(new_n272), .o1(new_n303));
  oai012aa1n03x5               g208(.a(new_n293), .b(new_n303), .c(new_n300), .o1(new_n304));
  nona22aa1n03x5               g209(.a(new_n304), .b(new_n297), .c(new_n296), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n298), .b(new_n305), .o1(\s[28] ));
  norb02aa1n03x5               g211(.a(new_n293), .b(new_n297), .out0(new_n307));
  tech160nm_fioai012aa1n04x5   g212(.a(new_n307), .b(new_n303), .c(new_n300), .o1(new_n308));
  xorc02aa1n12x5               g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  inv000aa1d42x5               g214(.a(\a[28] ), .o1(new_n310));
  inv000aa1d42x5               g215(.a(\b[27] ), .o1(new_n311));
  aoi112aa1n02x5               g216(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n312));
  aoi112aa1n02x5               g217(.a(new_n309), .b(new_n312), .c(new_n310), .d(new_n311), .o1(new_n313));
  aoi012aa1n03x5               g218(.a(new_n290), .b(new_n273), .c(new_n284), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n307), .o1(new_n315));
  oao003aa1n06x5               g220(.a(new_n310), .b(new_n311), .c(new_n296), .carry(new_n316));
  inv000aa1d42x5               g221(.a(new_n316), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n315), .c(new_n314), .d(new_n286), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n318), .b(new_n309), .c(new_n308), .d(new_n313), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g225(.a(new_n297), .b(new_n293), .c(new_n309), .out0(new_n321));
  oai012aa1n03x5               g226(.a(new_n321), .b(new_n303), .c(new_n300), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  inv000aa1d42x5               g228(.a(\a[29] ), .o1(new_n324));
  inv000aa1d42x5               g229(.a(\b[28] ), .o1(new_n325));
  oabi12aa1n02x5               g230(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n326));
  oaoi13aa1n02x5               g231(.a(new_n326), .b(new_n316), .c(new_n324), .d(new_n325), .o1(new_n327));
  inv000aa1n02x5               g232(.a(new_n321), .o1(new_n328));
  tech160nm_fioaoi03aa1n03p5x5 g233(.a(new_n324), .b(new_n325), .c(new_n316), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n328), .c(new_n314), .d(new_n286), .o1(new_n330));
  aoi022aa1n03x5               g235(.a(new_n330), .b(new_n323), .c(new_n322), .d(new_n327), .o1(\s[30] ));
  nand03aa1n02x5               g236(.a(new_n307), .b(new_n309), .c(new_n323), .o1(new_n332));
  oabi12aa1n03x5               g237(.a(new_n332), .b(new_n303), .c(new_n300), .out0(new_n333));
  xorc02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  oao003aa1n03x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n329), .carry(new_n335));
  norb02aa1n03x4               g240(.a(new_n335), .b(new_n334), .out0(new_n336));
  aoai13aa1n03x5               g241(.a(new_n335), .b(new_n332), .c(new_n314), .d(new_n286), .o1(new_n337));
  aoi022aa1n03x5               g242(.a(new_n337), .b(new_n334), .c(new_n333), .d(new_n336), .o1(\s[31] ));
  xnbna2aa1n03x5               g243(.a(new_n118), .b(new_n112), .c(new_n113), .out0(\s[3] ));
  orn002aa1n02x5               g244(.a(new_n118), .b(new_n114), .o(new_n340));
  xorc02aa1n02x5               g245(.a(\a[4] ), .b(\b[3] ), .out0(new_n341));
  norb02aa1n02x5               g246(.a(new_n112), .b(new_n341), .out0(new_n342));
  aoi022aa1n02x5               g247(.a(new_n340), .b(new_n342), .c(new_n119), .d(new_n341), .o1(\s[4] ));
  nano22aa1n02x4               g248(.a(new_n105), .b(new_n120), .c(new_n121), .out0(new_n344));
  nanb02aa1n02x5               g249(.a(new_n105), .b(new_n120), .out0(new_n345));
  nanp02aa1n02x5               g250(.a(new_n119), .b(new_n121), .o1(new_n346));
  aoi022aa1n02x5               g251(.a(new_n346), .b(new_n345), .c(new_n119), .d(new_n344), .o1(\s[5] ));
  aoi012aa1n02x5               g252(.a(new_n105), .b(new_n119), .c(new_n344), .o1(new_n348));
  xnrb03aa1n02x5               g253(.a(new_n348), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aob012aa1n02x5               g254(.a(new_n106), .b(new_n119), .c(new_n123), .out0(new_n350));
  xorb03aa1n02x5               g255(.a(new_n350), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g256(.a(new_n99), .b(new_n350), .c(new_n100), .o1(new_n352));
  xnrb03aa1n02x5               g257(.a(new_n352), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g258(.a(new_n134), .b(new_n131), .c(new_n130), .out0(\s[9] ));
endmodule


