// Benchmark "adder" written by ABC on Thu Jul 18 03:39:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n172, new_n173, new_n174, new_n175, new_n176, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n350, new_n351,
    new_n353, new_n354, new_n356, new_n357, new_n358, new_n360, new_n361,
    new_n362, new_n364, new_n366, new_n367, new_n369;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1n06x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nor042aa1n09x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n09x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor042aa1d18x5               g006(.a(new_n100), .b(new_n101), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nor042aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb03aa1n12x5               g009(.a(new_n104), .b(new_n99), .c(new_n103), .out0(new_n105));
  oab012aa1n04x5               g010(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .out0(new_n106));
  aoai13aa1n12x5               g011(.a(new_n106), .b(new_n105), .c(new_n99), .d(new_n102), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[5] ), .o1(new_n108));
  nanb02aa1n12x5               g013(.a(\a[6] ), .b(new_n108), .out0(new_n109));
  nanp02aa1n04x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  oai112aa1n03x5               g015(.a(new_n109), .b(new_n110), .c(\b[7] ), .d(\a[8] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  oai012aa1n02x5               g017(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .o1(new_n113));
  aoi022aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nor042aa1d18x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  inv000aa1n02x5               g021(.a(new_n116), .o1(new_n117));
  nand23aa1n03x5               g022(.a(new_n114), .b(new_n117), .c(new_n115), .o1(new_n118));
  nor043aa1n03x5               g023(.a(new_n118), .b(new_n111), .c(new_n113), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[7] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[6] ), .o1(new_n121));
  norp02aa1n03x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  aoai13aa1n03x5               g027(.a(new_n112), .b(new_n122), .c(new_n120), .d(new_n121), .o1(new_n123));
  oai122aa1n06x5               g028(.a(new_n110), .b(new_n120), .c(new_n121), .d(\a[8] ), .e(\b[7] ), .o1(new_n124));
  nor042aa1n02x5               g029(.a(\b[5] ), .b(\a[6] ), .o1(new_n125));
  nanp02aa1n02x5               g030(.a(new_n121), .b(new_n120), .o1(new_n126));
  oai112aa1n04x5               g031(.a(new_n126), .b(new_n112), .c(new_n125), .d(new_n116), .o1(new_n127));
  oai012aa1n12x5               g032(.a(new_n123), .b(new_n127), .c(new_n124), .o1(new_n128));
  xnrc02aa1n12x5               g033(.a(\b[8] ), .b(\a[9] ), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n128), .c(new_n119), .d(new_n107), .o1(new_n131));
  nor042aa1n04x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nand02aa1d16x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  norb02aa1n09x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  xnbna2aa1n03x5               g039(.a(new_n134), .b(new_n131), .c(new_n98), .out0(\s[10] ));
  nano23aa1n09x5               g040(.a(new_n102), .b(new_n104), .c(new_n103), .d(new_n99), .out0(new_n136));
  oai022aa1n02x5               g041(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n137));
  oai012aa1n06x5               g042(.a(new_n119), .b(new_n136), .c(new_n137), .o1(new_n138));
  inv040aa1n02x5               g043(.a(new_n128), .o1(new_n139));
  nanp02aa1n03x5               g044(.a(new_n138), .b(new_n139), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n134), .b(new_n97), .c(new_n140), .d(new_n130), .o1(new_n141));
  oai012aa1n02x5               g046(.a(new_n133), .b(new_n132), .c(new_n97), .o1(new_n142));
  nor022aa1n06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nand02aa1n03x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n141), .c(new_n142), .out0(\s[11] ));
  inv040aa1n02x5               g051(.a(new_n134), .o1(new_n147));
  aoai13aa1n02x5               g052(.a(new_n142), .b(new_n147), .c(new_n131), .d(new_n98), .o1(new_n148));
  aoi012aa1n02x5               g053(.a(new_n143), .b(new_n148), .c(new_n144), .o1(new_n149));
  nor002aa1n06x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nand02aa1d04x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nanb02aa1n02x5               g056(.a(new_n150), .b(new_n151), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n143), .b(new_n153), .c(new_n148), .d(new_n145), .o1(new_n154));
  oab012aa1n02x4               g059(.a(new_n154), .b(new_n149), .c(new_n152), .out0(\s[12] ));
  nona23aa1n03x5               g060(.a(new_n151), .b(new_n144), .c(new_n143), .d(new_n150), .out0(new_n156));
  nor043aa1n06x5               g061(.a(new_n156), .b(new_n147), .c(new_n129), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n128), .c(new_n119), .d(new_n107), .o1(new_n158));
  nano22aa1n03x7               g063(.a(new_n150), .b(new_n144), .c(new_n151), .out0(new_n159));
  oai122aa1n03x5               g064(.a(new_n133), .b(new_n132), .c(new_n97), .d(\b[10] ), .e(\a[11] ), .o1(new_n160));
  aoi012aa1n02x7               g065(.a(new_n150), .b(new_n143), .c(new_n151), .o1(new_n161));
  oaib12aa1n09x5               g066(.a(new_n161), .b(new_n160), .c(new_n159), .out0(new_n162));
  nanb02aa1n02x5               g067(.a(new_n162), .b(new_n158), .out0(new_n163));
  nor022aa1n06x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nand02aa1n03x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  oai012aa1n02x7               g071(.a(new_n133), .b(\b[10] ), .c(\a[11] ), .o1(new_n167));
  oab012aa1n06x5               g072(.a(new_n167), .b(new_n97), .c(new_n132), .out0(new_n168));
  inv000aa1n03x5               g073(.a(new_n161), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(new_n169), .b(new_n166), .c(new_n168), .d(new_n159), .o1(new_n170));
  aoi022aa1n02x5               g075(.a(new_n163), .b(new_n166), .c(new_n158), .d(new_n170), .o1(\s[13] ));
  nor022aa1n04x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nand42aa1n02x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n174), .b(new_n164), .c(new_n163), .d(new_n165), .o1(new_n175));
  aoi112aa1n02x5               g080(.a(new_n164), .b(new_n174), .c(new_n163), .d(new_n166), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n175), .b(new_n176), .out0(\s[14] ));
  nano23aa1n06x5               g082(.a(new_n164), .b(new_n172), .c(new_n173), .d(new_n165), .out0(new_n178));
  aoai13aa1n03x5               g083(.a(new_n178), .b(new_n162), .c(new_n140), .d(new_n157), .o1(new_n179));
  oaih12aa1n02x5               g084(.a(new_n173), .b(new_n172), .c(new_n164), .o1(new_n180));
  nor002aa1n20x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  nanp02aa1n04x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nanb02aa1n02x5               g087(.a(new_n181), .b(new_n182), .out0(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n179), .c(new_n180), .out0(\s[15] ));
  inv000aa1n02x5               g090(.a(new_n180), .o1(new_n186));
  aoai13aa1n02x5               g091(.a(new_n184), .b(new_n186), .c(new_n163), .d(new_n178), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n181), .o1(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n183), .c(new_n179), .d(new_n180), .o1(new_n189));
  nor002aa1n06x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nand02aa1n04x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  nanb02aa1n02x5               g096(.a(new_n190), .b(new_n191), .out0(new_n192));
  aoib12aa1n02x5               g097(.a(new_n181), .b(new_n191), .c(new_n190), .out0(new_n193));
  aboi22aa1n03x5               g098(.a(new_n192), .b(new_n189), .c(new_n193), .d(new_n187), .out0(\s[16] ));
  nona23aa1n02x4               g099(.a(new_n173), .b(new_n165), .c(new_n164), .d(new_n172), .out0(new_n195));
  nona23aa1d24x5               g100(.a(new_n191), .b(new_n182), .c(new_n181), .d(new_n190), .out0(new_n196));
  nona22aa1n09x5               g101(.a(new_n157), .b(new_n195), .c(new_n196), .out0(new_n197));
  aoi012aa1d18x5               g102(.a(new_n197), .b(new_n138), .c(new_n139), .o1(new_n198));
  aoai13aa1n04x5               g103(.a(new_n178), .b(new_n169), .c(new_n168), .d(new_n159), .o1(new_n199));
  tech160nm_fiaoi012aa1n03p5x5 g104(.a(new_n190), .b(new_n181), .c(new_n191), .o1(new_n200));
  aoai13aa1n12x5               g105(.a(new_n200), .b(new_n196), .c(new_n199), .d(new_n180), .o1(new_n201));
  tech160nm_fixorc02aa1n02p5x5 g106(.a(\a[17] ), .b(\b[16] ), .out0(new_n202));
  tech160nm_fioai012aa1n03p5x5 g107(.a(new_n202), .b(new_n201), .c(new_n198), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n196), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n186), .c(new_n162), .d(new_n178), .o1(new_n205));
  nano23aa1n02x4               g110(.a(new_n202), .b(new_n198), .c(new_n205), .d(new_n200), .out0(new_n206));
  norb02aa1n02x5               g111(.a(new_n203), .b(new_n206), .out0(\s[17] ));
  nor002aa1d32x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  nor042aa1n06x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nand02aa1d08x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  norb02aa1n06x4               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n203), .c(new_n209), .out0(\s[18] ));
  and002aa1n02x5               g118(.a(new_n202), .b(new_n212), .o(new_n214));
  tech160nm_fioai012aa1n03p5x5 g119(.a(new_n214), .b(new_n201), .c(new_n198), .o1(new_n215));
  oaoi03aa1n02x5               g120(.a(\a[18] ), .b(\b[17] ), .c(new_n209), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  nor042aa1d18x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nand02aa1n06x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  norb02aa1n06x4               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  xnbna2aa1n03x5               g125(.a(new_n220), .b(new_n215), .c(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g126(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoi012aa1n06x5               g127(.a(new_n128), .b(new_n119), .c(new_n107), .o1(new_n223));
  oai112aa1n06x5               g128(.a(new_n205), .b(new_n200), .c(new_n197), .d(new_n223), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n220), .b(new_n216), .c(new_n224), .d(new_n214), .o1(new_n225));
  inv040aa1n02x5               g130(.a(new_n218), .o1(new_n226));
  inv000aa1n03x5               g131(.a(new_n220), .o1(new_n227));
  aoai13aa1n02x5               g132(.a(new_n226), .b(new_n227), .c(new_n215), .d(new_n217), .o1(new_n228));
  nor042aa1n06x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  nand02aa1d28x5               g134(.a(\b[19] ), .b(\a[20] ), .o1(new_n230));
  norb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  inv000aa1d42x5               g136(.a(\a[19] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\b[18] ), .o1(new_n233));
  aboi22aa1n03x5               g138(.a(new_n229), .b(new_n230), .c(new_n232), .d(new_n233), .out0(new_n234));
  aoi022aa1n03x5               g139(.a(new_n228), .b(new_n231), .c(new_n225), .d(new_n234), .o1(\s[20] ));
  nano32aa1n03x7               g140(.a(new_n227), .b(new_n202), .c(new_n231), .d(new_n212), .out0(new_n236));
  oaih12aa1n02x5               g141(.a(new_n236), .b(new_n201), .c(new_n198), .o1(new_n237));
  nanb03aa1n09x5               g142(.a(new_n229), .b(new_n230), .c(new_n219), .out0(new_n238));
  oai112aa1n06x5               g143(.a(new_n226), .b(new_n211), .c(new_n210), .d(new_n208), .o1(new_n239));
  aoi012aa1n06x5               g144(.a(new_n229), .b(new_n218), .c(new_n230), .o1(new_n240));
  oaih12aa1n12x5               g145(.a(new_n240), .b(new_n239), .c(new_n238), .o1(new_n241));
  xnrc02aa1n12x5               g146(.a(\b[20] ), .b(\a[21] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n241), .c(new_n224), .d(new_n236), .o1(new_n244));
  nano22aa1n02x4               g149(.a(new_n229), .b(new_n219), .c(new_n230), .out0(new_n245));
  oai012aa1n02x5               g150(.a(new_n211), .b(\b[18] ), .c(\a[19] ), .o1(new_n246));
  oab012aa1n02x5               g151(.a(new_n246), .b(new_n208), .c(new_n210), .out0(new_n247));
  inv020aa1n02x5               g152(.a(new_n240), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n243), .b(new_n248), .c(new_n247), .d(new_n245), .o1(new_n249));
  aobi12aa1n03x7               g154(.a(new_n244), .b(new_n249), .c(new_n237), .out0(\s[21] ));
  inv000aa1d42x5               g155(.a(new_n241), .o1(new_n251));
  nor042aa1n06x5               g156(.a(\b[20] ), .b(\a[21] ), .o1(new_n252));
  inv000aa1n06x5               g157(.a(new_n252), .o1(new_n253));
  aoai13aa1n02x7               g158(.a(new_n253), .b(new_n242), .c(new_n237), .d(new_n251), .o1(new_n254));
  xnrc02aa1n12x5               g159(.a(\b[21] ), .b(\a[22] ), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n255), .b(new_n252), .out0(new_n257));
  aoi022aa1n03x5               g162(.a(new_n254), .b(new_n256), .c(new_n244), .d(new_n257), .o1(\s[22] ));
  nor042aa1n06x5               g163(.a(new_n255), .b(new_n242), .o1(new_n259));
  and002aa1n02x5               g164(.a(new_n236), .b(new_n259), .o(new_n260));
  oaih12aa1n02x5               g165(.a(new_n260), .b(new_n201), .c(new_n198), .o1(new_n261));
  oao003aa1n06x5               g166(.a(\a[22] ), .b(\b[21] ), .c(new_n253), .carry(new_n262));
  inv040aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  aoi012aa1d18x5               g168(.a(new_n263), .b(new_n241), .c(new_n259), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n12x5               g170(.a(\a[23] ), .b(\b[22] ), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n265), .c(new_n224), .d(new_n260), .o1(new_n267));
  aoi112aa1n02x5               g172(.a(new_n266), .b(new_n263), .c(new_n241), .d(new_n259), .o1(new_n268));
  aobi12aa1n02x7               g173(.a(new_n267), .b(new_n268), .c(new_n261), .out0(\s[23] ));
  nor042aa1n06x5               g174(.a(\b[22] ), .b(\a[23] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n266), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n271), .b(new_n272), .c(new_n261), .d(new_n264), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[24] ), .b(\b[23] ), .out0(new_n274));
  norp02aa1n02x5               g179(.a(new_n274), .b(new_n270), .o1(new_n275));
  aoi022aa1n02x7               g180(.a(new_n273), .b(new_n274), .c(new_n267), .d(new_n275), .o1(\s[24] ));
  inv000aa1n02x5               g181(.a(new_n236), .o1(new_n277));
  and002aa1n06x5               g182(.a(new_n274), .b(new_n266), .o(new_n278));
  nano22aa1n02x4               g183(.a(new_n277), .b(new_n278), .c(new_n259), .out0(new_n279));
  oaih12aa1n02x5               g184(.a(new_n279), .b(new_n201), .c(new_n198), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n259), .b(new_n248), .c(new_n247), .d(new_n245), .o1(new_n281));
  inv000aa1n02x5               g186(.a(new_n278), .o1(new_n282));
  oao003aa1n02x5               g187(.a(\a[24] ), .b(\b[23] ), .c(new_n271), .carry(new_n283));
  aoai13aa1n12x5               g188(.a(new_n283), .b(new_n282), .c(new_n281), .d(new_n262), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n284), .c(new_n224), .d(new_n279), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n278), .b(new_n263), .c(new_n241), .d(new_n259), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  and003aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n283), .o(new_n289));
  aobi12aa1n03x7               g194(.a(new_n286), .b(new_n289), .c(new_n280), .out0(\s[25] ));
  inv000aa1d42x5               g195(.a(new_n284), .o1(new_n291));
  nor042aa1n03x5               g196(.a(\b[24] ), .b(\a[25] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n288), .c(new_n280), .d(new_n291), .o1(new_n294));
  xorc02aa1n02x5               g199(.a(\a[26] ), .b(\b[25] ), .out0(new_n295));
  norp02aa1n02x5               g200(.a(new_n295), .b(new_n292), .o1(new_n296));
  aoi022aa1n03x5               g201(.a(new_n294), .b(new_n295), .c(new_n286), .d(new_n296), .o1(\s[26] ));
  and002aa1n02x7               g202(.a(new_n295), .b(new_n285), .o(new_n298));
  nano32aa1n03x7               g203(.a(new_n277), .b(new_n298), .c(new_n259), .d(new_n278), .out0(new_n299));
  tech160nm_fioai012aa1n03p5x5 g204(.a(new_n299), .b(new_n201), .c(new_n198), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n298), .o1(new_n301));
  oao003aa1n02x5               g206(.a(\a[26] ), .b(\b[25] ), .c(new_n293), .carry(new_n302));
  aoai13aa1n04x5               g207(.a(new_n302), .b(new_n301), .c(new_n287), .d(new_n283), .o1(new_n303));
  xorc02aa1n12x5               g208(.a(\a[27] ), .b(\b[26] ), .out0(new_n304));
  aoai13aa1n06x5               g209(.a(new_n304), .b(new_n303), .c(new_n224), .d(new_n299), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n302), .o1(new_n306));
  aoi112aa1n02x5               g211(.a(new_n304), .b(new_n306), .c(new_n284), .d(new_n298), .o1(new_n307));
  aobi12aa1n02x7               g212(.a(new_n305), .b(new_n307), .c(new_n300), .out0(\s[27] ));
  aoi012aa1n09x5               g213(.a(new_n306), .b(new_n284), .c(new_n298), .o1(new_n309));
  norp02aa1n02x5               g214(.a(\b[26] ), .b(\a[27] ), .o1(new_n310));
  inv000aa1n03x5               g215(.a(new_n310), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n304), .o1(new_n312));
  aoai13aa1n03x5               g217(.a(new_n311), .b(new_n312), .c(new_n309), .d(new_n300), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[28] ), .b(\b[27] ), .out0(new_n314));
  norp02aa1n02x5               g219(.a(new_n314), .b(new_n310), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n305), .d(new_n315), .o1(\s[28] ));
  and002aa1n02x5               g221(.a(new_n314), .b(new_n304), .o(new_n317));
  aoai13aa1n02x5               g222(.a(new_n317), .b(new_n303), .c(new_n224), .d(new_n299), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[28] ), .b(\b[27] ), .c(new_n311), .carry(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n309), .d(new_n300), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n320), .b(new_n322), .out0(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g230(.a(new_n312), .b(new_n314), .c(new_n322), .out0(new_n326));
  aoai13aa1n06x5               g231(.a(new_n326), .b(new_n303), .c(new_n224), .d(new_n299), .o1(new_n327));
  inv000aa1n02x5               g232(.a(new_n326), .o1(new_n328));
  inv000aa1d42x5               g233(.a(\b[28] ), .o1(new_n329));
  inv000aa1d42x5               g234(.a(\a[29] ), .o1(new_n330));
  oaib12aa1n02x5               g235(.a(new_n320), .b(\b[28] ), .c(new_n330), .out0(new_n331));
  oaib12aa1n02x5               g236(.a(new_n331), .b(new_n329), .c(\a[29] ), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n328), .c(new_n309), .d(new_n300), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[30] ), .b(\b[29] ), .out0(new_n334));
  oaoi13aa1n02x5               g239(.a(new_n334), .b(new_n331), .c(new_n330), .d(new_n329), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n333), .b(new_n334), .c(new_n327), .d(new_n335), .o1(\s[30] ));
  nanb02aa1n02x5               g241(.a(\b[30] ), .b(\a[31] ), .out0(new_n337));
  nanb02aa1n02x5               g242(.a(\a[31] ), .b(\b[30] ), .out0(new_n338));
  nanp02aa1n02x5               g243(.a(new_n338), .b(new_n337), .o1(new_n339));
  nano32aa1n06x5               g244(.a(new_n312), .b(new_n334), .c(new_n314), .d(new_n322), .out0(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n303), .c(new_n224), .d(new_n299), .o1(new_n341));
  inv000aa1d42x5               g246(.a(new_n340), .o1(new_n342));
  norp02aa1n02x5               g247(.a(\b[29] ), .b(\a[30] ), .o1(new_n343));
  aoi022aa1n02x5               g248(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n344));
  aoi012aa1n02x5               g249(.a(new_n343), .b(new_n331), .c(new_n344), .o1(new_n345));
  aoai13aa1n03x5               g250(.a(new_n345), .b(new_n342), .c(new_n309), .d(new_n300), .o1(new_n346));
  oai112aa1n02x5               g251(.a(new_n337), .b(new_n338), .c(\b[29] ), .d(\a[30] ), .o1(new_n347));
  aoi012aa1n02x5               g252(.a(new_n347), .b(new_n331), .c(new_n344), .o1(new_n348));
  aoi022aa1n03x5               g253(.a(new_n346), .b(new_n339), .c(new_n341), .d(new_n348), .o1(\s[31] ));
  inv000aa1d42x5               g254(.a(new_n102), .o1(new_n350));
  aboi22aa1n03x5               g255(.a(new_n104), .b(new_n103), .c(new_n350), .d(new_n99), .out0(new_n351));
  norp02aa1n02x5               g256(.a(new_n351), .b(new_n136), .o1(\s[3] ));
  xorc02aa1n02x5               g257(.a(\a[4] ), .b(\b[3] ), .out0(new_n353));
  norp02aa1n02x5               g258(.a(new_n353), .b(new_n104), .o1(new_n354));
  aboi22aa1n03x5               g259(.a(new_n136), .b(new_n354), .c(new_n107), .d(new_n353), .out0(\s[4] ));
  aoi022aa1n02x5               g260(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n356));
  and002aa1n02x5               g261(.a(\b[3] ), .b(\a[4] ), .o(new_n357));
  aboi22aa1n03x5               g262(.a(new_n357), .b(new_n107), .c(new_n117), .d(new_n115), .out0(new_n358));
  aoi013aa1n02x4               g263(.a(new_n358), .b(new_n356), .c(new_n117), .d(new_n107), .o1(\s[5] ));
  norb02aa1n02x5               g264(.a(new_n110), .b(new_n125), .out0(new_n360));
  aoai13aa1n02x5               g265(.a(new_n360), .b(new_n116), .c(new_n107), .d(new_n356), .o1(new_n361));
  aoi112aa1n02x5               g266(.a(new_n116), .b(new_n360), .c(new_n107), .d(new_n356), .o1(new_n362));
  norb02aa1n02x5               g267(.a(new_n361), .b(new_n362), .out0(\s[6] ));
  xorc02aa1n02x5               g268(.a(\a[7] ), .b(\b[6] ), .out0(new_n364));
  xnbna2aa1n03x5               g269(.a(new_n364), .b(new_n361), .c(new_n109), .out0(\s[7] ));
  aob012aa1n02x5               g270(.a(new_n364), .b(new_n361), .c(new_n109), .out0(new_n366));
  norb02aa1n02x5               g271(.a(new_n112), .b(new_n122), .out0(new_n367));
  xnbna2aa1n03x5               g272(.a(new_n367), .b(new_n366), .c(new_n126), .out0(\s[8] ));
  oai112aa1n02x5               g273(.a(new_n123), .b(new_n129), .c(new_n127), .d(new_n124), .o1(new_n369));
  aboi22aa1n03x5               g274(.a(new_n369), .b(new_n138), .c(new_n140), .d(new_n130), .out0(\s[9] ));
endmodule


