// Benchmark "adder" written by ABC on Thu Jul 18 02:46:48 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n247, new_n248, new_n249, new_n250, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n323, new_n326,
    new_n327, new_n328, new_n330, new_n331, new_n332, new_n333, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  nand42aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nor042aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oaih12aa1n06x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  nor022aa1n08x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n09x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n104), .b(new_n103), .c(new_n105), .d(new_n102), .out0(new_n106));
  tech160nm_fiaoi012aa1n03p5x5 g011(.a(new_n105), .b(new_n102), .c(new_n104), .o1(new_n107));
  oai012aa1n12x5               g012(.a(new_n107), .b(new_n106), .c(new_n101), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\a[6] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\b[5] ), .o1(new_n111));
  norp02aa1n12x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  aoi012aa1n02x5               g017(.a(new_n112), .b(new_n110), .c(new_n111), .o1(new_n113));
  nor042aa1n06x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nor042aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nona23aa1n09x5               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nanp02aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano32aa1n03x7               g024(.a(new_n118), .b(new_n113), .c(new_n109), .d(new_n119), .out0(new_n120));
  oaoi03aa1n02x5               g025(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n121));
  oai012aa1n02x5               g026(.a(new_n116), .b(new_n117), .c(new_n114), .o1(new_n122));
  oai012aa1n06x5               g027(.a(new_n122), .b(new_n118), .c(new_n121), .o1(new_n123));
  nor042aa1d18x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nand42aa1n08x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  aoai13aa1n03x5               g031(.a(new_n126), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n127));
  nor042aa1d18x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand02aa1d28x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n06x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n97), .out0(\s[10] ));
  nor002aa1d32x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand02aa1n12x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nanb02aa1n02x5               g038(.a(new_n132), .b(new_n133), .out0(new_n134));
  nona22aa1n02x4               g039(.a(new_n127), .b(new_n128), .c(new_n124), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n134), .b(new_n135), .c(new_n129), .out0(\s[11] ));
  aoi013aa1n02x4               g041(.a(new_n132), .b(new_n135), .c(new_n133), .d(new_n129), .o1(new_n137));
  xnrb03aa1n03x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norb03aa1n12x5               g043(.a(new_n125), .b(new_n124), .c(new_n132), .out0(new_n139));
  nor002aa1d32x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nano22aa1n12x5               g046(.a(new_n140), .b(new_n133), .c(new_n141), .out0(new_n142));
  nand23aa1d12x5               g047(.a(new_n142), .b(new_n139), .c(new_n130), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n143), .o1(new_n144));
  aoai13aa1n03x5               g049(.a(new_n144), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n145));
  nanb03aa1n12x5               g050(.a(new_n140), .b(new_n141), .c(new_n133), .out0(new_n146));
  inv020aa1n06x5               g051(.a(new_n132), .o1(new_n147));
  oai112aa1n06x5               g052(.a(new_n147), .b(new_n129), .c(new_n128), .d(new_n124), .o1(new_n148));
  oai012aa1d24x5               g053(.a(new_n141), .b(new_n140), .c(new_n132), .o1(new_n149));
  oai012aa1n18x5               g054(.a(new_n149), .b(new_n148), .c(new_n146), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n145), .b(new_n151), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n09x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand42aa1d28x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n154), .b(new_n152), .c(new_n155), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand42aa1d28x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nano23aa1d15x5               g064(.a(new_n154), .b(new_n158), .c(new_n159), .d(new_n155), .out0(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoi012aa1d18x5               g066(.a(new_n158), .b(new_n154), .c(new_n159), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n161), .c(new_n145), .d(new_n151), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n09x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand42aa1d28x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nor042aa1n06x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nand42aa1d28x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  aoai13aa1n03x5               g074(.a(new_n169), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n165), .b(new_n169), .c(new_n163), .d(new_n166), .o1(new_n171));
  norb02aa1n03x4               g076(.a(new_n170), .b(new_n171), .out0(\s[16] ));
  nano23aa1d15x5               g077(.a(new_n165), .b(new_n167), .c(new_n168), .d(new_n166), .out0(new_n173));
  nano22aa1d15x5               g078(.a(new_n143), .b(new_n160), .c(new_n173), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n123), .c(new_n108), .d(new_n120), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n162), .o1(new_n176));
  aoai13aa1n09x5               g081(.a(new_n173), .b(new_n176), .c(new_n150), .d(new_n160), .o1(new_n177));
  oai012aa1n18x5               g082(.a(new_n168), .b(new_n167), .c(new_n165), .o1(new_n178));
  nand23aa1n06x5               g083(.a(new_n175), .b(new_n177), .c(new_n178), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  inv030aa1d32x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n03x5               g088(.a(new_n182), .b(new_n183), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  inv040aa1n02x5               g090(.a(new_n123), .o1(new_n186));
  aob012aa1d15x5               g091(.a(new_n186), .b(new_n108), .c(new_n120), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n173), .o1(new_n188));
  oai012aa1n02x5               g093(.a(new_n129), .b(\b[10] ), .c(\a[11] ), .o1(new_n189));
  oab012aa1n02x4               g094(.a(new_n189), .b(new_n124), .c(new_n128), .out0(new_n190));
  inv000aa1d42x5               g095(.a(new_n149), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n160), .b(new_n191), .c(new_n190), .d(new_n142), .o1(new_n192));
  aoai13aa1n09x5               g097(.a(new_n178), .b(new_n188), .c(new_n192), .d(new_n162), .o1(new_n193));
  xroi22aa1d06x4               g098(.a(new_n182), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n193), .c(new_n187), .d(new_n174), .o1(new_n195));
  nor042aa1d18x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nor042aa1n06x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  nand02aa1d28x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  aoi012aa1d24x5               g103(.a(new_n197), .b(new_n196), .c(new_n198), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\a[19] ), .o1(new_n200));
  nanb02aa1d36x5               g105(.a(\b[18] ), .b(new_n200), .out0(new_n201));
  nanp02aa1n02x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand22aa1n04x5               g107(.a(new_n201), .b(new_n202), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n195), .c(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g111(.a(new_n199), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n204), .b(new_n207), .c(new_n179), .d(new_n194), .o1(new_n208));
  xnrc02aa1n02x5               g113(.a(\b[19] ), .b(\a[20] ), .out0(new_n209));
  aoi012aa1n02x7               g114(.a(new_n209), .b(new_n208), .c(new_n201), .o1(new_n210));
  tech160nm_fiaoi012aa1n03p5x5 g115(.a(new_n203), .b(new_n195), .c(new_n199), .o1(new_n211));
  nano22aa1n03x7               g116(.a(new_n211), .b(new_n201), .c(new_n209), .out0(new_n212));
  nor002aa1n02x5               g117(.a(new_n210), .b(new_n212), .o1(\s[20] ));
  nona22aa1d18x5               g118(.a(new_n194), .b(new_n203), .c(new_n209), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n193), .c(new_n187), .d(new_n174), .o1(new_n216));
  inv000aa1d42x5               g121(.a(\b[19] ), .o1(new_n217));
  oa0022aa1n12x5               g122(.a(\a[20] ), .b(\b[19] ), .c(\a[19] ), .d(\b[18] ), .o(new_n218));
  aoai13aa1n12x5               g123(.a(new_n218), .b(new_n199), .c(\a[19] ), .d(\b[18] ), .o1(new_n219));
  oaib12aa1n12x5               g124(.a(new_n219), .b(new_n217), .c(\a[20] ), .out0(new_n220));
  nor002aa1d32x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  tech160nm_finand02aa1n05x5   g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n216), .c(new_n220), .out0(\s[21] ));
  inv020aa1n02x5               g129(.a(new_n221), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n220), .o1(new_n226));
  aoai13aa1n03x5               g131(.a(new_n223), .b(new_n226), .c(new_n179), .d(new_n215), .o1(new_n227));
  nor022aa1n16x5               g132(.a(\b[21] ), .b(\a[22] ), .o1(new_n228));
  nand42aa1n04x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  nanb02aa1n02x5               g134(.a(new_n228), .b(new_n229), .out0(new_n230));
  tech160nm_fiaoi012aa1n02p5x5 g135(.a(new_n230), .b(new_n227), .c(new_n225), .o1(new_n231));
  inv000aa1n02x5               g136(.a(new_n223), .o1(new_n232));
  aoi012aa1n03x5               g137(.a(new_n232), .b(new_n216), .c(new_n220), .o1(new_n233));
  nano22aa1n02x4               g138(.a(new_n233), .b(new_n225), .c(new_n230), .out0(new_n234));
  norp02aa1n03x5               g139(.a(new_n231), .b(new_n234), .o1(\s[22] ));
  xnrc02aa1n12x5               g140(.a(\b[22] ), .b(\a[23] ), .out0(new_n236));
  nona23aa1d24x5               g141(.a(new_n229), .b(new_n222), .c(new_n221), .d(new_n228), .out0(new_n237));
  nor042aa1n03x5               g142(.a(new_n214), .b(new_n237), .o1(new_n238));
  oaoi03aa1n03x5               g143(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .o1(new_n239));
  oabi12aa1n06x5               g144(.a(new_n239), .b(new_n220), .c(new_n237), .out0(new_n240));
  aoai13aa1n02x5               g145(.a(new_n236), .b(new_n240), .c(new_n179), .d(new_n238), .o1(new_n241));
  norp02aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  and002aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o(new_n243));
  aoai13aa1n03x5               g148(.a(new_n238), .b(new_n193), .c(new_n187), .d(new_n174), .o1(new_n244));
  nona32aa1n03x5               g149(.a(new_n244), .b(new_n240), .c(new_n243), .d(new_n242), .out0(new_n245));
  nanp02aa1n02x5               g150(.a(new_n241), .b(new_n245), .o1(\s[23] ));
  aoi112aa1n03x5               g151(.a(new_n236), .b(new_n240), .c(new_n179), .d(new_n238), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[24] ), .b(\b[23] ), .out0(new_n248));
  oai012aa1n03x5               g153(.a(new_n248), .b(new_n247), .c(new_n243), .o1(new_n249));
  nona22aa1n03x5               g154(.a(new_n245), .b(new_n248), .c(new_n243), .out0(new_n250));
  nanp02aa1n03x5               g155(.a(new_n249), .b(new_n250), .o1(\s[24] ));
  inv000aa1d42x5               g156(.a(new_n237), .o1(new_n252));
  norb02aa1n12x5               g157(.a(new_n248), .b(new_n236), .out0(new_n253));
  nano22aa1n03x7               g158(.a(new_n214), .b(new_n253), .c(new_n252), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n193), .c(new_n187), .d(new_n174), .o1(new_n255));
  and002aa1n02x5               g160(.a(\b[19] ), .b(\a[20] ), .o(new_n256));
  nona23aa1d18x5               g161(.a(new_n253), .b(new_n219), .c(new_n256), .d(new_n237), .out0(new_n257));
  aob012aa1n02x5               g162(.a(new_n242), .b(\b[23] ), .c(\a[24] ), .out0(new_n258));
  oai012aa1n02x5               g163(.a(new_n258), .b(\b[23] ), .c(\a[24] ), .o1(new_n259));
  aoi012aa1n12x5               g164(.a(new_n259), .b(new_n253), .c(new_n239), .o1(new_n260));
  nand02aa1d16x5               g165(.a(new_n260), .b(new_n257), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  xnrc02aa1n12x5               g167(.a(\b[24] ), .b(\a[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n255), .c(new_n262), .out0(\s[25] ));
  norp02aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n264), .b(new_n261), .c(new_n179), .d(new_n254), .o1(new_n268));
  xnrc02aa1n12x5               g173(.a(\b[25] ), .b(\a[26] ), .out0(new_n269));
  tech160nm_fiaoi012aa1n02p5x5 g174(.a(new_n269), .b(new_n268), .c(new_n267), .o1(new_n270));
  tech160nm_fiaoi012aa1n03p5x5 g175(.a(new_n263), .b(new_n255), .c(new_n262), .o1(new_n271));
  nano22aa1n02x4               g176(.a(new_n271), .b(new_n267), .c(new_n269), .out0(new_n272));
  norp02aa1n03x5               g177(.a(new_n270), .b(new_n272), .o1(\s[26] ));
  nor022aa1n04x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  nand42aa1n03x5               g179(.a(\b[26] ), .b(\a[27] ), .o1(new_n275));
  nanb02aa1n12x5               g180(.a(new_n274), .b(new_n275), .out0(new_n276));
  nor042aa1n09x5               g181(.a(new_n269), .b(new_n263), .o1(new_n277));
  nano32aa1d12x5               g182(.a(new_n214), .b(new_n277), .c(new_n252), .d(new_n253), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n193), .c(new_n187), .d(new_n174), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(\b[25] ), .b(\a[26] ), .o1(new_n280));
  oai022aa1n02x5               g185(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n281));
  aoi022aa1n12x5               g186(.a(new_n261), .b(new_n277), .c(new_n280), .d(new_n281), .o1(new_n282));
  xobna2aa1n03x5               g187(.a(new_n276), .b(new_n279), .c(new_n282), .out0(\s[27] ));
  xorc02aa1n12x5               g188(.a(\a[28] ), .b(\b[27] ), .out0(new_n284));
  inv000aa1d42x5               g189(.a(new_n277), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n281), .b(new_n280), .o1(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n285), .c(new_n260), .d(new_n257), .o1(new_n287));
  nona22aa1n02x5               g192(.a(new_n279), .b(new_n287), .c(new_n274), .out0(new_n288));
  aoi012aa1n03x5               g193(.a(new_n284), .b(new_n288), .c(new_n275), .o1(new_n289));
  aoi112aa1n03x4               g194(.a(new_n274), .b(new_n287), .c(new_n179), .d(new_n278), .o1(new_n290));
  nano22aa1n03x7               g195(.a(new_n290), .b(new_n275), .c(new_n284), .out0(new_n291));
  norp02aa1n03x5               g196(.a(new_n289), .b(new_n291), .o1(\s[28] ));
  norb02aa1n09x5               g197(.a(new_n284), .b(new_n276), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n293), .b(new_n287), .c(new_n179), .d(new_n278), .o1(new_n294));
  aoi112aa1n02x5               g199(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n295));
  oab012aa1n02x4               g200(.a(new_n295), .b(\a[28] ), .c(\b[27] ), .out0(new_n296));
  xnrc02aa1n12x5               g201(.a(\b[28] ), .b(\a[29] ), .out0(new_n297));
  tech160nm_fiaoi012aa1n02p5x5 g202(.a(new_n297), .b(new_n294), .c(new_n296), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n293), .o1(new_n299));
  aoi012aa1n02x7               g204(.a(new_n299), .b(new_n279), .c(new_n282), .o1(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n297), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n298), .b(new_n301), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n12x5               g208(.a(new_n284), .b(new_n276), .c(new_n297), .out0(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n287), .c(new_n179), .d(new_n278), .o1(new_n305));
  oao003aa1n02x5               g210(.a(\a[29] ), .b(\b[28] ), .c(new_n296), .carry(new_n306));
  xnrc02aa1n02x5               g211(.a(\b[29] ), .b(\a[30] ), .out0(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n307), .b(new_n305), .c(new_n306), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n304), .o1(new_n309));
  aoi012aa1n02x7               g214(.a(new_n309), .b(new_n279), .c(new_n282), .o1(new_n310));
  nano22aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n307), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n308), .b(new_n311), .o1(\s[30] ));
  norb02aa1n06x5               g217(.a(new_n304), .b(new_n307), .out0(new_n313));
  inv000aa1n02x5               g218(.a(new_n313), .o1(new_n314));
  aoi012aa1n02x7               g219(.a(new_n314), .b(new_n279), .c(new_n282), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .c(new_n306), .carry(new_n316));
  xnrc02aa1n02x5               g221(.a(\b[30] ), .b(\a[31] ), .out0(new_n317));
  nano22aa1n03x5               g222(.a(new_n315), .b(new_n316), .c(new_n317), .out0(new_n318));
  aoai13aa1n03x5               g223(.a(new_n313), .b(new_n287), .c(new_n179), .d(new_n278), .o1(new_n319));
  tech160nm_fiaoi012aa1n02p5x5 g224(.a(new_n317), .b(new_n319), .c(new_n316), .o1(new_n320));
  norp02aa1n03x5               g225(.a(new_n320), .b(new_n318), .o1(\s[31] ));
  xnrb03aa1n02x5               g226(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g227(.a(\a[3] ), .b(\b[2] ), .c(new_n101), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g229(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g230(.a(new_n119), .b(new_n112), .out0(new_n326));
  oai112aa1n02x5               g231(.a(new_n107), .b(new_n326), .c(new_n106), .d(new_n101), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[6] ), .b(\b[5] ), .out0(new_n328));
  xobna2aa1n03x5               g233(.a(new_n328), .b(new_n327), .c(new_n119), .out0(\s[6] ));
  nanb02aa1n02x5               g234(.a(new_n114), .b(new_n115), .out0(new_n330));
  nanp03aa1n02x5               g235(.a(new_n327), .b(new_n119), .c(new_n328), .o1(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n330), .b(new_n331), .c(\a[6] ), .d(\b[5] ), .o1(new_n332));
  oai112aa1n02x5               g237(.a(new_n331), .b(new_n330), .c(\b[5] ), .d(\a[6] ), .o1(new_n333));
  norb02aa1n02x5               g238(.a(new_n333), .b(new_n332), .out0(\s[7] ));
  norp02aa1n02x5               g239(.a(new_n332), .b(new_n114), .o1(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g241(.a(new_n187), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


