// Benchmark "adder" written by ABC on Thu Jul 18 07:50:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n276, new_n277, new_n278, new_n279, new_n280, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n334, new_n337, new_n338, new_n340, new_n342;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[1] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[0] ), .o1(new_n98));
  norp02aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n03x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oaoi13aa1n09x5               g005(.a(new_n99), .b(new_n100), .c(new_n97), .d(new_n98), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor002aa1d32x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norp02aa1n06x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n102), .b(new_n105), .c(new_n104), .d(new_n103), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\a[3] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[2] ), .o1(new_n108));
  aoai13aa1n04x5               g013(.a(new_n102), .b(new_n103), .c(new_n108), .d(new_n107), .o1(new_n109));
  oai012aa1n12x5               g014(.a(new_n109), .b(new_n106), .c(new_n101), .o1(new_n110));
  tech160nm_fixorc02aa1n02p5x5 g015(.a(\a[6] ), .b(\b[5] ), .out0(new_n111));
  tech160nm_fixorc02aa1n02p5x5 g016(.a(\a[5] ), .b(\b[4] ), .out0(new_n112));
  nor022aa1n08x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1d04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nanp02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nor002aa1n16x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n06x5               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  nano22aa1n03x7               g022(.a(new_n117), .b(new_n111), .c(new_n112), .out0(new_n118));
  inv000aa1d42x5               g023(.a(\a[6] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[5] ), .o1(new_n120));
  nor002aa1n03x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  tech160nm_fioaoi03aa1n03p5x5 g026(.a(new_n119), .b(new_n120), .c(new_n121), .o1(new_n122));
  ao0012aa1n03x7               g027(.a(new_n113), .b(new_n116), .c(new_n114), .o(new_n123));
  oabi12aa1n06x5               g028(.a(new_n123), .b(new_n117), .c(new_n122), .out0(new_n124));
  nor002aa1n12x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nand02aa1n10x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n124), .c(new_n118), .d(new_n110), .o1(new_n128));
  tech160nm_fioai012aa1n03p5x5 g033(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .o1(new_n129));
  xorb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1d24x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nand42aa1d28x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  and002aa1n03x5               g038(.a(\b[0] ), .b(\a[1] ), .o(new_n134));
  oaoi03aa1n02x5               g039(.a(\a[2] ), .b(\b[1] ), .c(new_n134), .o1(new_n135));
  norb02aa1n03x5               g040(.a(new_n102), .b(new_n103), .out0(new_n136));
  norb02aa1n02x5               g041(.a(new_n105), .b(new_n104), .out0(new_n137));
  nanp03aa1n02x5               g042(.a(new_n135), .b(new_n136), .c(new_n137), .o1(new_n138));
  nano23aa1n03x7               g043(.a(new_n116), .b(new_n113), .c(new_n114), .d(new_n115), .out0(new_n139));
  nanp03aa1n02x5               g044(.a(new_n139), .b(new_n111), .c(new_n112), .o1(new_n140));
  oao003aa1n02x5               g045(.a(new_n119), .b(new_n120), .c(new_n121), .carry(new_n141));
  tech160nm_fiaoi012aa1n04x5   g046(.a(new_n123), .b(new_n139), .c(new_n141), .o1(new_n142));
  aoai13aa1n04x5               g047(.a(new_n142), .b(new_n140), .c(new_n138), .d(new_n109), .o1(new_n143));
  aoai13aa1n03x5               g048(.a(new_n133), .b(new_n125), .c(new_n143), .d(new_n127), .o1(new_n144));
  nand42aa1n16x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  nor002aa1d32x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  nanb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n144), .c(new_n132), .out0(\s[11] ));
  aoai13aa1n02x5               g054(.a(new_n148), .b(new_n131), .c(new_n129), .d(new_n133), .o1(new_n150));
  nor002aa1d32x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nand42aa1d28x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  aoib12aa1n06x5               g058(.a(new_n146), .b(new_n152), .c(new_n151), .out0(new_n154));
  inv020aa1n03x5               g059(.a(new_n146), .o1(new_n155));
  aoai13aa1n02x5               g060(.a(new_n155), .b(new_n147), .c(new_n144), .d(new_n132), .o1(new_n156));
  aoi022aa1n02x5               g061(.a(new_n156), .b(new_n153), .c(new_n150), .d(new_n154), .o1(\s[12] ));
  oaib12aa1n09x5               g062(.a(new_n155), .b(new_n151), .c(new_n152), .out0(new_n158));
  norb03aa1n09x5               g063(.a(new_n126), .b(new_n131), .c(new_n125), .out0(new_n159));
  nano22aa1n09x5               g064(.a(new_n146), .b(new_n133), .c(new_n145), .out0(new_n160));
  nand23aa1n09x5               g065(.a(new_n158), .b(new_n160), .c(new_n159), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n06x5               g067(.a(new_n162), .b(new_n124), .c(new_n118), .d(new_n110), .o1(new_n163));
  nanb03aa1n12x5               g068(.a(new_n146), .b(new_n133), .c(new_n145), .out0(new_n164));
  norb03aa1n09x5               g069(.a(new_n133), .b(new_n131), .c(new_n125), .out0(new_n165));
  tech160nm_fiaoi012aa1n03p5x5 g070(.a(new_n151), .b(new_n146), .c(new_n152), .o1(new_n166));
  oai013aa1d12x5               g071(.a(new_n166), .b(new_n154), .c(new_n165), .d(new_n164), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  and002aa1n02x5               g073(.a(\b[12] ), .b(\a[13] ), .o(new_n169));
  nor002aa1d32x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  nor042aa1n04x5               g075(.a(new_n169), .b(new_n170), .o1(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n163), .c(new_n168), .out0(\s[13] ));
  inv000aa1d42x5               g077(.a(new_n170), .o1(new_n173));
  aoai13aa1n02x5               g078(.a(new_n171), .b(new_n167), .c(new_n143), .d(new_n162), .o1(new_n174));
  xorc02aa1n12x5               g079(.a(\a[14] ), .b(\b[13] ), .out0(new_n175));
  xnbna2aa1n03x5               g080(.a(new_n175), .b(new_n174), .c(new_n173), .out0(\s[14] ));
  nanp02aa1n02x5               g081(.a(new_n175), .b(new_n171), .o1(new_n177));
  norp02aa1n02x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  aoi012aa1n02x5               g084(.a(new_n178), .b(new_n170), .c(new_n179), .o1(new_n180));
  aoai13aa1n06x5               g085(.a(new_n180), .b(new_n177), .c(new_n163), .d(new_n168), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  nanp02aa1n09x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norb02aa1n02x5               g089(.a(new_n184), .b(new_n183), .out0(new_n185));
  nor042aa1n04x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  nanp02aa1n09x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nanb02aa1n02x5               g092(.a(new_n186), .b(new_n187), .out0(new_n188));
  aoai13aa1n02x5               g093(.a(new_n188), .b(new_n183), .c(new_n181), .d(new_n185), .o1(new_n189));
  nanp02aa1n02x5               g094(.a(new_n181), .b(new_n185), .o1(new_n190));
  nona22aa1n02x4               g095(.a(new_n190), .b(new_n188), .c(new_n183), .out0(new_n191));
  nanp02aa1n03x5               g096(.a(new_n191), .b(new_n189), .o1(\s[16] ));
  nano23aa1n06x5               g097(.a(new_n186), .b(new_n183), .c(new_n187), .d(new_n184), .out0(new_n193));
  nano32aa1d12x5               g098(.a(new_n161), .b(new_n193), .c(new_n171), .d(new_n175), .out0(new_n194));
  aoai13aa1n12x5               g099(.a(new_n194), .b(new_n124), .c(new_n118), .d(new_n110), .o1(new_n195));
  nand03aa1n02x5               g100(.a(new_n193), .b(new_n171), .c(new_n175), .o1(new_n196));
  inv000aa1n03x5               g101(.a(new_n196), .o1(new_n197));
  oa0012aa1n02x5               g102(.a(new_n187), .b(new_n186), .c(new_n183), .o(new_n198));
  aoib12aa1n06x5               g103(.a(new_n198), .b(new_n193), .c(new_n180), .out0(new_n199));
  aobi12aa1d24x5               g104(.a(new_n199), .b(new_n197), .c(new_n167), .out0(new_n200));
  xorc02aa1n02x5               g105(.a(\a[17] ), .b(\b[16] ), .out0(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n195), .c(new_n200), .out0(\s[17] ));
  inv040aa1d32x5               g107(.a(\a[18] ), .o1(new_n203));
  inv040aa1d30x5               g108(.a(\a[17] ), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\b[16] ), .o1(new_n205));
  nanp02aa1n09x5               g110(.a(new_n195), .b(new_n200), .o1(new_n206));
  oaoi03aa1n03x5               g111(.a(new_n204), .b(new_n205), .c(new_n206), .o1(new_n207));
  xorb03aa1n02x5               g112(.a(new_n207), .b(\b[17] ), .c(new_n203), .out0(\s[18] ));
  xroi22aa1d06x4               g113(.a(new_n204), .b(\b[16] ), .c(new_n203), .d(\b[17] ), .out0(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor042aa1n02x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  aoi112aa1n09x5               g116(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n212));
  norp02aa1n02x5               g117(.a(new_n212), .b(new_n211), .o1(new_n213));
  aoai13aa1n06x5               g118(.a(new_n213), .b(new_n210), .c(new_n195), .d(new_n200), .o1(new_n214));
  xorb03aa1n02x5               g119(.a(new_n214), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n04x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nor042aa1n04x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nor042aa1n06x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand42aa1n16x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  norb02aa1d21x5               g125(.a(new_n220), .b(new_n219), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n222), .b(new_n218), .c(new_n214), .d(new_n217), .o1(new_n223));
  norb02aa1n03x5               g128(.a(new_n217), .b(new_n218), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n214), .b(new_n224), .o1(new_n225));
  nona22aa1n02x5               g130(.a(new_n225), .b(new_n222), .c(new_n218), .out0(new_n226));
  nanp02aa1n03x5               g131(.a(new_n226), .b(new_n223), .o1(\s[20] ));
  nano23aa1n06x5               g132(.a(new_n219), .b(new_n218), .c(new_n220), .d(new_n217), .out0(new_n228));
  nand02aa1d04x5               g133(.a(new_n209), .b(new_n228), .o1(new_n229));
  oai112aa1n06x5               g134(.a(new_n224), .b(new_n221), .c(new_n212), .d(new_n211), .o1(new_n230));
  oai012aa1n06x5               g135(.a(new_n220), .b(new_n219), .c(new_n218), .o1(new_n231));
  nand02aa1d06x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n229), .c(new_n195), .d(new_n200), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  tech160nm_fixorc02aa1n04x5   g141(.a(\a[21] ), .b(\b[20] ), .out0(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[21] ), .b(\a[22] ), .out0(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n236), .c(new_n234), .d(new_n237), .o1(new_n239));
  nand02aa1n02x5               g144(.a(new_n234), .b(new_n237), .o1(new_n240));
  nona22aa1n02x5               g145(.a(new_n240), .b(new_n238), .c(new_n236), .out0(new_n241));
  nand42aa1n02x5               g146(.a(new_n241), .b(new_n239), .o1(\s[22] ));
  norb02aa1n03x5               g147(.a(new_n237), .b(new_n238), .out0(new_n243));
  nanp03aa1n02x5               g148(.a(new_n243), .b(new_n209), .c(new_n228), .o1(new_n244));
  orn002aa1n02x5               g149(.a(\a[21] ), .b(\b[20] ), .o(new_n245));
  oaoi03aa1n09x5               g150(.a(\a[22] ), .b(\b[21] ), .c(new_n245), .o1(new_n246));
  tech160nm_fiaoi012aa1n02p5x5 g151(.a(new_n246), .b(new_n232), .c(new_n243), .o1(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n244), .c(new_n195), .d(new_n200), .o1(new_n248));
  xorb03aa1n02x5               g153(.a(new_n248), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g154(.a(\b[22] ), .b(\a[23] ), .o1(new_n250));
  nand42aa1n02x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  norb02aa1n02x5               g156(.a(new_n251), .b(new_n250), .out0(new_n252));
  nor042aa1n03x5               g157(.a(\b[23] ), .b(\a[24] ), .o1(new_n253));
  nand42aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n03x5               g161(.a(new_n256), .b(new_n250), .c(new_n248), .d(new_n252), .o1(new_n257));
  nand02aa1n02x5               g162(.a(new_n248), .b(new_n252), .o1(new_n258));
  nona22aa1n02x5               g163(.a(new_n258), .b(new_n256), .c(new_n250), .out0(new_n259));
  nanp02aa1n03x5               g164(.a(new_n259), .b(new_n257), .o1(\s[24] ));
  xorc02aa1n02x5               g165(.a(\a[22] ), .b(\b[21] ), .out0(new_n261));
  nanp02aa1n02x5               g166(.a(new_n261), .b(new_n237), .o1(new_n262));
  nano23aa1n09x5               g167(.a(new_n250), .b(new_n253), .c(new_n254), .d(new_n251), .out0(new_n263));
  inv000aa1n02x5               g168(.a(new_n263), .o1(new_n264));
  nona32aa1n02x4               g169(.a(new_n206), .b(new_n264), .c(new_n262), .d(new_n229), .out0(new_n265));
  nanb03aa1n03x5               g170(.a(new_n229), .b(new_n263), .c(new_n243), .out0(new_n266));
  aoi112aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n267));
  nanp02aa1n06x5               g172(.a(new_n263), .b(new_n246), .o1(new_n268));
  nona22aa1d18x5               g173(.a(new_n268), .b(new_n267), .c(new_n253), .out0(new_n269));
  aoi013aa1n03x5               g174(.a(new_n269), .b(new_n232), .c(new_n243), .d(new_n263), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n270), .b(new_n266), .c(new_n195), .d(new_n200), .o1(new_n271));
  xorc02aa1n12x5               g176(.a(\a[25] ), .b(\b[24] ), .out0(new_n272));
  aoi112aa1n03x5               g177(.a(new_n264), .b(new_n262), .c(new_n230), .d(new_n231), .o1(new_n273));
  norp03aa1n02x5               g178(.a(new_n273), .b(new_n272), .c(new_n269), .o1(new_n274));
  aoi022aa1n02x5               g179(.a(new_n274), .b(new_n265), .c(new_n271), .d(new_n272), .o1(\s[25] ));
  nor002aa1n02x5               g180(.a(\b[24] ), .b(\a[25] ), .o1(new_n276));
  xnrc02aa1n12x5               g181(.a(\b[25] ), .b(\a[26] ), .out0(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n276), .c(new_n271), .d(new_n272), .o1(new_n278));
  nand02aa1n02x5               g183(.a(new_n271), .b(new_n272), .o1(new_n279));
  nona22aa1n02x5               g184(.a(new_n279), .b(new_n277), .c(new_n276), .out0(new_n280));
  nanp02aa1n03x5               g185(.a(new_n280), .b(new_n278), .o1(\s[26] ));
  nanb03aa1n02x5               g186(.a(new_n165), .b(new_n158), .c(new_n160), .out0(new_n282));
  aoai13aa1n02x5               g187(.a(new_n199), .b(new_n196), .c(new_n282), .d(new_n166), .o1(new_n283));
  norb02aa1n06x5               g188(.a(new_n272), .b(new_n277), .out0(new_n284));
  nano32aa1d12x5               g189(.a(new_n229), .b(new_n284), .c(new_n243), .d(new_n263), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n283), .c(new_n143), .d(new_n194), .o1(new_n286));
  inv000aa1d42x5               g191(.a(\a[26] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(\b[25] ), .o1(new_n288));
  oao003aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n276), .carry(new_n289));
  oaoi13aa1n09x5               g194(.a(new_n289), .b(new_n284), .c(new_n273), .d(new_n269), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnbna2aa1n03x5               g196(.a(new_n291), .b(new_n286), .c(new_n290), .out0(\s[27] ));
  xnrc02aa1n02x5               g197(.a(\b[27] ), .b(\a[28] ), .out0(new_n293));
  nor042aa1n03x5               g198(.a(\b[26] ), .b(\a[27] ), .o1(new_n294));
  inv000aa1n03x5               g199(.a(new_n294), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n291), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n295), .b(new_n296), .c(new_n286), .d(new_n290), .o1(new_n297));
  nand02aa1n02x5               g202(.a(new_n297), .b(new_n293), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n269), .o1(new_n299));
  nona22aa1n09x5               g204(.a(new_n232), .b(new_n264), .c(new_n262), .out0(new_n300));
  inv000aa1d42x5               g205(.a(new_n284), .o1(new_n301));
  inv000aa1n02x5               g206(.a(new_n289), .o1(new_n302));
  aoai13aa1n12x5               g207(.a(new_n302), .b(new_n301), .c(new_n299), .d(new_n300), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n291), .b(new_n303), .c(new_n206), .d(new_n285), .o1(new_n304));
  nona22aa1n02x5               g209(.a(new_n304), .b(new_n293), .c(new_n294), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n298), .b(new_n305), .o1(\s[28] ));
  norb02aa1n09x5               g211(.a(new_n291), .b(new_n293), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n206), .d(new_n285), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n307), .o1(new_n309));
  oao003aa1n03x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n310));
  aoai13aa1n02x7               g215(.a(new_n310), .b(new_n309), .c(new_n286), .d(new_n290), .o1(new_n311));
  tech160nm_fixorc02aa1n03p5x5 g216(.a(\a[29] ), .b(\b[28] ), .out0(new_n312));
  norb02aa1n02x5               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n308), .d(new_n313), .o1(\s[29] ));
  xnrb03aa1n02x5               g219(.a(new_n134), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g220(.a(new_n293), .b(new_n291), .c(new_n312), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n303), .c(new_n206), .d(new_n285), .o1(new_n317));
  inv000aa1n02x5               g222(.a(new_n316), .o1(new_n318));
  oaoi03aa1n02x5               g223(.a(\a[29] ), .b(\b[28] ), .c(new_n310), .o1(new_n319));
  inv000aa1n03x5               g224(.a(new_n319), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n318), .c(new_n286), .d(new_n290), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  norp02aa1n02x5               g227(.a(new_n319), .b(new_n322), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n317), .d(new_n323), .o1(\s[30] ));
  nano22aa1d33x5               g229(.a(new_n309), .b(new_n312), .c(new_n322), .out0(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n303), .c(new_n206), .d(new_n285), .o1(new_n326));
  xorc02aa1n02x5               g231(.a(\a[31] ), .b(\b[30] ), .out0(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n320), .carry(new_n328));
  norb02aa1n02x5               g233(.a(new_n328), .b(new_n327), .out0(new_n329));
  inv000aa1d42x5               g234(.a(new_n325), .o1(new_n330));
  aoai13aa1n02x7               g235(.a(new_n328), .b(new_n330), .c(new_n286), .d(new_n290), .o1(new_n331));
  aoi022aa1n03x5               g236(.a(new_n331), .b(new_n327), .c(new_n326), .d(new_n329), .o1(\s[31] ));
  xorb03aa1n02x5               g237(.a(new_n101), .b(\b[2] ), .c(new_n107), .out0(\s[3] ));
  aoi112aa1n02x5               g238(.a(new_n104), .b(new_n136), .c(new_n135), .d(new_n105), .o1(new_n334));
  aoib12aa1n02x5               g239(.a(new_n334), .b(new_n110), .c(new_n103), .out0(\s[4] ));
  xorb03aa1n02x5               g240(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n03x5               g241(.a(new_n111), .b(new_n121), .c(new_n110), .d(new_n112), .o1(new_n337));
  aoi112aa1n02x5               g242(.a(new_n121), .b(new_n111), .c(new_n110), .d(new_n112), .o1(new_n338));
  norb02aa1n02x5               g243(.a(new_n337), .b(new_n338), .out0(\s[6] ));
  nanp02aa1n03x5               g244(.a(new_n337), .b(new_n122), .o1(new_n340));
  xorb03aa1n02x5               g245(.a(new_n340), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g246(.a(new_n116), .b(new_n340), .c(new_n115), .o1(new_n342));
  xnrb03aa1n03x5               g247(.a(new_n342), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g248(.a(new_n143), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


