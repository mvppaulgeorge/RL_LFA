// Benchmark "adder" written by ABC on Thu Jul 18 02:59:40 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n176, new_n177, new_n178, new_n179, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n293, new_n296, new_n298, new_n299,
    new_n301;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nand42aa1n04x5               g001(.a(\b[3] ), .b(\a[4] ), .o1(new_n97));
  nor022aa1n16x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  nor002aa1n12x5               g003(.a(\b[2] ), .b(\a[3] ), .o1(new_n99));
  oa0012aa1n03x5               g004(.a(new_n97), .b(new_n98), .c(new_n99), .o(new_n100));
  inv000aa1d42x5               g005(.a(\a[2] ), .o1(new_n101));
  inv030aa1d32x5               g006(.a(\b[1] ), .o1(new_n102));
  nand42aa1n08x5               g007(.a(\b[0] ), .b(\a[1] ), .o1(new_n103));
  tech160nm_fioaoi03aa1n03p5x5 g008(.a(new_n101), .b(new_n102), .c(new_n103), .o1(new_n104));
  nand42aa1n03x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n09x5               g010(.a(new_n97), .b(new_n105), .c(new_n99), .d(new_n98), .out0(new_n106));
  oabi12aa1n12x5               g011(.a(new_n100), .b(new_n104), .c(new_n106), .out0(new_n107));
  tech160nm_fixnrc02aa1n02p5x5 g012(.a(\b[5] ), .b(\a[6] ), .out0(new_n108));
  xnrc02aa1n02x5               g013(.a(\b[4] ), .b(\a[5] ), .out0(new_n109));
  nand42aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor022aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  norp02aa1n04x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n09x5               g018(.a(new_n112), .b(new_n110), .c(new_n113), .d(new_n111), .out0(new_n114));
  nor043aa1n03x5               g019(.a(new_n114), .b(new_n109), .c(new_n108), .o1(new_n115));
  orn002aa1n03x5               g020(.a(\a[5] ), .b(\b[4] ), .o(new_n116));
  tech160nm_fioaoi03aa1n02p5x5 g021(.a(\a[6] ), .b(\b[5] ), .c(new_n116), .o1(new_n117));
  oai012aa1n02x5               g022(.a(new_n112), .b(new_n113), .c(new_n111), .o1(new_n118));
  oaib12aa1n06x5               g023(.a(new_n118), .b(new_n114), .c(new_n117), .out0(new_n119));
  aoi012aa1n02x5               g024(.a(new_n119), .b(new_n107), .c(new_n115), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[9] ), .b(\b[8] ), .c(new_n120), .o1(new_n121));
  xorb03aa1n02x5               g026(.a(new_n121), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  norp02aa1n06x5               g027(.a(\b[10] ), .b(\a[11] ), .o1(new_n123));
  nand42aa1n03x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  inv040aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  nor002aa1n06x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nor002aa1n06x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1n20x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  tech160nm_fioai012aa1n04x5   g034(.a(new_n129), .b(new_n128), .c(new_n127), .o1(new_n130));
  nand42aa1d28x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nano23aa1d15x5               g036(.a(new_n127), .b(new_n128), .c(new_n129), .d(new_n131), .out0(new_n132));
  inv000aa1d42x5               g037(.a(new_n132), .o1(new_n133));
  oaoi13aa1n03x5               g038(.a(new_n126), .b(new_n130), .c(new_n120), .d(new_n133), .o1(new_n134));
  oai112aa1n02x5               g039(.a(new_n130), .b(new_n126), .c(new_n120), .d(new_n133), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(\s[11] ));
  norp02aa1n03x5               g041(.a(new_n134), .b(new_n123), .o1(new_n137));
  nor002aa1d32x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n138), .o1(new_n139));
  tech160nm_finand02aa1n03p5x5 g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n137), .b(new_n140), .c(new_n139), .out0(\s[12] ));
  nona23aa1n09x5               g046(.a(new_n140), .b(new_n124), .c(new_n123), .d(new_n138), .out0(new_n142));
  norb02aa1n02x5               g047(.a(new_n132), .b(new_n142), .out0(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n119), .c(new_n107), .d(new_n115), .o1(new_n144));
  nanp02aa1n02x5               g049(.a(new_n123), .b(new_n140), .o1(new_n145));
  oai112aa1n06x5               g050(.a(new_n145), .b(new_n139), .c(new_n142), .d(new_n130), .o1(new_n146));
  nanb02aa1n03x5               g051(.a(new_n146), .b(new_n144), .out0(new_n147));
  xorb03aa1n02x5               g052(.a(new_n147), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nand42aa1n03x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  aoi012aa1n02x5               g055(.a(new_n149), .b(new_n147), .c(new_n150), .o1(new_n151));
  xnrb03aa1n02x5               g056(.a(new_n151), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n12x5               g057(.a(\b[13] ), .b(\a[14] ), .o1(new_n153));
  nand42aa1n04x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nano23aa1n06x5               g059(.a(new_n149), .b(new_n153), .c(new_n154), .d(new_n150), .out0(new_n155));
  oaih12aa1n06x5               g060(.a(new_n154), .b(new_n153), .c(new_n149), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  xorc02aa1n12x5               g062(.a(\a[15] ), .b(\b[14] ), .out0(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n157), .c(new_n147), .d(new_n155), .o1(new_n159));
  aoi112aa1n02x5               g064(.a(new_n158), .b(new_n157), .c(new_n147), .d(new_n155), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(\s[15] ));
  xnrc02aa1n02x5               g066(.a(\b[15] ), .b(\a[16] ), .out0(new_n162));
  oai112aa1n02x5               g067(.a(new_n159), .b(new_n162), .c(\b[14] ), .d(\a[15] ), .o1(new_n163));
  oaoi13aa1n06x5               g068(.a(new_n162), .b(new_n159), .c(\a[15] ), .d(\b[14] ), .o1(new_n164));
  norb02aa1n02x7               g069(.a(new_n163), .b(new_n164), .out0(\s[16] ));
  xorc02aa1n03x5               g070(.a(\a[16] ), .b(\b[15] ), .out0(new_n166));
  nand22aa1n03x5               g071(.a(new_n166), .b(new_n158), .o1(new_n167));
  nano23aa1n06x5               g072(.a(new_n167), .b(new_n142), .c(new_n132), .d(new_n155), .out0(new_n168));
  aoai13aa1n06x5               g073(.a(new_n168), .b(new_n119), .c(new_n107), .d(new_n115), .o1(new_n169));
  norb02aa1n02x7               g074(.a(new_n155), .b(new_n167), .out0(new_n170));
  aoi112aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n171));
  oai022aa1n03x5               g076(.a(new_n167), .b(new_n156), .c(\b[15] ), .d(\a[16] ), .o1(new_n172));
  aoi112aa1n09x5               g077(.a(new_n172), .b(new_n171), .c(new_n146), .d(new_n170), .o1(new_n173));
  nanp02aa1n12x5               g078(.a(new_n173), .b(new_n169), .o1(new_n174));
  xorb03aa1n02x5               g079(.a(new_n174), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g080(.a(\a[18] ), .o1(new_n176));
  inv000aa1d42x5               g081(.a(\a[17] ), .o1(new_n177));
  inv000aa1d42x5               g082(.a(\b[16] ), .o1(new_n178));
  oaoi03aa1n02x5               g083(.a(new_n177), .b(new_n178), .c(new_n174), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[17] ), .c(new_n176), .out0(\s[18] ));
  xroi22aa1d04x5               g085(.a(new_n177), .b(\b[16] ), .c(new_n176), .d(\b[17] ), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n178), .b(new_n177), .o1(new_n182));
  oaoi03aa1n02x5               g087(.a(\a[18] ), .b(\b[17] ), .c(new_n182), .o1(new_n183));
  nor022aa1n08x5               g088(.a(\b[18] ), .b(\a[19] ), .o1(new_n184));
  nand42aa1d28x5               g089(.a(\b[18] ), .b(\a[19] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n183), .c(new_n174), .d(new_n181), .o1(new_n187));
  aoi112aa1n02x5               g092(.a(new_n186), .b(new_n183), .c(new_n174), .d(new_n181), .o1(new_n188));
  norb02aa1n02x5               g093(.a(new_n187), .b(new_n188), .out0(\s[19] ));
  xnrc02aa1n02x5               g094(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n04x5               g095(.a(\b[19] ), .b(\a[20] ), .o1(new_n191));
  nand42aa1n10x5               g096(.a(\b[19] ), .b(\a[20] ), .o1(new_n192));
  norb02aa1n02x5               g097(.a(new_n192), .b(new_n191), .out0(new_n193));
  nona22aa1n03x5               g098(.a(new_n187), .b(new_n193), .c(new_n184), .out0(new_n194));
  orn002aa1n06x5               g099(.a(\a[19] ), .b(\b[18] ), .o(new_n195));
  aobi12aa1n03x5               g100(.a(new_n193), .b(new_n187), .c(new_n195), .out0(new_n196));
  norb02aa1n03x4               g101(.a(new_n194), .b(new_n196), .out0(\s[20] ));
  nano23aa1n03x5               g102(.a(new_n184), .b(new_n191), .c(new_n192), .d(new_n185), .out0(new_n198));
  nanp02aa1n02x5               g103(.a(new_n181), .b(new_n198), .o1(new_n199));
  oai022aa1n02x5               g104(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n200));
  oaib12aa1n02x5               g105(.a(new_n200), .b(new_n176), .c(\b[17] ), .out0(new_n201));
  nona23aa1n12x5               g106(.a(new_n192), .b(new_n185), .c(new_n184), .d(new_n191), .out0(new_n202));
  oaoi03aa1n02x5               g107(.a(\a[20] ), .b(\b[19] ), .c(new_n195), .o1(new_n203));
  oabi12aa1n12x5               g108(.a(new_n203), .b(new_n202), .c(new_n201), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  aoai13aa1n03x5               g110(.a(new_n205), .b(new_n199), .c(new_n173), .d(new_n169), .o1(new_n206));
  xorb03aa1n02x5               g111(.a(new_n206), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g112(.a(\b[20] ), .b(\a[21] ), .o1(new_n208));
  xorc02aa1n02x5               g113(.a(\a[21] ), .b(\b[20] ), .out0(new_n209));
  xorc02aa1n02x5               g114(.a(\a[22] ), .b(\b[21] ), .out0(new_n210));
  aoi112aa1n02x7               g115(.a(new_n208), .b(new_n210), .c(new_n206), .d(new_n209), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n210), .b(new_n208), .c(new_n206), .d(new_n209), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(\s[22] ));
  inv000aa1d42x5               g118(.a(\a[21] ), .o1(new_n214));
  inv000aa1d42x5               g119(.a(\a[22] ), .o1(new_n215));
  xroi22aa1d04x5               g120(.a(new_n214), .b(\b[20] ), .c(new_n215), .d(\b[21] ), .out0(new_n216));
  nanp03aa1n03x5               g121(.a(new_n216), .b(new_n181), .c(new_n198), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[21] ), .o1(new_n218));
  oaoi03aa1n09x5               g123(.a(new_n215), .b(new_n218), .c(new_n208), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  aoi012aa1n02x5               g125(.a(new_n220), .b(new_n204), .c(new_n216), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n217), .c(new_n173), .d(new_n169), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g128(.a(\b[22] ), .b(\a[23] ), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[23] ), .b(\b[22] ), .out0(new_n225));
  xorc02aa1n02x5               g130(.a(\a[24] ), .b(\b[23] ), .out0(new_n226));
  aoi112aa1n02x5               g131(.a(new_n224), .b(new_n226), .c(new_n222), .d(new_n225), .o1(new_n227));
  aoai13aa1n03x5               g132(.a(new_n226), .b(new_n224), .c(new_n222), .d(new_n225), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(\s[24] ));
  and002aa1n02x5               g134(.a(new_n226), .b(new_n225), .o(new_n230));
  inv000aa1n02x5               g135(.a(new_n230), .o1(new_n231));
  nano32aa1n02x4               g136(.a(new_n231), .b(new_n216), .c(new_n181), .d(new_n198), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n216), .b(new_n203), .c(new_n198), .d(new_n183), .o1(new_n233));
  aoi112aa1n02x5               g138(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n234));
  oab012aa1n02x4               g139(.a(new_n234), .b(\a[24] ), .c(\b[23] ), .out0(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n231), .c(new_n233), .d(new_n219), .o1(new_n236));
  tech160nm_fixorc02aa1n04x5   g141(.a(\a[25] ), .b(\b[24] ), .out0(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n236), .c(new_n174), .d(new_n232), .o1(new_n238));
  aoi112aa1n02x5               g143(.a(new_n237), .b(new_n236), .c(new_n174), .d(new_n232), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n238), .b(new_n239), .out0(\s[25] ));
  nor042aa1n03x5               g145(.a(\b[24] ), .b(\a[25] ), .o1(new_n241));
  tech160nm_fixorc02aa1n04x5   g146(.a(\a[26] ), .b(\b[25] ), .out0(new_n242));
  nona22aa1n03x5               g147(.a(new_n238), .b(new_n242), .c(new_n241), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n241), .o1(new_n244));
  aobi12aa1n03x5               g149(.a(new_n242), .b(new_n238), .c(new_n244), .out0(new_n245));
  norb02aa1n03x4               g150(.a(new_n243), .b(new_n245), .out0(\s[26] ));
  and002aa1n06x5               g151(.a(new_n242), .b(new_n237), .o(new_n247));
  nano22aa1n03x7               g152(.a(new_n217), .b(new_n230), .c(new_n247), .out0(new_n248));
  nanp02aa1n09x5               g153(.a(new_n174), .b(new_n248), .o1(new_n249));
  oao003aa1n02x5               g154(.a(\a[26] ), .b(\b[25] ), .c(new_n244), .carry(new_n250));
  aobi12aa1n12x5               g155(.a(new_n250), .b(new_n236), .c(new_n247), .out0(new_n251));
  xorc02aa1n02x5               g156(.a(\a[27] ), .b(\b[26] ), .out0(new_n252));
  xnbna2aa1n06x5               g157(.a(new_n252), .b(new_n249), .c(new_n251), .out0(\s[27] ));
  norp02aa1n02x5               g158(.a(\b[26] ), .b(\a[27] ), .o1(new_n254));
  inv040aa1n03x5               g159(.a(new_n254), .o1(new_n255));
  aobi12aa1n06x5               g160(.a(new_n252), .b(new_n249), .c(new_n251), .out0(new_n256));
  xnrc02aa1n02x5               g161(.a(\b[27] ), .b(\a[28] ), .out0(new_n257));
  nano22aa1n03x5               g162(.a(new_n256), .b(new_n255), .c(new_n257), .out0(new_n258));
  inv020aa1n03x5               g163(.a(new_n248), .o1(new_n259));
  aoi012aa1n06x5               g164(.a(new_n259), .b(new_n173), .c(new_n169), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n230), .b(new_n220), .c(new_n204), .d(new_n216), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n247), .o1(new_n262));
  aoai13aa1n06x5               g167(.a(new_n250), .b(new_n262), .c(new_n261), .d(new_n235), .o1(new_n263));
  oaih12aa1n02x5               g168(.a(new_n252), .b(new_n263), .c(new_n260), .o1(new_n264));
  aoi012aa1n03x5               g169(.a(new_n257), .b(new_n264), .c(new_n255), .o1(new_n265));
  norp02aa1n03x5               g170(.a(new_n265), .b(new_n258), .o1(\s[28] ));
  xnrc02aa1n02x5               g171(.a(\b[28] ), .b(\a[29] ), .out0(new_n267));
  norb02aa1n02x5               g172(.a(new_n252), .b(new_n257), .out0(new_n268));
  aobi12aa1n06x5               g173(.a(new_n268), .b(new_n249), .c(new_n251), .out0(new_n269));
  oao003aa1n02x5               g174(.a(\a[28] ), .b(\b[27] ), .c(new_n255), .carry(new_n270));
  nano22aa1n03x7               g175(.a(new_n269), .b(new_n267), .c(new_n270), .out0(new_n271));
  oaih12aa1n02x5               g176(.a(new_n268), .b(new_n263), .c(new_n260), .o1(new_n272));
  aoi012aa1n02x5               g177(.a(new_n267), .b(new_n272), .c(new_n270), .o1(new_n273));
  norp02aa1n03x5               g178(.a(new_n273), .b(new_n271), .o1(\s[29] ));
  xorb03aa1n02x5               g179(.a(new_n103), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g180(.a(new_n252), .b(new_n267), .c(new_n257), .out0(new_n276));
  oaih12aa1n02x5               g181(.a(new_n276), .b(new_n263), .c(new_n260), .o1(new_n277));
  oao003aa1n02x5               g182(.a(\a[29] ), .b(\b[28] ), .c(new_n270), .carry(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[29] ), .b(\a[30] ), .out0(new_n279));
  aoi012aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n278), .o1(new_n280));
  aobi12aa1n06x5               g185(.a(new_n276), .b(new_n249), .c(new_n251), .out0(new_n281));
  nano22aa1n03x7               g186(.a(new_n281), .b(new_n278), .c(new_n279), .out0(new_n282));
  norp02aa1n03x5               g187(.a(new_n280), .b(new_n282), .o1(\s[30] ));
  xnrc02aa1n02x5               g188(.a(\b[30] ), .b(\a[31] ), .out0(new_n284));
  norb02aa1n02x5               g189(.a(new_n276), .b(new_n279), .out0(new_n285));
  aobi12aa1n06x5               g190(.a(new_n285), .b(new_n249), .c(new_n251), .out0(new_n286));
  oao003aa1n02x5               g191(.a(\a[30] ), .b(\b[29] ), .c(new_n278), .carry(new_n287));
  nano22aa1n03x7               g192(.a(new_n286), .b(new_n284), .c(new_n287), .out0(new_n288));
  oaih12aa1n02x5               g193(.a(new_n285), .b(new_n263), .c(new_n260), .o1(new_n289));
  aoi012aa1n02x5               g194(.a(new_n284), .b(new_n289), .c(new_n287), .o1(new_n290));
  norp02aa1n03x5               g195(.a(new_n290), .b(new_n288), .o1(\s[31] ));
  xnrb03aa1n02x5               g196(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g197(.a(\a[3] ), .b(\b[2] ), .c(new_n104), .o1(new_n293));
  xorb03aa1n02x5               g198(.a(new_n293), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g199(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g200(.a(new_n109), .b(new_n107), .out0(new_n296));
  xobna2aa1n03x5               g201(.a(new_n108), .b(new_n296), .c(new_n116), .out0(\s[6] ));
  norp02aa1n02x5               g202(.a(new_n109), .b(new_n108), .o1(new_n298));
  aoi012aa1n02x5               g203(.a(new_n117), .b(new_n107), .c(new_n298), .o1(new_n299));
  xnrb03aa1n02x5               g204(.a(new_n299), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g205(.a(\a[7] ), .b(\b[6] ), .c(new_n299), .o1(new_n301));
  xorb03aa1n02x5               g206(.a(new_n301), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g207(.a(new_n120), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


