// Benchmark "adder" written by ABC on Wed Jul 17 16:18:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n337, new_n340,
    new_n342, new_n343, new_n344, new_n345, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv040aa1d32x5               g001(.a(\a[10] ), .o1(new_n97));
  nor022aa1n16x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  and002aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n02x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor002aa1d24x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano23aa1n02x4               g009(.a(new_n101), .b(new_n103), .c(new_n104), .d(new_n102), .out0(new_n105));
  inv000aa1n03x5               g010(.a(new_n103), .o1(new_n106));
  tech160nm_fioaoi03aa1n05x5   g011(.a(\a[4] ), .b(\b[3] ), .c(new_n106), .o1(new_n107));
  aoi012aa1n03x5               g012(.a(new_n107), .b(new_n105), .c(new_n100), .o1(new_n108));
  nor042aa1n12x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nanp02aa1n04x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nanb02aa1n03x5               g015(.a(new_n109), .b(new_n110), .out0(new_n111));
  nor002aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand02aa1d28x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nanb02aa1n09x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  nor002aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nand02aa1n08x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor002aa1d24x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand02aa1d10x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nano23aa1n02x4               g023(.a(new_n115), .b(new_n117), .c(new_n118), .d(new_n116), .out0(new_n119));
  nona22aa1n02x4               g024(.a(new_n119), .b(new_n114), .c(new_n111), .out0(new_n120));
  inv000aa1d42x5               g025(.a(\b[6] ), .o1(new_n121));
  nanb02aa1n02x5               g026(.a(\a[7] ), .b(new_n121), .out0(new_n122));
  aoai13aa1n06x5               g027(.a(new_n116), .b(new_n112), .c(new_n109), .d(new_n113), .o1(new_n123));
  nand22aa1n03x5               g028(.a(new_n123), .b(new_n122), .o1(new_n124));
  aoi012aa1n12x5               g029(.a(new_n117), .b(new_n124), .c(new_n118), .o1(new_n125));
  tech160nm_fioai012aa1n04x5   g030(.a(new_n125), .b(new_n108), .c(new_n120), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  aoi012aa1n02x5               g032(.a(new_n98), .b(new_n126), .c(new_n127), .o1(new_n128));
  xorb03aa1n02x5               g033(.a(new_n128), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  inv020aa1n08x5               g034(.a(\a[1] ), .o1(new_n130));
  inv040aa1d32x5               g035(.a(\b[0] ), .o1(new_n131));
  nor022aa1n12x5               g036(.a(\b[1] ), .b(\a[2] ), .o1(new_n132));
  nand02aa1n03x5               g037(.a(\b[1] ), .b(\a[2] ), .o1(new_n133));
  oaoi13aa1n12x5               g038(.a(new_n132), .b(new_n133), .c(new_n130), .d(new_n131), .o1(new_n134));
  nona23aa1d18x5               g039(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n135));
  oabi12aa1n18x5               g040(.a(new_n107), .b(new_n135), .c(new_n134), .out0(new_n136));
  nona23aa1d18x5               g041(.a(new_n118), .b(new_n116), .c(new_n115), .d(new_n117), .out0(new_n137));
  nor043aa1n09x5               g042(.a(new_n137), .b(new_n114), .c(new_n111), .o1(new_n138));
  nanp02aa1n09x5               g043(.a(new_n136), .b(new_n138), .o1(new_n139));
  tech160nm_fixorc02aa1n03p5x5 g044(.a(\a[10] ), .b(\b[9] ), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n127), .b(new_n140), .o1(new_n141));
  inv040aa1d32x5               g046(.a(\b[9] ), .o1(new_n142));
  oaoi03aa1n12x5               g047(.a(new_n97), .b(new_n142), .c(new_n98), .o1(new_n143));
  aoai13aa1n03x5               g048(.a(new_n143), .b(new_n141), .c(new_n139), .d(new_n125), .o1(new_n144));
  xorb03aa1n02x5               g049(.a(new_n144), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g050(.a(\a[12] ), .o1(new_n146));
  nor002aa1d24x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  nand42aa1n08x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  aoi012aa1n03x5               g053(.a(new_n147), .b(new_n144), .c(new_n148), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[11] ), .c(new_n146), .out0(\s[12] ));
  inv000aa1d42x5               g055(.a(new_n117), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n118), .o1(new_n152));
  aoai13aa1n06x5               g057(.a(new_n151), .b(new_n152), .c(new_n123), .d(new_n122), .o1(new_n153));
  nor002aa1d32x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  nand02aa1d24x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nona23aa1d18x5               g060(.a(new_n155), .b(new_n148), .c(new_n147), .d(new_n154), .out0(new_n156));
  nano22aa1n02x5               g061(.a(new_n156), .b(new_n140), .c(new_n127), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n153), .c(new_n136), .d(new_n138), .o1(new_n158));
  aoi012aa1n09x5               g063(.a(new_n154), .b(new_n147), .c(new_n155), .o1(new_n159));
  oai012aa1d24x5               g064(.a(new_n159), .b(new_n156), .c(new_n143), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  nanp02aa1n02x5               g066(.a(new_n158), .b(new_n161), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv000aa1d42x5               g068(.a(\a[14] ), .o1(new_n164));
  norp02aa1n24x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nand02aa1d20x5               g070(.a(\b[12] ), .b(\a[13] ), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n165), .b(new_n162), .c(new_n166), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[13] ), .c(new_n164), .out0(\s[14] ));
  nor002aa1d32x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1d16x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nona23aa1n09x5               g075(.a(new_n170), .b(new_n166), .c(new_n165), .d(new_n169), .out0(new_n171));
  aoi012aa1n12x5               g076(.a(new_n169), .b(new_n165), .c(new_n170), .o1(new_n172));
  aoai13aa1n06x5               g077(.a(new_n172), .b(new_n171), .c(new_n158), .d(new_n161), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  tech160nm_fixorc02aa1n04x5   g080(.a(\a[15] ), .b(\b[14] ), .out0(new_n176));
  xnrc02aa1n12x5               g081(.a(\b[15] ), .b(\a[16] ), .out0(new_n177));
  aoai13aa1n03x5               g082(.a(new_n177), .b(new_n175), .c(new_n173), .d(new_n176), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(new_n173), .b(new_n176), .o1(new_n179));
  nona22aa1n02x4               g084(.a(new_n179), .b(new_n177), .c(new_n175), .out0(new_n180));
  nanp02aa1n02x5               g085(.a(new_n180), .b(new_n178), .o1(\s[16] ));
  nano23aa1n06x5               g086(.a(new_n147), .b(new_n154), .c(new_n155), .d(new_n148), .out0(new_n182));
  nano23aa1n03x7               g087(.a(new_n165), .b(new_n169), .c(new_n170), .d(new_n166), .out0(new_n183));
  xorc02aa1n02x5               g088(.a(\a[16] ), .b(\b[15] ), .out0(new_n184));
  nand23aa1n03x5               g089(.a(new_n183), .b(new_n176), .c(new_n184), .o1(new_n185));
  nano32aa1n03x7               g090(.a(new_n185), .b(new_n182), .c(new_n127), .d(new_n140), .out0(new_n186));
  aoai13aa1n12x5               g091(.a(new_n186), .b(new_n153), .c(new_n136), .d(new_n138), .o1(new_n187));
  xnrc02aa1n12x5               g092(.a(\b[14] ), .b(\a[15] ), .out0(new_n188));
  norp03aa1d12x5               g093(.a(new_n171), .b(new_n188), .c(new_n177), .o1(new_n189));
  orn002aa1n03x5               g094(.a(\a[15] ), .b(\b[14] ), .o(new_n190));
  oao003aa1n06x5               g095(.a(\a[16] ), .b(\b[15] ), .c(new_n190), .carry(new_n191));
  oai013aa1d12x5               g096(.a(new_n191), .b(new_n188), .c(new_n177), .d(new_n172), .o1(new_n192));
  aoi012aa1d24x5               g097(.a(new_n192), .b(new_n160), .c(new_n189), .o1(new_n193));
  xorc02aa1n02x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n187), .c(new_n193), .out0(\s[17] ));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  nand22aa1n02x5               g101(.a(new_n157), .b(new_n189), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n193), .b(new_n197), .c(new_n139), .d(new_n125), .o1(new_n198));
  norp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  tech160nm_fiaoi012aa1n05x5   g104(.a(new_n199), .b(new_n198), .c(new_n194), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[17] ), .c(new_n196), .out0(\s[18] ));
  inv000aa1d42x5               g106(.a(\a[17] ), .o1(new_n202));
  xroi22aa1d06x4               g107(.a(new_n202), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n203));
  inv030aa1n02x5               g108(.a(new_n203), .o1(new_n204));
  nor042aa1n03x5               g109(.a(\b[17] ), .b(\a[18] ), .o1(new_n205));
  aoi112aa1n09x5               g110(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n206));
  norp02aa1n02x5               g111(.a(new_n206), .b(new_n205), .o1(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n204), .c(new_n187), .d(new_n193), .o1(new_n208));
  xorb03aa1n03x5               g113(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g114(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanp02aa1n04x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nor002aa1n16x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d28x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1d27x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n211), .c(new_n208), .d(new_n212), .o1(new_n217));
  inv000aa1n02x5               g122(.a(new_n207), .o1(new_n218));
  norb02aa1n09x5               g123(.a(new_n212), .b(new_n211), .out0(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n218), .c(new_n198), .d(new_n203), .o1(new_n220));
  nona22aa1n03x5               g125(.a(new_n220), .b(new_n216), .c(new_n211), .out0(new_n221));
  nanp02aa1n03x5               g126(.a(new_n217), .b(new_n221), .o1(\s[20] ));
  nano23aa1n06x5               g127(.a(new_n211), .b(new_n213), .c(new_n214), .d(new_n212), .out0(new_n223));
  nand02aa1d04x5               g128(.a(new_n203), .b(new_n223), .o1(new_n224));
  oai112aa1n06x5               g129(.a(new_n219), .b(new_n215), .c(new_n206), .d(new_n205), .o1(new_n225));
  aoi012aa1n06x5               g130(.a(new_n213), .b(new_n211), .c(new_n214), .o1(new_n226));
  nand02aa1d10x5               g131(.a(new_n225), .b(new_n226), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n224), .c(new_n187), .d(new_n193), .o1(new_n229));
  xorb03aa1n02x5               g134(.a(new_n229), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  nanp02aa1n06x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  nor042aa1n06x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  nand22aa1n12x5               g139(.a(\b[21] ), .b(\a[22] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n235), .b(new_n234), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n231), .c(new_n229), .d(new_n233), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n224), .o1(new_n239));
  aoai13aa1n03x5               g144(.a(new_n233), .b(new_n227), .c(new_n198), .d(new_n239), .o1(new_n240));
  nona22aa1n03x5               g145(.a(new_n240), .b(new_n237), .c(new_n231), .out0(new_n241));
  nanp02aa1n03x5               g146(.a(new_n238), .b(new_n241), .o1(\s[22] ));
  nano23aa1d12x5               g147(.a(new_n231), .b(new_n234), .c(new_n235), .d(new_n232), .out0(new_n243));
  nand23aa1d12x5               g148(.a(new_n203), .b(new_n223), .c(new_n243), .o1(new_n244));
  ao0012aa1n03x7               g149(.a(new_n234), .b(new_n231), .c(new_n235), .o(new_n245));
  tech160nm_fiaoi012aa1n05x5   g150(.a(new_n245), .b(new_n227), .c(new_n243), .o1(new_n246));
  aoai13aa1n04x5               g151(.a(new_n246), .b(new_n244), .c(new_n187), .d(new_n193), .o1(new_n247));
  nor042aa1n06x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  nand22aa1n12x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  inv030aa1n02x5               g155(.a(new_n244), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n246), .o1(new_n252));
  aoi112aa1n03x4               g157(.a(new_n250), .b(new_n252), .c(new_n198), .d(new_n251), .o1(new_n253));
  aoi012aa1n02x5               g158(.a(new_n253), .b(new_n247), .c(new_n250), .o1(\s[23] ));
  nor022aa1n16x5               g159(.a(\b[23] ), .b(\a[24] ), .o1(new_n255));
  nand22aa1n04x5               g160(.a(\b[23] ), .b(\a[24] ), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n03x5               g163(.a(new_n258), .b(new_n248), .c(new_n247), .d(new_n250), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n250), .b(new_n252), .c(new_n198), .d(new_n251), .o1(new_n260));
  nona22aa1n03x5               g165(.a(new_n260), .b(new_n258), .c(new_n248), .out0(new_n261));
  nanp02aa1n03x5               g166(.a(new_n259), .b(new_n261), .o1(\s[24] ));
  inv000aa1d42x5               g167(.a(new_n192), .o1(new_n263));
  aob012aa1n02x5               g168(.a(new_n263), .b(new_n160), .c(new_n189), .out0(new_n264));
  nano23aa1n09x5               g169(.a(new_n248), .b(new_n255), .c(new_n256), .d(new_n249), .out0(new_n265));
  nano32aa1n03x7               g170(.a(new_n204), .b(new_n265), .c(new_n223), .d(new_n243), .out0(new_n266));
  aoai13aa1n02x5               g171(.a(new_n266), .b(new_n264), .c(new_n126), .d(new_n186), .o1(new_n267));
  inv000aa1n02x5               g172(.a(new_n266), .o1(new_n268));
  nona23aa1n02x4               g173(.a(new_n235), .b(new_n232), .c(new_n231), .d(new_n234), .out0(new_n269));
  nona23aa1n02x4               g174(.a(new_n256), .b(new_n249), .c(new_n248), .d(new_n255), .out0(new_n270));
  nor042aa1n04x5               g175(.a(new_n269), .b(new_n270), .o1(new_n271));
  aoi112aa1n02x5               g176(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n272));
  nand42aa1n06x5               g177(.a(new_n265), .b(new_n245), .o1(new_n273));
  nona22aa1n12x5               g178(.a(new_n273), .b(new_n272), .c(new_n255), .out0(new_n274));
  aoi012aa1d24x5               g179(.a(new_n274), .b(new_n227), .c(new_n271), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n275), .b(new_n268), .c(new_n187), .d(new_n193), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  aoi112aa1n02x5               g182(.a(new_n274), .b(new_n277), .c(new_n227), .d(new_n271), .o1(new_n278));
  aoi022aa1n02x5               g183(.a(new_n276), .b(new_n277), .c(new_n267), .d(new_n278), .o1(\s[25] ));
  nor002aa1n02x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  xnrc02aa1n02x5               g185(.a(\b[25] ), .b(\a[26] ), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n280), .c(new_n276), .d(new_n277), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n275), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n277), .b(new_n283), .c(new_n198), .d(new_n266), .o1(new_n284));
  nona22aa1n03x5               g189(.a(new_n284), .b(new_n281), .c(new_n280), .out0(new_n285));
  nanp02aa1n03x5               g190(.a(new_n282), .b(new_n285), .o1(\s[26] ));
  norb02aa1n06x4               g191(.a(new_n277), .b(new_n281), .out0(new_n287));
  nano22aa1n06x5               g192(.a(new_n244), .b(new_n265), .c(new_n287), .out0(new_n288));
  inv020aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  nand22aa1n03x5               g194(.a(new_n265), .b(new_n243), .o1(new_n290));
  aoi012aa1n03x5               g195(.a(new_n290), .b(new_n225), .c(new_n226), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\a[26] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\b[25] ), .o1(new_n293));
  oaoi03aa1n02x5               g198(.a(new_n292), .b(new_n293), .c(new_n280), .o1(new_n294));
  inv000aa1n02x5               g199(.a(new_n294), .o1(new_n295));
  oaoi13aa1n09x5               g200(.a(new_n295), .b(new_n287), .c(new_n291), .d(new_n274), .o1(new_n296));
  aoai13aa1n09x5               g201(.a(new_n296), .b(new_n289), .c(new_n187), .d(new_n193), .o1(new_n297));
  xorb03aa1n03x5               g202(.a(new_n297), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  xorc02aa1n12x5               g204(.a(\a[27] ), .b(\b[26] ), .out0(new_n300));
  xnrc02aa1n12x5               g205(.a(\b[27] ), .b(\a[28] ), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n299), .c(new_n297), .d(new_n300), .o1(new_n302));
  oaib12aa1n12x5               g207(.a(new_n294), .b(new_n275), .c(new_n287), .out0(new_n303));
  aoai13aa1n04x5               g208(.a(new_n300), .b(new_n303), .c(new_n198), .d(new_n288), .o1(new_n304));
  nona22aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n299), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n302), .b(new_n305), .o1(\s[28] ));
  norb02aa1n03x5               g211(.a(new_n300), .b(new_n301), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n198), .d(new_n288), .o1(new_n308));
  aoai13aa1n06x5               g213(.a(new_n288), .b(new_n264), .c(new_n126), .d(new_n186), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n307), .o1(new_n310));
  orn002aa1n02x5               g215(.a(\a[27] ), .b(\b[26] ), .o(new_n311));
  oao003aa1n03x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n311), .carry(new_n312));
  aoai13aa1n02x7               g217(.a(new_n312), .b(new_n310), .c(new_n309), .d(new_n296), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .out0(new_n314));
  norb02aa1n02x5               g219(.a(new_n312), .b(new_n314), .out0(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n308), .d(new_n315), .o1(\s[29] ));
  xnrb03aa1n02x5               g221(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g222(.a(new_n301), .b(new_n314), .c(new_n300), .out0(new_n318));
  nanb02aa1n03x5               g223(.a(new_n318), .b(new_n297), .out0(new_n319));
  oaoi03aa1n09x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .o1(new_n320));
  inv000aa1n06x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n02x7               g226(.a(new_n321), .b(new_n318), .c(new_n309), .d(new_n296), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(\b[28] ), .b(\a[29] ), .o(new_n324));
  oabi12aa1n02x5               g229(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n325));
  oab012aa1n02x4               g230(.a(new_n325), .b(new_n312), .c(new_n324), .out0(new_n326));
  aoi022aa1n03x5               g231(.a(new_n322), .b(new_n323), .c(new_n319), .d(new_n326), .o1(\s[30] ));
  nanp03aa1n02x5               g232(.a(new_n307), .b(new_n314), .c(new_n323), .o1(new_n328));
  nanb02aa1n03x5               g233(.a(new_n328), .b(new_n297), .out0(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  oao003aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n331));
  norb02aa1n02x5               g236(.a(new_n331), .b(new_n330), .out0(new_n332));
  aoai13aa1n02x7               g237(.a(new_n331), .b(new_n328), .c(new_n309), .d(new_n296), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n333), .b(new_n330), .c(new_n329), .d(new_n332), .o1(\s[31] ));
  xnbna2aa1n03x5               g239(.a(new_n134), .b(new_n104), .c(new_n106), .out0(\s[3] ));
  inv000aa1d42x5               g240(.a(new_n101), .o1(new_n336));
  aoi122aa1n02x5               g241(.a(new_n103), .b(new_n336), .c(new_n102), .d(new_n100), .e(new_n104), .o1(new_n337));
  aoi012aa1n02x5               g242(.a(new_n337), .b(new_n336), .c(new_n136), .o1(\s[4] ));
  xorb03aa1n02x5               g243(.a(new_n136), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g244(.a(\a[5] ), .b(\b[4] ), .c(new_n108), .o1(new_n340));
  xnrc02aa1n02x5               g245(.a(new_n340), .b(new_n114), .out0(\s[6] ));
  inv000aa1d42x5               g246(.a(new_n113), .o1(new_n342));
  nanp02aa1n02x5               g247(.a(new_n122), .b(new_n116), .o1(new_n343));
  aoi112aa1n03x5               g248(.a(new_n109), .b(new_n114), .c(new_n136), .d(new_n110), .o1(new_n344));
  nano32aa1n03x7               g249(.a(new_n344), .b(new_n116), .c(new_n122), .d(new_n113), .out0(new_n345));
  oaoi13aa1n02x5               g250(.a(new_n345), .b(new_n343), .c(new_n342), .d(new_n344), .o1(\s[7] ));
  nor042aa1n03x5               g251(.a(new_n345), .b(new_n115), .o1(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n347), .b(new_n151), .c(new_n118), .out0(\s[8] ));
  xnbna2aa1n03x5               g253(.a(new_n127), .b(new_n139), .c(new_n125), .out0(\s[9] ));
endmodule


