// Benchmark "adder" written by ABC on Thu Jul 18 04:53:20 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n315, new_n318, new_n320,
    new_n321, new_n323;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  nand42aa1n10x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  norp02aa1n06x5               g003(.a(\b[8] ), .b(\a[9] ), .o1(new_n99));
  and002aa1n03x5               g004(.a(\b[1] ), .b(\a[2] ), .o(new_n100));
  nor042aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n09x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  norp02aa1n03x5               g007(.a(new_n101), .b(new_n102), .o1(new_n103));
  nor002aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand42aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n02x7               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor042aa1n04x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nona23aa1n06x5               g014(.a(new_n106), .b(new_n109), .c(new_n103), .d(new_n100), .out0(new_n110));
  tech160nm_fioai012aa1n03p5x5 g015(.a(new_n105), .b(new_n107), .c(new_n104), .o1(new_n111));
  nor022aa1n16x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand22aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n16x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n09x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nand42aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1n04x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  inv040aa1d32x5               g024(.a(\a[5] ), .o1(new_n120));
  inv000aa1d48x5               g025(.a(\b[4] ), .o1(new_n121));
  nand22aa1n04x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  nand42aa1n02x5               g028(.a(new_n122), .b(new_n123), .o1(new_n124));
  nona22aa1n03x5               g029(.a(new_n116), .b(new_n119), .c(new_n124), .out0(new_n125));
  oaoi03aa1n02x5               g030(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n126));
  inv000aa1d42x5               g031(.a(\a[7] ), .o1(new_n127));
  inv000aa1d42x5               g032(.a(\b[6] ), .o1(new_n128));
  aoai13aa1n02x7               g033(.a(new_n113), .b(new_n112), .c(new_n127), .d(new_n128), .o1(new_n129));
  aobi12aa1n06x5               g034(.a(new_n129), .b(new_n116), .c(new_n126), .out0(new_n130));
  aoai13aa1n12x5               g035(.a(new_n130), .b(new_n125), .c(new_n110), .d(new_n111), .o1(new_n131));
  tech160nm_fioai012aa1n05x5   g036(.a(new_n98), .b(new_n131), .c(new_n99), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  oaoi03aa1n02x5               g038(.a(\a[10] ), .b(\b[9] ), .c(new_n132), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand42aa1n06x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  nor042aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand42aa1n06x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n136), .c(new_n134), .d(new_n138), .o1(new_n142));
  nand42aa1n08x5               g047(.a(\b[9] ), .b(\a[10] ), .o1(new_n143));
  oaib12aa1n02x5               g048(.a(new_n132), .b(\b[9] ), .c(new_n97), .out0(new_n144));
  nanp03aa1n02x5               g049(.a(new_n144), .b(new_n143), .c(new_n138), .o1(new_n145));
  nona22aa1n02x4               g050(.a(new_n145), .b(new_n141), .c(new_n136), .out0(new_n146));
  nanp02aa1n02x5               g051(.a(new_n142), .b(new_n146), .o1(\s[12] ));
  nano23aa1d15x5               g052(.a(new_n136), .b(new_n139), .c(new_n140), .d(new_n137), .out0(new_n148));
  nor042aa1n06x5               g053(.a(\b[9] ), .b(\a[10] ), .o1(new_n149));
  tech160nm_fioai012aa1n05x5   g054(.a(new_n143), .b(new_n99), .c(new_n149), .o1(new_n150));
  inv040aa1n03x5               g055(.a(new_n150), .o1(new_n151));
  tech160nm_fioai012aa1n04x5   g056(.a(new_n140), .b(new_n139), .c(new_n136), .o1(new_n152));
  aobi12aa1n06x5               g057(.a(new_n152), .b(new_n148), .c(new_n151), .out0(new_n153));
  nano23aa1n06x5               g058(.a(new_n99), .b(new_n149), .c(new_n143), .d(new_n98), .out0(new_n154));
  nanp02aa1n02x5               g059(.a(new_n154), .b(new_n148), .o1(new_n155));
  nanb02aa1n06x5               g060(.a(new_n155), .b(new_n131), .out0(new_n156));
  nanp02aa1n06x5               g061(.a(new_n156), .b(new_n153), .o1(new_n157));
  xorb03aa1n02x5               g062(.a(new_n157), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n09x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand42aa1d28x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  tech160nm_fiaoi012aa1n05x5   g065(.a(new_n159), .b(new_n157), .c(new_n160), .o1(new_n161));
  xnrb03aa1n03x5               g066(.a(new_n161), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  nand42aa1n20x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nano23aa1d15x5               g069(.a(new_n159), .b(new_n163), .c(new_n164), .d(new_n160), .out0(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  aoi012aa1n02x5               g071(.a(new_n163), .b(new_n159), .c(new_n164), .o1(new_n167));
  aoai13aa1n04x5               g072(.a(new_n167), .b(new_n166), .c(new_n156), .d(new_n153), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor022aa1n08x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nand02aa1d16x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  nor002aa1n04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand02aa1d08x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  aoai13aa1n03x5               g080(.a(new_n175), .b(new_n170), .c(new_n168), .d(new_n172), .o1(new_n176));
  nanp02aa1n02x5               g081(.a(new_n168), .b(new_n172), .o1(new_n177));
  nona22aa1n02x4               g082(.a(new_n177), .b(new_n175), .c(new_n170), .out0(new_n178));
  nanp02aa1n03x5               g083(.a(new_n178), .b(new_n176), .o1(\s[16] ));
  oabi12aa1n12x5               g084(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n180));
  nona23aa1n03x5               g085(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n181));
  oai012aa1n06x5               g086(.a(new_n111), .b(new_n181), .c(new_n180), .o1(new_n182));
  nona23aa1n02x5               g087(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n183));
  nor043aa1n03x5               g088(.a(new_n183), .b(new_n119), .c(new_n124), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n117), .b(new_n118), .c(new_n121), .d(new_n120), .o1(new_n185));
  oaih12aa1n02x5               g090(.a(new_n129), .b(new_n183), .c(new_n185), .o1(new_n186));
  nano23aa1n09x5               g091(.a(new_n170), .b(new_n173), .c(new_n174), .d(new_n171), .out0(new_n187));
  nand22aa1n09x5               g092(.a(new_n187), .b(new_n165), .o1(new_n188));
  nano22aa1d15x5               g093(.a(new_n188), .b(new_n148), .c(new_n154), .out0(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n186), .c(new_n182), .d(new_n184), .o1(new_n190));
  nona23aa1n03x5               g095(.a(new_n140), .b(new_n137), .c(new_n136), .d(new_n139), .out0(new_n191));
  tech160nm_fioai012aa1n04x5   g096(.a(new_n152), .b(new_n191), .c(new_n150), .o1(new_n192));
  oa0012aa1n02x5               g097(.a(new_n164), .b(new_n163), .c(new_n159), .o(new_n193));
  oai012aa1n02x5               g098(.a(new_n174), .b(new_n173), .c(new_n170), .o1(new_n194));
  aob012aa1n06x5               g099(.a(new_n194), .b(new_n187), .c(new_n193), .out0(new_n195));
  aoib12aa1n12x5               g100(.a(new_n195), .b(new_n192), .c(new_n188), .out0(new_n196));
  xorc02aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n190), .c(new_n196), .out0(\s[17] ));
  inv040aa1d32x5               g103(.a(\a[18] ), .o1(new_n199));
  nanp02aa1n06x5               g104(.a(new_n190), .b(new_n196), .o1(new_n200));
  nor042aa1n03x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  tech160nm_fiaoi012aa1n05x5   g106(.a(new_n201), .b(new_n200), .c(new_n197), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[17] ), .c(new_n199), .out0(\s[18] ));
  inv000aa1d42x5               g108(.a(\a[17] ), .o1(new_n204));
  xroi22aa1d06x4               g109(.a(new_n204), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[17] ), .o1(new_n207));
  oaoi03aa1n09x5               g112(.a(new_n199), .b(new_n207), .c(new_n201), .o1(new_n208));
  aoai13aa1n04x5               g113(.a(new_n208), .b(new_n206), .c(new_n190), .d(new_n196), .o1(new_n209));
  xorb03aa1n02x5               g114(.a(new_n209), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nand02aa1n06x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nor042aa1n06x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand42aa1n04x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nanb02aa1n02x5               g120(.a(new_n214), .b(new_n215), .out0(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n212), .c(new_n209), .d(new_n213), .o1(new_n217));
  aoi112aa1n03x4               g122(.a(new_n212), .b(new_n216), .c(new_n209), .d(new_n213), .o1(new_n218));
  nanb02aa1n03x5               g123(.a(new_n218), .b(new_n217), .out0(\s[20] ));
  nona23aa1d18x5               g124(.a(new_n215), .b(new_n213), .c(new_n212), .d(new_n214), .out0(new_n220));
  oa0012aa1n06x5               g125(.a(new_n215), .b(new_n214), .c(new_n212), .o(new_n221));
  inv000aa1n09x5               g126(.a(new_n221), .o1(new_n222));
  oai012aa1d24x5               g127(.a(new_n222), .b(new_n220), .c(new_n208), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  nano23aa1n09x5               g129(.a(new_n212), .b(new_n214), .c(new_n215), .d(new_n213), .out0(new_n225));
  nanp02aa1n02x5               g130(.a(new_n205), .b(new_n225), .o1(new_n226));
  aoai13aa1n04x5               g131(.a(new_n224), .b(new_n226), .c(new_n190), .d(new_n196), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  tech160nm_fixnrc02aa1n05x5   g136(.a(\b[21] ), .b(\a[22] ), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n229), .c(new_n227), .d(new_n231), .o1(new_n233));
  aoi112aa1n03x4               g138(.a(new_n229), .b(new_n232), .c(new_n227), .d(new_n231), .o1(new_n234));
  nanb02aa1n03x5               g139(.a(new_n234), .b(new_n233), .out0(\s[22] ));
  nor042aa1n06x5               g140(.a(new_n232), .b(new_n230), .o1(new_n236));
  orn002aa1n02x5               g141(.a(\a[21] ), .b(\b[20] ), .o(new_n237));
  oao003aa1n02x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n237), .carry(new_n238));
  aobi12aa1n09x5               g143(.a(new_n238), .b(new_n223), .c(new_n236), .out0(new_n239));
  nand23aa1n06x5               g144(.a(new_n205), .b(new_n236), .c(new_n225), .o1(new_n240));
  aoai13aa1n04x5               g145(.a(new_n239), .b(new_n240), .c(new_n190), .d(new_n196), .o1(new_n241));
  xorb03aa1n02x5               g146(.a(new_n241), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  tech160nm_fixnrc02aa1n02p5x5 g149(.a(\b[23] ), .b(\a[24] ), .out0(new_n245));
  aoai13aa1n03x5               g150(.a(new_n245), .b(new_n243), .c(new_n241), .d(new_n244), .o1(new_n246));
  aoi112aa1n03x4               g151(.a(new_n243), .b(new_n245), .c(new_n241), .d(new_n244), .o1(new_n247));
  nanb02aa1n03x5               g152(.a(new_n247), .b(new_n246), .out0(\s[24] ));
  aobi12aa1n02x5               g153(.a(new_n194), .b(new_n187), .c(new_n193), .out0(new_n249));
  tech160nm_fioai012aa1n05x5   g154(.a(new_n249), .b(new_n153), .c(new_n188), .o1(new_n250));
  norb02aa1n03x4               g155(.a(new_n244), .b(new_n245), .out0(new_n251));
  inv030aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  nano32aa1n03x7               g157(.a(new_n252), .b(new_n205), .c(new_n236), .d(new_n225), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n250), .c(new_n131), .d(new_n189), .o1(new_n254));
  oao003aa1n02x5               g159(.a(new_n199), .b(new_n207), .c(new_n201), .carry(new_n255));
  aoai13aa1n06x5               g160(.a(new_n236), .b(new_n221), .c(new_n225), .d(new_n255), .o1(new_n256));
  oai022aa1n02x5               g161(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n257));
  aob012aa1n02x5               g162(.a(new_n257), .b(\b[23] ), .c(\a[24] ), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n252), .c(new_n256), .d(new_n238), .o1(new_n259));
  nanb02aa1n06x5               g164(.a(new_n259), .b(new_n254), .out0(new_n260));
  xorb03aa1n02x5               g165(.a(new_n260), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  xorc02aa1n03x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  xnrc02aa1n12x5               g168(.a(\b[25] ), .b(\a[26] ), .out0(new_n264));
  aoai13aa1n03x5               g169(.a(new_n264), .b(new_n262), .c(new_n260), .d(new_n263), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n263), .b(new_n259), .c(new_n200), .d(new_n253), .o1(new_n266));
  nona22aa1n02x5               g171(.a(new_n266), .b(new_n264), .c(new_n262), .out0(new_n267));
  nanp02aa1n03x5               g172(.a(new_n265), .b(new_n267), .o1(\s[26] ));
  norb02aa1n09x5               g173(.a(new_n263), .b(new_n264), .out0(new_n269));
  nand42aa1n03x5               g174(.a(new_n259), .b(new_n269), .o1(new_n270));
  nano22aa1n03x7               g175(.a(new_n240), .b(new_n251), .c(new_n269), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n250), .c(new_n131), .d(new_n189), .o1(new_n272));
  oai022aa1n02x5               g177(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n273));
  aob012aa1n02x5               g178(.a(new_n273), .b(\b[25] ), .c(\a[26] ), .out0(new_n274));
  nanp03aa1n06x5               g179(.a(new_n270), .b(new_n272), .c(new_n274), .o1(new_n275));
  xorb03aa1n02x5               g180(.a(new_n275), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xnrc02aa1n02x5               g183(.a(\b[27] ), .b(\a[28] ), .out0(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n277), .c(new_n275), .d(new_n278), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n269), .o1(new_n281));
  oaoi13aa1n04x5               g186(.a(new_n281), .b(new_n258), .c(new_n239), .d(new_n252), .o1(new_n282));
  inv020aa1n03x5               g187(.a(new_n271), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n274), .b(new_n283), .c(new_n190), .d(new_n196), .o1(new_n284));
  tech160nm_fioai012aa1n04x5   g189(.a(new_n278), .b(new_n284), .c(new_n282), .o1(new_n285));
  nona22aa1n02x5               g190(.a(new_n285), .b(new_n279), .c(new_n277), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n280), .b(new_n286), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n278), .b(new_n279), .out0(new_n288));
  oai012aa1n03x5               g193(.a(new_n288), .b(new_n284), .c(new_n282), .o1(new_n289));
  inv000aa1n03x5               g194(.a(new_n277), .o1(new_n290));
  oaoi03aa1n02x5               g195(.a(\a[28] ), .b(\b[27] ), .c(new_n290), .o1(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[28] ), .b(\a[29] ), .out0(new_n292));
  nona22aa1n02x5               g197(.a(new_n289), .b(new_n291), .c(new_n292), .out0(new_n293));
  aoai13aa1n03x5               g198(.a(new_n292), .b(new_n291), .c(new_n275), .d(new_n288), .o1(new_n294));
  nanp02aa1n03x5               g199(.a(new_n294), .b(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g201(.a(new_n278), .b(new_n292), .c(new_n279), .out0(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n290), .carry(new_n298));
  oaoi03aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .o1(new_n299));
  tech160nm_fixorc02aa1n03p5x5 g204(.a(\a[30] ), .b(\b[29] ), .out0(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n299), .c(new_n275), .d(new_n297), .o1(new_n302));
  oai012aa1n03x5               g207(.a(new_n297), .b(new_n284), .c(new_n282), .o1(new_n303));
  nona22aa1n02x5               g208(.a(new_n303), .b(new_n299), .c(new_n301), .out0(new_n304));
  nanp02aa1n03x5               g209(.a(new_n302), .b(new_n304), .o1(\s[30] ));
  nano23aa1n02x4               g210(.a(new_n292), .b(new_n279), .c(new_n300), .d(new_n278), .out0(new_n306));
  oai012aa1n03x5               g211(.a(new_n306), .b(new_n284), .c(new_n282), .o1(new_n307));
  nanp02aa1n02x5               g212(.a(new_n299), .b(new_n300), .o1(new_n308));
  oai012aa1n02x5               g213(.a(new_n308), .b(\b[29] ), .c(\a[30] ), .o1(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  nona22aa1n02x5               g215(.a(new_n307), .b(new_n309), .c(new_n310), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n310), .b(new_n309), .c(new_n275), .d(new_n306), .o1(new_n312));
  nanp02aa1n03x5               g217(.a(new_n312), .b(new_n311), .o1(\s[31] ));
  xnrc02aa1n02x5               g218(.a(new_n180), .b(new_n109), .out0(\s[3] ));
  oaoi03aa1n02x5               g219(.a(\a[3] ), .b(\b[2] ), .c(new_n180), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g221(.a(new_n182), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n02x5               g222(.a(new_n122), .b(new_n124), .c(new_n110), .d(new_n111), .o1(new_n318));
  xorb03aa1n02x5               g223(.a(new_n318), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  orn002aa1n02x5               g224(.a(new_n119), .b(new_n124), .o(new_n320));
  aoai13aa1n02x5               g225(.a(new_n185), .b(new_n320), .c(new_n110), .d(new_n111), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g227(.a(new_n127), .b(new_n128), .c(new_n321), .o1(new_n323));
  xnrb03aa1n02x5               g228(.a(new_n323), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g229(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


