// Benchmark "adder" written by ABC on Thu Jul 18 02:15:27 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n329, new_n331,
    new_n334, new_n335, new_n336, new_n338, new_n339, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand22aa1n09x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  oai112aa1n06x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .d(new_n100), .o1(new_n104));
  oa0022aa1n09x5               g009(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n105));
  aoi022aa1d18x5               g010(.a(new_n104), .b(new_n105), .c(\b[3] ), .d(\a[4] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nand02aa1d04x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nor042aa1n04x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  norb02aa1n02x5               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  nor042aa1n03x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor042aa1n04x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  nano22aa1n06x5               g022(.a(new_n117), .b(new_n109), .c(new_n112), .out0(new_n118));
  nanb02aa1n06x5               g023(.a(new_n107), .b(new_n108), .out0(new_n119));
  nanb02aa1n06x5               g024(.a(new_n110), .b(new_n111), .out0(new_n120));
  oai012aa1n02x7               g025(.a(new_n108), .b(new_n110), .c(new_n107), .o1(new_n121));
  tech160nm_fioai012aa1n05x5   g026(.a(new_n114), .b(new_n115), .c(new_n113), .o1(new_n122));
  oai013aa1n03x5               g027(.a(new_n121), .b(new_n122), .c(new_n119), .d(new_n120), .o1(new_n123));
  tech160nm_fixorc02aa1n04x5   g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n123), .c(new_n106), .d(new_n118), .o1(new_n125));
  nor002aa1d32x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand42aa1n08x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1d21x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n125), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g034(.a(new_n126), .o1(new_n130));
  inv000aa1d42x5               g035(.a(new_n128), .o1(new_n131));
  aoai13aa1n04x5               g036(.a(new_n130), .b(new_n131), .c(new_n125), .d(new_n99), .o1(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n16x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand22aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nor002aa1n20x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand42aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aoi112aa1n02x5               g043(.a(new_n134), .b(new_n138), .c(new_n132), .d(new_n135), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n138), .b(new_n134), .c(new_n132), .d(new_n135), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(\s[12] ));
  nona23aa1n09x5               g046(.a(new_n137), .b(new_n135), .c(new_n134), .d(new_n136), .out0(new_n142));
  nano22aa1n02x5               g047(.a(new_n142), .b(new_n124), .c(new_n128), .out0(new_n143));
  aoai13aa1n06x5               g048(.a(new_n143), .b(new_n123), .c(new_n106), .d(new_n118), .o1(new_n144));
  nano23aa1n06x5               g049(.a(new_n134), .b(new_n136), .c(new_n137), .d(new_n135), .out0(new_n145));
  tech160nm_fioai012aa1n03p5x5 g050(.a(new_n137), .b(new_n136), .c(new_n134), .o1(new_n146));
  aoai13aa1n12x5               g051(.a(new_n127), .b(new_n126), .c(new_n97), .d(new_n98), .o1(new_n147));
  inv000aa1n02x5               g052(.a(new_n147), .o1(new_n148));
  aobi12aa1n12x5               g053(.a(new_n146), .b(new_n145), .c(new_n148), .out0(new_n149));
  nanp02aa1n03x5               g054(.a(new_n144), .b(new_n149), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1n16x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand22aa1n03x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  aoi012aa1n02x5               g058(.a(new_n152), .b(new_n150), .c(new_n153), .o1(new_n154));
  xnrb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nand02aa1n06x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nona23aa1n12x5               g062(.a(new_n157), .b(new_n153), .c(new_n152), .d(new_n156), .out0(new_n158));
  oa0012aa1n02x5               g063(.a(new_n157), .b(new_n156), .c(new_n152), .o(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  aoai13aa1n04x5               g065(.a(new_n160), .b(new_n158), .c(new_n144), .d(new_n149), .o1(new_n161));
  xorb03aa1n02x5               g066(.a(new_n161), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  nanp02aa1n06x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nor042aa1n04x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nand42aa1n20x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  norb02aa1n12x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  aoi112aa1n02x5               g072(.a(new_n163), .b(new_n167), .c(new_n161), .d(new_n164), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n167), .b(new_n163), .c(new_n161), .d(new_n164), .o1(new_n169));
  norb02aa1n02x7               g074(.a(new_n169), .b(new_n168), .out0(\s[16] ));
  nand02aa1d04x5               g075(.a(new_n106), .b(new_n118), .o1(new_n171));
  nor003aa1n03x5               g076(.a(new_n122), .b(new_n119), .c(new_n120), .o1(new_n172));
  norb02aa1n03x5               g077(.a(new_n121), .b(new_n172), .out0(new_n173));
  norb02aa1n02x7               g078(.a(new_n164), .b(new_n163), .out0(new_n174));
  nano22aa1n12x5               g079(.a(new_n158), .b(new_n174), .c(new_n167), .out0(new_n175));
  nand02aa1d04x5               g080(.a(new_n143), .b(new_n175), .o1(new_n176));
  oai012aa1n06x5               g081(.a(new_n146), .b(new_n142), .c(new_n147), .o1(new_n177));
  oai112aa1n02x7               g082(.a(new_n157), .b(new_n164), .c(new_n156), .d(new_n152), .o1(new_n178));
  nona22aa1n03x5               g083(.a(new_n178), .b(new_n165), .c(new_n163), .out0(new_n179));
  aoi022aa1d18x5               g084(.a(new_n177), .b(new_n175), .c(new_n166), .d(new_n179), .o1(new_n180));
  aoai13aa1n12x5               g085(.a(new_n180), .b(new_n176), .c(new_n171), .d(new_n173), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nano23aa1n06x5               g087(.a(new_n152), .b(new_n156), .c(new_n157), .d(new_n153), .out0(new_n183));
  nand23aa1n03x5               g088(.a(new_n183), .b(new_n174), .c(new_n167), .o1(new_n184));
  nano32aa1n03x7               g089(.a(new_n184), .b(new_n145), .c(new_n128), .d(new_n124), .out0(new_n185));
  aoai13aa1n06x5               g090(.a(new_n185), .b(new_n123), .c(new_n106), .d(new_n118), .o1(new_n186));
  nor042aa1n06x5               g091(.a(\b[16] ), .b(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  xnrc02aa1n12x5               g093(.a(\b[16] ), .b(\a[17] ), .out0(new_n189));
  aoai13aa1n03x5               g094(.a(new_n188), .b(new_n189), .c(new_n186), .d(new_n180), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  tech160nm_fixnrc02aa1n04x5   g096(.a(\b[17] ), .b(\a[18] ), .out0(new_n192));
  nor042aa1n09x5               g097(.a(new_n192), .b(new_n189), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  oaoi03aa1n12x5               g099(.a(\a[18] ), .b(\b[17] ), .c(new_n188), .o1(new_n195));
  inv000aa1d42x5               g100(.a(new_n195), .o1(new_n196));
  aoai13aa1n04x5               g101(.a(new_n196), .b(new_n194), .c(new_n186), .d(new_n180), .o1(new_n197));
  xorb03aa1n02x5               g102(.a(new_n197), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g103(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n24x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand22aa1n09x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  xnrc02aa1n12x5               g106(.a(\b[19] ), .b(\a[20] ), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  aoi112aa1n03x4               g108(.a(new_n200), .b(new_n203), .c(new_n197), .d(new_n201), .o1(new_n204));
  inv000aa1d42x5               g109(.a(new_n200), .o1(new_n205));
  nanb02aa1d24x5               g110(.a(new_n200), .b(new_n201), .out0(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n207), .b(new_n195), .c(new_n181), .d(new_n193), .o1(new_n208));
  aoi012aa1n03x5               g113(.a(new_n202), .b(new_n208), .c(new_n205), .o1(new_n209));
  norp02aa1n03x5               g114(.a(new_n209), .b(new_n204), .o1(\s[20] ));
  nona22aa1n12x5               g115(.a(new_n193), .b(new_n206), .c(new_n202), .out0(new_n211));
  nanp02aa1n02x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  oaih22aa1d12x5               g117(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n213));
  nand23aa1n04x5               g118(.a(new_n213), .b(new_n212), .c(new_n201), .o1(new_n214));
  oab012aa1n09x5               g119(.a(new_n200), .b(\a[20] ), .c(\b[19] ), .out0(new_n215));
  aoi022aa1d18x5               g120(.a(new_n214), .b(new_n215), .c(\b[19] ), .d(\a[20] ), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n211), .c(new_n186), .d(new_n180), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  nand42aa1n03x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  nor022aa1n16x5               g127(.a(\b[21] ), .b(\a[22] ), .o1(new_n223));
  nanp02aa1n04x5               g128(.a(\b[21] ), .b(\a[22] ), .o1(new_n224));
  norb02aa1n09x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  aoi112aa1n03x4               g130(.a(new_n220), .b(new_n225), .c(new_n218), .d(new_n222), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n220), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n211), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n222), .b(new_n216), .c(new_n181), .d(new_n228), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n225), .o1(new_n230));
  tech160nm_fiaoi012aa1n02p5x5 g135(.a(new_n230), .b(new_n229), .c(new_n227), .o1(new_n231));
  nor002aa1n02x5               g136(.a(new_n231), .b(new_n226), .o1(\s[22] ));
  nona23aa1d18x5               g137(.a(new_n224), .b(new_n221), .c(new_n220), .d(new_n223), .out0(new_n233));
  nona23aa1d24x5               g138(.a(new_n193), .b(new_n203), .c(new_n233), .d(new_n206), .out0(new_n234));
  and002aa1n02x5               g139(.a(\b[19] ), .b(\a[20] ), .o(new_n235));
  aoi112aa1n06x5               g140(.a(new_n233), .b(new_n235), .c(new_n214), .d(new_n215), .o1(new_n236));
  tech160nm_fioai012aa1n04x5   g141(.a(new_n224), .b(new_n223), .c(new_n220), .o1(new_n237));
  norb02aa1n12x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n234), .c(new_n186), .d(new_n180), .o1(new_n239));
  xorb03aa1n02x5               g144(.a(new_n239), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n04x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  xnrc02aa1n12x5               g146(.a(\b[22] ), .b(\a[23] ), .out0(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[23] ), .b(\a[24] ), .out0(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  aoi112aa1n03x4               g150(.a(new_n241), .b(new_n245), .c(new_n239), .d(new_n243), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n241), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n234), .o1(new_n248));
  inv040aa1n03x5               g153(.a(new_n238), .o1(new_n249));
  aoai13aa1n03x5               g154(.a(new_n243), .b(new_n249), .c(new_n181), .d(new_n248), .o1(new_n250));
  aoi012aa1n03x5               g155(.a(new_n244), .b(new_n250), .c(new_n247), .o1(new_n251));
  norp02aa1n03x5               g156(.a(new_n251), .b(new_n246), .o1(\s[24] ));
  nor042aa1n09x5               g157(.a(new_n244), .b(new_n242), .o1(new_n253));
  nano32aa1n06x5               g158(.a(new_n211), .b(new_n253), .c(new_n222), .d(new_n225), .out0(new_n254));
  inv040aa1n03x5               g159(.a(new_n254), .o1(new_n255));
  tech160nm_finand02aa1n03p5x5 g160(.a(new_n214), .b(new_n215), .o1(new_n256));
  nona23aa1n08x5               g161(.a(new_n256), .b(new_n253), .c(new_n233), .d(new_n235), .out0(new_n257));
  orn002aa1n02x5               g162(.a(\a[24] ), .b(\b[23] ), .o(new_n258));
  aob012aa1n02x5               g163(.a(new_n241), .b(\b[23] ), .c(\a[24] ), .out0(new_n259));
  nor003aa1n04x5               g164(.a(new_n244), .b(new_n242), .c(new_n237), .o1(new_n260));
  nano22aa1n03x7               g165(.a(new_n260), .b(new_n258), .c(new_n259), .out0(new_n261));
  nand22aa1n12x5               g166(.a(new_n257), .b(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n255), .c(new_n186), .d(new_n180), .o1(new_n264));
  xorb03aa1n02x5               g169(.a(new_n264), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  xorc02aa1n12x5               g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  xorc02aa1n12x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  aoi112aa1n03x4               g173(.a(new_n266), .b(new_n268), .c(new_n264), .d(new_n267), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n266), .o1(new_n270));
  aoai13aa1n03x5               g175(.a(new_n267), .b(new_n262), .c(new_n181), .d(new_n254), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n268), .o1(new_n272));
  aoi012aa1n02x7               g177(.a(new_n272), .b(new_n271), .c(new_n270), .o1(new_n273));
  nor002aa1n02x5               g178(.a(new_n273), .b(new_n269), .o1(\s[26] ));
  nanp02aa1n02x5               g179(.a(\b[3] ), .b(\a[4] ), .o1(new_n275));
  nanp02aa1n02x5               g180(.a(new_n104), .b(new_n105), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(new_n276), .b(new_n275), .o1(new_n277));
  nano23aa1n02x4               g182(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n278));
  nona22aa1n02x4               g183(.a(new_n278), .b(new_n119), .c(new_n120), .out0(new_n279));
  oai012aa1n02x7               g184(.a(new_n173), .b(new_n277), .c(new_n279), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(new_n179), .b(new_n166), .o1(new_n281));
  tech160nm_fioai012aa1n04x5   g186(.a(new_n281), .b(new_n149), .c(new_n184), .o1(new_n282));
  and002aa1n24x5               g187(.a(new_n268), .b(new_n267), .o(new_n283));
  nano22aa1d15x5               g188(.a(new_n234), .b(new_n283), .c(new_n253), .out0(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n282), .c(new_n280), .d(new_n185), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .c(new_n270), .carry(new_n286));
  aobi12aa1n18x5               g191(.a(new_n286), .b(new_n262), .c(new_n283), .out0(new_n287));
  nor042aa1n06x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  nanb02aa1n06x5               g194(.a(new_n288), .b(new_n289), .out0(new_n290));
  xobna2aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n287), .out0(\s[27] ));
  inv000aa1d42x5               g196(.a(new_n288), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n283), .o1(new_n293));
  aoai13aa1n06x5               g198(.a(new_n286), .b(new_n293), .c(new_n257), .d(new_n261), .o1(new_n294));
  aoai13aa1n03x5               g199(.a(new_n289), .b(new_n294), .c(new_n181), .d(new_n284), .o1(new_n295));
  xnrc02aa1n12x5               g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  aoi012aa1n03x5               g201(.a(new_n296), .b(new_n295), .c(new_n292), .o1(new_n297));
  aoi022aa1n03x5               g202(.a(new_n285), .b(new_n287), .c(\b[26] ), .d(\a[27] ), .o1(new_n298));
  nano22aa1n03x5               g203(.a(new_n298), .b(new_n292), .c(new_n296), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[28] ));
  nor042aa1n03x5               g205(.a(new_n296), .b(new_n290), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n294), .c(new_n181), .d(new_n284), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  aoi012aa1n02x7               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n301), .o1(new_n306));
  tech160nm_fiaoi012aa1n02p5x5 g211(.a(new_n306), .b(new_n285), .c(new_n287), .o1(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n304), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n305), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nor043aa1n03x5               g215(.a(new_n304), .b(new_n296), .c(new_n290), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n294), .c(new_n181), .d(new_n284), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[29] ), .b(\a[30] ), .out0(new_n314));
  tech160nm_fiaoi012aa1n02p5x5 g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n316), .b(new_n285), .c(new_n287), .o1(new_n317));
  nano22aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n314), .out0(new_n318));
  norp02aa1n03x5               g223(.a(new_n315), .b(new_n318), .o1(\s[30] ));
  xnrc02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  norb03aa1n02x7               g225(.a(new_n301), .b(new_n314), .c(new_n304), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n294), .c(new_n181), .d(new_n284), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n323));
  aoi012aa1n03x5               g228(.a(new_n320), .b(new_n322), .c(new_n323), .o1(new_n324));
  inv000aa1n02x5               g229(.a(new_n321), .o1(new_n325));
  tech160nm_fiaoi012aa1n02p5x5 g230(.a(new_n325), .b(new_n285), .c(new_n287), .o1(new_n326));
  nano22aa1n03x5               g231(.a(new_n326), .b(new_n320), .c(new_n323), .out0(new_n327));
  norp02aa1n03x5               g232(.a(new_n324), .b(new_n327), .o1(\s[31] ));
  oai012aa1n02x5               g233(.a(new_n101), .b(new_n102), .c(new_n100), .o1(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g235(.a(\a[3] ), .b(\b[2] ), .c(new_n329), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g237(.a(new_n106), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g238(.a(new_n114), .b(new_n113), .out0(new_n334));
  oaoi13aa1n02x5               g239(.a(new_n334), .b(new_n116), .c(new_n106), .d(new_n115), .o1(new_n335));
  oai112aa1n03x5               g240(.a(new_n116), .b(new_n334), .c(new_n106), .d(new_n115), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n336), .b(new_n335), .out0(\s[6] ));
  oaoi13aa1n02x5               g242(.a(new_n120), .b(new_n336), .c(\a[6] ), .d(\b[5] ), .o1(new_n338));
  nona22aa1n02x4               g243(.a(new_n336), .b(new_n113), .c(new_n112), .out0(new_n339));
  norb02aa1n02x5               g244(.a(new_n339), .b(new_n338), .out0(\s[7] ));
  norp02aa1n03x5               g245(.a(new_n338), .b(new_n110), .o1(new_n341));
  xnrc02aa1n02x5               g246(.a(new_n341), .b(new_n109), .out0(\s[8] ));
  xnbna2aa1n03x5               g247(.a(new_n124), .b(new_n171), .c(new_n173), .out0(\s[9] ));
endmodule


