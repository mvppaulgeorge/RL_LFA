// Benchmark "adder" written by ABC on Wed Jul 17 15:28:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n309, new_n310,
    new_n313, new_n315, new_n317;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n05x5   g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  orn002aa1n02x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  nor042aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nand22aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor022aa1n12x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor022aa1n08x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n103), .b(new_n106), .c(new_n105), .d(new_n104), .out0(new_n107));
  tech160nm_fiaoi012aa1n04x5   g012(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n108));
  oai012aa1n12x5               g013(.a(new_n108), .b(new_n107), .c(new_n102), .o1(new_n109));
  xorc02aa1n12x5               g014(.a(\a[7] ), .b(\b[6] ), .out0(new_n110));
  nand42aa1n06x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  norp02aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanb02aa1n06x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nor042aa1n06x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nor022aa1n06x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand22aa1n12x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nona23aa1n09x5               g022(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n118));
  norb03aa1n12x5               g023(.a(new_n110), .b(new_n118), .c(new_n113), .out0(new_n119));
  nanp02aa1n02x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  orn002aa1n24x5               g025(.a(\a[7] ), .b(\b[6] ), .o(new_n121));
  tech160nm_finand02aa1n05x5   g026(.a(new_n114), .b(new_n117), .o1(new_n122));
  oai112aa1n06x5               g027(.a(new_n122), .b(new_n121), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  nanp03aa1n06x5               g028(.a(new_n123), .b(new_n120), .c(new_n111), .o1(new_n124));
  oai012aa1n12x5               g029(.a(new_n124), .b(\b[7] ), .c(\a[8] ), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n97), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  aobi12aa1n06x5               g033(.a(new_n97), .b(new_n127), .c(new_n98), .out0(new_n129));
  oai022aa1d24x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  aob012aa1d24x5               g035(.a(new_n130), .b(\b[9] ), .c(\a[10] ), .out0(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1d08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  tech160nm_fioai012aa1n04x5   g040(.a(new_n135), .b(new_n129), .c(new_n132), .o1(new_n136));
  norp03aa1n02x5               g041(.a(new_n129), .b(new_n132), .c(new_n135), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n136), .b(new_n137), .out0(\s[11] ));
  nor042aa1n06x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n09x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  nona22aa1n02x4               g046(.a(new_n136), .b(new_n141), .c(new_n133), .out0(new_n142));
  inv040aa1n04x5               g047(.a(new_n133), .o1(new_n143));
  aobi12aa1n06x5               g048(.a(new_n141), .b(new_n136), .c(new_n143), .out0(new_n144));
  norb02aa1n03x4               g049(.a(new_n142), .b(new_n144), .out0(\s[12] ));
  nanp02aa1n06x5               g050(.a(new_n119), .b(new_n109), .o1(new_n146));
  aoi013aa1n06x4               g051(.a(new_n112), .b(new_n123), .c(new_n120), .d(new_n111), .o1(new_n147));
  nano23aa1n06x5               g052(.a(new_n133), .b(new_n139), .c(new_n140), .d(new_n134), .out0(new_n148));
  nand23aa1n04x5               g053(.a(new_n148), .b(new_n97), .c(new_n126), .o1(new_n149));
  nona23aa1d16x5               g054(.a(new_n140), .b(new_n134), .c(new_n133), .d(new_n139), .out0(new_n150));
  oaoi03aa1n03x5               g055(.a(\a[12] ), .b(\b[11] ), .c(new_n143), .o1(new_n151));
  oabi12aa1n18x5               g056(.a(new_n151), .b(new_n150), .c(new_n131), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n06x5               g058(.a(new_n153), .b(new_n149), .c(new_n146), .d(new_n147), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n12x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand42aa1n16x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  aoi012aa1n02x5               g062(.a(new_n156), .b(new_n154), .c(new_n157), .o1(new_n158));
  xnrb03aa1n03x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1d18x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n10x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nano23aa1d15x5               g066(.a(new_n156), .b(new_n160), .c(new_n161), .d(new_n157), .out0(new_n162));
  oa0012aa1n02x5               g067(.a(new_n161), .b(new_n160), .c(new_n156), .o(new_n163));
  nor002aa1d32x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand42aa1n06x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nanb02aa1d36x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoai13aa1n06x5               g072(.a(new_n167), .b(new_n163), .c(new_n154), .d(new_n162), .o1(new_n168));
  aoi112aa1n02x5               g073(.a(new_n167), .b(new_n163), .c(new_n154), .d(new_n162), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(\s[15] ));
  inv000aa1d42x5               g075(.a(new_n164), .o1(new_n171));
  nor022aa1n16x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand42aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nanb02aa1n12x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  nanp03aa1n03x5               g079(.a(new_n168), .b(new_n171), .c(new_n174), .o1(new_n175));
  tech160nm_fiaoi012aa1n04x5   g080(.a(new_n174), .b(new_n168), .c(new_n171), .o1(new_n176));
  norb02aa1n03x4               g081(.a(new_n175), .b(new_n176), .out0(\s[16] ));
  nona22aa1n09x5               g082(.a(new_n162), .b(new_n166), .c(new_n174), .out0(new_n178));
  nor042aa1n06x5               g083(.a(new_n149), .b(new_n178), .o1(new_n179));
  aoai13aa1n12x5               g084(.a(new_n179), .b(new_n125), .c(new_n109), .d(new_n119), .o1(new_n180));
  nona23aa1n02x5               g085(.a(new_n161), .b(new_n157), .c(new_n156), .d(new_n160), .out0(new_n181));
  nor003aa1n03x5               g086(.a(new_n181), .b(new_n166), .c(new_n174), .o1(new_n182));
  oaoi13aa1n02x7               g087(.a(new_n164), .b(new_n161), .c(new_n156), .d(new_n160), .o1(new_n183));
  nano22aa1n03x5               g088(.a(new_n183), .b(new_n165), .c(new_n173), .out0(new_n184));
  aoi112aa1n09x5               g089(.a(new_n184), .b(new_n172), .c(new_n152), .d(new_n182), .o1(new_n185));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n180), .c(new_n185), .out0(\s[17] ));
  inv000aa1d42x5               g092(.a(\a[17] ), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[16] ), .o1(new_n189));
  nand42aa1n02x5               g094(.a(new_n189), .b(new_n188), .o1(new_n190));
  nand02aa1n04x5               g095(.a(new_n146), .b(new_n147), .o1(new_n191));
  nanp02aa1n02x5               g096(.a(new_n152), .b(new_n182), .o1(new_n192));
  nona22aa1n03x5               g097(.a(new_n192), .b(new_n184), .c(new_n172), .out0(new_n193));
  aoai13aa1n02x5               g098(.a(new_n186), .b(new_n193), .c(new_n191), .d(new_n179), .o1(new_n194));
  nor002aa1d32x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nand42aa1n08x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nanb02aa1n12x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  xobna2aa1n03x5               g102(.a(new_n197), .b(new_n194), .c(new_n190), .out0(\s[18] ));
  nanp02aa1n02x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  nano22aa1n12x5               g104(.a(new_n197), .b(new_n190), .c(new_n199), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n196), .b(new_n195), .c(new_n188), .d(new_n189), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n201), .c(new_n180), .d(new_n185), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand22aa1n09x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nor042aa1n06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand22aa1n09x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi112aa1n03x5               g115(.a(new_n206), .b(new_n210), .c(new_n203), .d(new_n207), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n210), .b(new_n206), .c(new_n203), .d(new_n207), .o1(new_n212));
  norb02aa1n03x4               g117(.a(new_n212), .b(new_n211), .out0(\s[20] ));
  nano23aa1n06x5               g118(.a(new_n206), .b(new_n208), .c(new_n209), .d(new_n207), .out0(new_n214));
  nanp02aa1n02x5               g119(.a(new_n200), .b(new_n214), .o1(new_n215));
  nona23aa1d18x5               g120(.a(new_n209), .b(new_n207), .c(new_n206), .d(new_n208), .out0(new_n216));
  aoi012aa1n12x5               g121(.a(new_n208), .b(new_n206), .c(new_n209), .o1(new_n217));
  oai012aa1d24x5               g122(.a(new_n217), .b(new_n216), .c(new_n202), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n06x5               g124(.a(new_n219), .b(new_n215), .c(new_n180), .d(new_n185), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[21] ), .b(\b[20] ), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[22] ), .b(\b[21] ), .out0(new_n224));
  aoi112aa1n03x5               g129(.a(new_n222), .b(new_n224), .c(new_n220), .d(new_n223), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n224), .b(new_n222), .c(new_n220), .d(new_n223), .o1(new_n226));
  norb02aa1n03x4               g131(.a(new_n226), .b(new_n225), .out0(\s[22] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  nand23aa1n02x5               g135(.a(new_n230), .b(new_n200), .c(new_n214), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\b[21] ), .o1(new_n232));
  oaoi03aa1n12x5               g137(.a(new_n229), .b(new_n232), .c(new_n222), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoi012aa1n02x5               g139(.a(new_n234), .b(new_n218), .c(new_n230), .o1(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n231), .c(new_n180), .d(new_n185), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  tech160nm_fixorc02aa1n02p5x5 g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  xorc02aa1n03x5               g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  aoi112aa1n02x5               g145(.a(new_n238), .b(new_n240), .c(new_n236), .d(new_n239), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n238), .c(new_n236), .d(new_n239), .o1(new_n242));
  norb02aa1n03x4               g147(.a(new_n242), .b(new_n241), .out0(\s[24] ));
  nanp02aa1n06x5               g148(.a(new_n180), .b(new_n185), .o1(new_n244));
  and002aa1n02x5               g149(.a(new_n240), .b(new_n239), .o(new_n245));
  inv000aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  nor002aa1n02x5               g151(.a(new_n231), .b(new_n246), .o1(new_n247));
  inv040aa1n03x5               g152(.a(new_n202), .o1(new_n248));
  inv040aa1n03x5               g153(.a(new_n217), .o1(new_n249));
  aoai13aa1n06x5               g154(.a(new_n230), .b(new_n249), .c(new_n214), .d(new_n248), .o1(new_n250));
  orn002aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .o(new_n251));
  oao003aa1n02x5               g156(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .carry(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n246), .c(new_n250), .d(new_n233), .o1(new_n253));
  xorc02aa1n12x5               g158(.a(\a[25] ), .b(\b[24] ), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n253), .c(new_n244), .d(new_n247), .o1(new_n255));
  aoi112aa1n02x5               g160(.a(new_n254), .b(new_n253), .c(new_n244), .d(new_n247), .o1(new_n256));
  norb02aa1n03x4               g161(.a(new_n255), .b(new_n256), .out0(\s[25] ));
  nor042aa1n03x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  tech160nm_fixorc02aa1n04x5   g163(.a(\a[26] ), .b(\b[25] ), .out0(new_n259));
  nona22aa1n02x5               g164(.a(new_n255), .b(new_n259), .c(new_n258), .out0(new_n260));
  inv000aa1d42x5               g165(.a(new_n258), .o1(new_n261));
  aobi12aa1n06x5               g166(.a(new_n259), .b(new_n255), .c(new_n261), .out0(new_n262));
  norb02aa1n03x4               g167(.a(new_n260), .b(new_n262), .out0(\s[26] ));
  and002aa1n06x5               g168(.a(new_n259), .b(new_n254), .o(new_n264));
  nano22aa1n03x7               g169(.a(new_n231), .b(new_n245), .c(new_n264), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n193), .c(new_n191), .d(new_n179), .o1(new_n266));
  oao003aa1n02x5               g171(.a(\a[26] ), .b(\b[25] ), .c(new_n261), .carry(new_n267));
  aobi12aa1n06x5               g172(.a(new_n267), .b(new_n253), .c(new_n264), .out0(new_n268));
  xorc02aa1n12x5               g173(.a(\a[27] ), .b(\b[26] ), .out0(new_n269));
  xnbna2aa1n03x5               g174(.a(new_n269), .b(new_n268), .c(new_n266), .out0(\s[27] ));
  norp02aa1n02x5               g175(.a(\b[26] ), .b(\a[27] ), .o1(new_n271));
  inv040aa1n03x5               g176(.a(new_n271), .o1(new_n272));
  aobi12aa1n03x5               g177(.a(new_n269), .b(new_n268), .c(new_n266), .out0(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[27] ), .b(\a[28] ), .out0(new_n274));
  nano22aa1n02x4               g179(.a(new_n273), .b(new_n272), .c(new_n274), .out0(new_n275));
  aobi12aa1n06x5               g180(.a(new_n265), .b(new_n180), .c(new_n185), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n245), .b(new_n234), .c(new_n218), .d(new_n230), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n264), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n267), .b(new_n278), .c(new_n277), .d(new_n252), .o1(new_n279));
  oaih12aa1n02x5               g184(.a(new_n269), .b(new_n279), .c(new_n276), .o1(new_n280));
  aoi012aa1n03x5               g185(.a(new_n274), .b(new_n280), .c(new_n272), .o1(new_n281));
  nor002aa1n02x5               g186(.a(new_n281), .b(new_n275), .o1(\s[28] ));
  norb02aa1n02x5               g187(.a(new_n269), .b(new_n274), .out0(new_n283));
  oaih12aa1n02x5               g188(.a(new_n283), .b(new_n279), .c(new_n276), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[28] ), .b(\b[27] ), .c(new_n272), .carry(new_n285));
  xnrc02aa1n02x5               g190(.a(\b[28] ), .b(\a[29] ), .out0(new_n286));
  aoi012aa1n03x5               g191(.a(new_n286), .b(new_n284), .c(new_n285), .o1(new_n287));
  aobi12aa1n06x5               g192(.a(new_n283), .b(new_n268), .c(new_n266), .out0(new_n288));
  nano22aa1n03x5               g193(.a(new_n288), .b(new_n285), .c(new_n286), .out0(new_n289));
  norp02aa1n03x5               g194(.a(new_n287), .b(new_n289), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g196(.a(new_n269), .b(new_n286), .c(new_n274), .out0(new_n292));
  oaih12aa1n02x5               g197(.a(new_n292), .b(new_n279), .c(new_n276), .o1(new_n293));
  oao003aa1n02x5               g198(.a(\a[29] ), .b(\b[28] ), .c(new_n285), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .out0(new_n295));
  aoi012aa1n03x5               g200(.a(new_n295), .b(new_n293), .c(new_n294), .o1(new_n296));
  aobi12aa1n02x7               g201(.a(new_n292), .b(new_n268), .c(new_n266), .out0(new_n297));
  nano22aa1n03x5               g202(.a(new_n297), .b(new_n294), .c(new_n295), .out0(new_n298));
  nor002aa1n02x5               g203(.a(new_n296), .b(new_n298), .o1(\s[30] ));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n292), .b(new_n295), .out0(new_n301));
  aobi12aa1n02x7               g206(.a(new_n301), .b(new_n268), .c(new_n266), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n294), .carry(new_n303));
  nano22aa1n03x5               g208(.a(new_n302), .b(new_n300), .c(new_n303), .out0(new_n304));
  oaih12aa1n02x5               g209(.a(new_n301), .b(new_n279), .c(new_n276), .o1(new_n305));
  aoi012aa1n03x5               g210(.a(new_n300), .b(new_n305), .c(new_n303), .o1(new_n306));
  norp02aa1n03x5               g211(.a(new_n306), .b(new_n304), .o1(\s[31] ));
  xnrb03aa1n02x5               g212(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nona22aa1n02x4               g213(.a(new_n106), .b(new_n102), .c(new_n105), .out0(new_n309));
  aoib12aa1n02x5               g214(.a(new_n105), .b(new_n103), .c(new_n104), .out0(new_n310));
  aboi22aa1n03x5               g215(.a(new_n104), .b(new_n109), .c(new_n309), .d(new_n310), .out0(\s[4] ));
  xorb03aa1n02x5               g216(.a(new_n109), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n03x5               g217(.a(new_n114), .b(new_n109), .c(new_n115), .o1(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb03aa1n02x5               g219(.a(new_n116), .b(new_n313), .c(new_n117), .out0(new_n315));
  xobna2aa1n03x5               g220(.a(new_n110), .b(new_n315), .c(new_n117), .out0(\s[7] ));
  nanp03aa1n02x5               g221(.a(new_n315), .b(new_n110), .c(new_n117), .o1(new_n317));
  xobna2aa1n03x5               g222(.a(new_n113), .b(new_n317), .c(new_n121), .out0(\s[8] ));
  xnbna2aa1n03x5               g223(.a(new_n126), .b(new_n146), .c(new_n147), .out0(\s[9] ));
endmodule


