// Benchmark "adder" written by ABC on Thu Jul 18 08:06:29 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n180, new_n181,
    new_n182, new_n183, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n326, new_n327,
    new_n328, new_n330, new_n331;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand02aa1d04x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nand02aa1d04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  aoi012aa1n06x5               g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  nor022aa1n06x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nanp02aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  tech160nm_fiaoi012aa1n03p5x5 g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  norp02aa1n09x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand22aa1n04x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand02aa1n03x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n09x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  nor022aa1n08x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nanp02aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nanb02aa1n02x5               g019(.a(new_n113), .b(new_n114), .out0(new_n115));
  tech160nm_fixnrc02aa1n04x5   g020(.a(\b[4] ), .b(\a[5] ), .out0(new_n116));
  nor043aa1n06x5               g021(.a(new_n112), .b(new_n115), .c(new_n116), .o1(new_n117));
  inv000aa1d42x5               g022(.a(\a[5] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[4] ), .o1(new_n119));
  aoai13aa1n02x5               g024(.a(new_n114), .b(new_n113), .c(new_n118), .d(new_n119), .o1(new_n120));
  aoi012aa1n02x7               g025(.a(new_n108), .b(new_n110), .c(new_n109), .o1(new_n121));
  oai012aa1n06x5               g026(.a(new_n121), .b(new_n112), .c(new_n120), .o1(new_n122));
  aoi012aa1n12x5               g027(.a(new_n122), .b(new_n107), .c(new_n117), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .c(new_n123), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1d32x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nand22aa1n04x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n126), .b(new_n127), .out0(new_n128));
  inv000aa1d42x5               g033(.a(\a[10] ), .o1(new_n129));
  inv000aa1d42x5               g034(.a(\b[8] ), .o1(new_n130));
  xroi22aa1d06x4               g035(.a(new_n129), .b(\b[9] ), .c(new_n130), .d(\a[9] ), .out0(new_n131));
  aoai13aa1n06x5               g036(.a(new_n131), .b(new_n122), .c(new_n107), .d(new_n117), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  oai022aa1d18x5               g038(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n134));
  nand02aa1n03x5               g039(.a(new_n134), .b(new_n133), .o1(new_n135));
  xobna2aa1n03x5               g040(.a(new_n128), .b(new_n132), .c(new_n135), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n126), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n137), .b(new_n128), .c(new_n132), .d(new_n135), .o1(new_n138));
  xorb03aa1n02x5               g043(.a(new_n138), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norp02aa1n12x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand02aa1d06x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nona23aa1d18x5               g046(.a(new_n141), .b(new_n127), .c(new_n126), .d(new_n140), .out0(new_n142));
  tech160nm_fiaoi012aa1n03p5x5 g047(.a(new_n140), .b(new_n126), .c(new_n141), .o1(new_n143));
  oai012aa1n12x5               g048(.a(new_n143), .b(new_n142), .c(new_n135), .o1(new_n144));
  oab012aa1n06x5               g049(.a(new_n144), .b(new_n132), .c(new_n142), .out0(new_n145));
  nor002aa1d32x5               g050(.a(\b[12] ), .b(\a[13] ), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  nand42aa1n08x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n145), .b(new_n148), .c(new_n147), .out0(\s[13] ));
  nanb02aa1n02x5               g054(.a(new_n146), .b(new_n148), .out0(new_n150));
  nor002aa1n16x5               g055(.a(\b[13] ), .b(\a[14] ), .o1(new_n151));
  nand42aa1n08x5               g056(.a(\b[13] ), .b(\a[14] ), .o1(new_n152));
  nanb02aa1n02x5               g057(.a(new_n151), .b(new_n152), .out0(new_n153));
  oai112aa1n03x5               g058(.a(new_n153), .b(new_n147), .c(new_n145), .d(new_n150), .o1(new_n154));
  oaoi13aa1n09x5               g059(.a(new_n153), .b(new_n147), .c(new_n145), .d(new_n150), .o1(new_n155));
  norb02aa1n03x4               g060(.a(new_n154), .b(new_n155), .out0(\s[14] ));
  inv040aa1n02x5               g061(.a(new_n142), .o1(new_n157));
  nano23aa1n09x5               g062(.a(new_n146), .b(new_n151), .c(new_n152), .d(new_n148), .out0(new_n158));
  nano32aa1n03x7               g063(.a(new_n123), .b(new_n158), .c(new_n131), .d(new_n157), .out0(new_n159));
  tech160nm_fioai012aa1n04x5   g064(.a(new_n152), .b(new_n151), .c(new_n146), .o1(new_n160));
  aob012aa1n02x5               g065(.a(new_n160), .b(new_n144), .c(new_n158), .out0(new_n161));
  norp02aa1n02x5               g066(.a(new_n159), .b(new_n161), .o1(new_n162));
  xorc02aa1n02x5               g067(.a(\a[15] ), .b(\b[14] ), .out0(new_n163));
  xnrc02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(\s[15] ));
  inv000aa1d42x5               g069(.a(\a[16] ), .o1(new_n165));
  norp02aa1n02x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  oaoi13aa1n03x5               g071(.a(new_n166), .b(new_n163), .c(new_n159), .d(new_n161), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[15] ), .c(new_n165), .out0(\s[16] ));
  nona23aa1n02x4               g073(.a(new_n152), .b(new_n148), .c(new_n146), .d(new_n151), .out0(new_n169));
  tech160nm_fixnrc02aa1n02p5x5 g074(.a(\b[14] ), .b(\a[15] ), .out0(new_n170));
  xnrc02aa1n06x5               g075(.a(\b[15] ), .b(\a[16] ), .out0(new_n171));
  nor042aa1n03x5               g076(.a(new_n171), .b(new_n170), .o1(new_n172));
  nona23aa1n06x5               g077(.a(new_n131), .b(new_n172), .c(new_n169), .d(new_n142), .out0(new_n173));
  aoi112aa1n02x5               g078(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n174));
  aoib12aa1n02x5               g079(.a(new_n174), .b(new_n165), .c(\b[15] ), .out0(new_n175));
  oai013aa1n02x5               g080(.a(new_n175), .b(new_n170), .c(new_n171), .d(new_n160), .o1(new_n176));
  aoi013aa1n09x5               g081(.a(new_n176), .b(new_n144), .c(new_n158), .d(new_n172), .o1(new_n177));
  oai012aa1n12x5               g082(.a(new_n177), .b(new_n123), .c(new_n173), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g084(.a(\a[18] ), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\a[17] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(\b[16] ), .o1(new_n182));
  oaoi03aa1n03x5               g087(.a(new_n181), .b(new_n182), .c(new_n178), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[17] ), .c(new_n180), .out0(\s[18] ));
  xorc02aa1n02x5               g089(.a(\a[16] ), .b(\b[15] ), .out0(new_n185));
  nand23aa1n03x5               g090(.a(new_n158), .b(new_n163), .c(new_n185), .o1(new_n186));
  nano22aa1n03x7               g091(.a(new_n186), .b(new_n131), .c(new_n157), .out0(new_n187));
  aoai13aa1n06x5               g092(.a(new_n187), .b(new_n122), .c(new_n107), .d(new_n117), .o1(new_n188));
  xroi22aa1d06x4               g093(.a(new_n181), .b(\b[16] ), .c(new_n180), .d(\b[17] ), .out0(new_n189));
  inv000aa1n02x5               g094(.a(new_n189), .o1(new_n190));
  oai022aa1d24x5               g095(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n191));
  oaib12aa1n18x5               g096(.a(new_n191), .b(new_n180), .c(\b[17] ), .out0(new_n192));
  aoai13aa1n02x7               g097(.a(new_n192), .b(new_n190), .c(new_n188), .d(new_n177), .o1(new_n193));
  xorb03aa1n02x5               g098(.a(new_n193), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  xorc02aa1n12x5               g101(.a(\a[19] ), .b(\b[18] ), .out0(new_n197));
  tech160nm_fixorc02aa1n05x5   g102(.a(\a[20] ), .b(\b[19] ), .out0(new_n198));
  aoi112aa1n03x4               g103(.a(new_n196), .b(new_n198), .c(new_n193), .d(new_n197), .o1(new_n199));
  inv000aa1n04x5               g104(.a(new_n196), .o1(new_n200));
  nor042aa1d18x5               g105(.a(\b[16] ), .b(\a[17] ), .o1(new_n201));
  inv020aa1n03x5               g106(.a(new_n201), .o1(new_n202));
  oaoi03aa1n02x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n197), .b(new_n203), .c(new_n178), .d(new_n189), .o1(new_n204));
  xnrc02aa1n12x5               g109(.a(\b[19] ), .b(\a[20] ), .out0(new_n205));
  tech160nm_fiaoi012aa1n02p5x5 g110(.a(new_n205), .b(new_n204), .c(new_n200), .o1(new_n206));
  nor002aa1n02x5               g111(.a(new_n206), .b(new_n199), .o1(\s[20] ));
  nand22aa1n03x5               g112(.a(new_n198), .b(new_n197), .o1(new_n208));
  norb02aa1n03x5               g113(.a(new_n189), .b(new_n208), .out0(new_n209));
  inv000aa1n02x5               g114(.a(new_n209), .o1(new_n210));
  xnrc02aa1n12x5               g115(.a(\b[18] ), .b(\a[19] ), .out0(new_n211));
  oao003aa1n09x5               g116(.a(\a[20] ), .b(\b[19] ), .c(new_n200), .carry(new_n212));
  oai013aa1d12x5               g117(.a(new_n212), .b(new_n211), .c(new_n205), .d(new_n192), .o1(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  aoai13aa1n04x5               g119(.a(new_n214), .b(new_n210), .c(new_n188), .d(new_n177), .o1(new_n215));
  xorb03aa1n02x5               g120(.a(new_n215), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  nand02aa1n04x5               g122(.a(\b[20] ), .b(\a[21] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  nor042aa1n04x5               g124(.a(\b[21] ), .b(\a[22] ), .o1(new_n220));
  nanp02aa1n04x5               g125(.a(\b[21] ), .b(\a[22] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  aoi112aa1n03x4               g127(.a(new_n217), .b(new_n222), .c(new_n215), .d(new_n219), .o1(new_n223));
  inv040aa1n03x5               g128(.a(new_n217), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n219), .b(new_n213), .c(new_n178), .d(new_n209), .o1(new_n225));
  inv000aa1d42x5               g130(.a(new_n222), .o1(new_n226));
  tech160nm_fiaoi012aa1n02p5x5 g131(.a(new_n226), .b(new_n225), .c(new_n224), .o1(new_n227));
  nor002aa1n02x5               g132(.a(new_n227), .b(new_n223), .o1(\s[22] ));
  nano23aa1d15x5               g133(.a(new_n217), .b(new_n220), .c(new_n221), .d(new_n218), .out0(new_n229));
  nano32aa1n03x7               g134(.a(new_n190), .b(new_n229), .c(new_n197), .d(new_n198), .out0(new_n230));
  inv000aa1n02x5               g135(.a(new_n230), .o1(new_n231));
  oaoi03aa1n09x5               g136(.a(\a[22] ), .b(\b[21] ), .c(new_n224), .o1(new_n232));
  aoi012aa1d18x5               g137(.a(new_n232), .b(new_n213), .c(new_n229), .o1(new_n233));
  aoai13aa1n04x5               g138(.a(new_n233), .b(new_n231), .c(new_n188), .d(new_n177), .o1(new_n234));
  xorb03aa1n02x5               g139(.a(new_n234), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n10x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  nand42aa1d28x5               g141(.a(\b[22] ), .b(\a[23] ), .o1(new_n237));
  norb02aa1n02x5               g142(.a(new_n237), .b(new_n236), .out0(new_n238));
  nor042aa1n04x5               g143(.a(\b[23] ), .b(\a[24] ), .o1(new_n239));
  nand42aa1n16x5               g144(.a(\b[23] ), .b(\a[24] ), .o1(new_n240));
  norb02aa1n02x5               g145(.a(new_n240), .b(new_n239), .out0(new_n241));
  aoi112aa1n03x4               g146(.a(new_n236), .b(new_n241), .c(new_n234), .d(new_n238), .o1(new_n242));
  inv030aa1n02x5               g147(.a(new_n236), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n233), .o1(new_n244));
  aoai13aa1n03x5               g149(.a(new_n238), .b(new_n244), .c(new_n178), .d(new_n230), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n241), .o1(new_n246));
  aoi012aa1n02x7               g151(.a(new_n246), .b(new_n245), .c(new_n243), .o1(new_n247));
  nor002aa1n02x5               g152(.a(new_n247), .b(new_n242), .o1(\s[24] ));
  nano23aa1d15x5               g153(.a(new_n236), .b(new_n239), .c(new_n240), .d(new_n237), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  nano23aa1n02x4               g155(.a(new_n250), .b(new_n208), .c(new_n189), .d(new_n229), .out0(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  nanp03aa1n02x5               g157(.a(new_n203), .b(new_n197), .c(new_n198), .o1(new_n253));
  nand02aa1d04x5               g158(.a(new_n249), .b(new_n229), .o1(new_n254));
  oaoi03aa1n03x5               g159(.a(\a[24] ), .b(\b[23] ), .c(new_n243), .o1(new_n255));
  aoi012aa1n12x5               g160(.a(new_n255), .b(new_n249), .c(new_n232), .o1(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n254), .c(new_n253), .d(new_n212), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n02x7               g163(.a(new_n258), .b(new_n252), .c(new_n188), .d(new_n177), .o1(new_n259));
  xorb03aa1n02x5               g164(.a(new_n259), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  tech160nm_fixorc02aa1n02p5x5 g166(.a(\a[25] ), .b(\b[24] ), .out0(new_n262));
  xorc02aa1n12x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  aoi112aa1n03x4               g168(.a(new_n261), .b(new_n263), .c(new_n259), .d(new_n262), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n261), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n262), .b(new_n257), .c(new_n178), .d(new_n251), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n263), .o1(new_n267));
  tech160nm_fiaoi012aa1n02p5x5 g172(.a(new_n267), .b(new_n266), .c(new_n265), .o1(new_n268));
  nor002aa1n02x5               g173(.a(new_n268), .b(new_n264), .o1(\s[26] ));
  and002aa1n06x5               g174(.a(new_n263), .b(new_n262), .o(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  nona22aa1n03x5               g176(.a(new_n230), .b(new_n250), .c(new_n271), .out0(new_n272));
  oao003aa1n02x5               g177(.a(\a[26] ), .b(\b[25] ), .c(new_n265), .carry(new_n273));
  aobi12aa1n06x5               g178(.a(new_n273), .b(new_n257), .c(new_n270), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n272), .c(new_n188), .d(new_n177), .o1(new_n275));
  xorb03aa1n03x5               g180(.a(new_n275), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n09x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  xorc02aa1n02x5               g182(.a(\a[27] ), .b(\b[26] ), .out0(new_n278));
  xorc02aa1n12x5               g183(.a(\a[28] ), .b(\b[27] ), .out0(new_n279));
  aoi112aa1n03x4               g184(.a(new_n277), .b(new_n279), .c(new_n275), .d(new_n278), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n277), .o1(new_n281));
  nano32aa1n02x5               g186(.a(new_n210), .b(new_n270), .c(new_n229), .d(new_n249), .out0(new_n282));
  inv030aa1n02x5               g187(.a(new_n254), .o1(new_n283));
  nanp02aa1n03x5               g188(.a(new_n283), .b(new_n213), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n273), .b(new_n271), .c(new_n284), .d(new_n256), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n278), .b(new_n285), .c(new_n178), .d(new_n282), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n279), .o1(new_n287));
  tech160nm_fiaoi012aa1n02p5x5 g192(.a(new_n287), .b(new_n286), .c(new_n281), .o1(new_n288));
  nor002aa1n02x5               g193(.a(new_n288), .b(new_n280), .o1(\s[28] ));
  and002aa1n02x5               g194(.a(new_n279), .b(new_n278), .o(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n178), .d(new_n282), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\a[28] ), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\b[27] ), .o1(new_n293));
  oaoi03aa1n09x5               g198(.a(new_n292), .b(new_n293), .c(new_n277), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[29] ), .b(\b[28] ), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  aoi012aa1n03x5               g201(.a(new_n296), .b(new_n291), .c(new_n294), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n294), .o1(new_n298));
  aoi112aa1n03x4               g203(.a(new_n295), .b(new_n298), .c(new_n275), .d(new_n290), .o1(new_n299));
  norp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g206(.a(new_n296), .b(new_n278), .c(new_n279), .out0(new_n302));
  aoai13aa1n03x5               g207(.a(new_n302), .b(new_n285), .c(new_n178), .d(new_n282), .o1(new_n303));
  tech160nm_fioaoi03aa1n03p5x5 g208(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .o1(new_n304));
  inv000aa1n02x5               g209(.a(new_n304), .o1(new_n305));
  xorc02aa1n12x5               g210(.a(\a[30] ), .b(\b[29] ), .out0(new_n306));
  inv000aa1d42x5               g211(.a(new_n306), .o1(new_n307));
  tech160nm_fiaoi012aa1n02p5x5 g212(.a(new_n307), .b(new_n303), .c(new_n305), .o1(new_n308));
  aoi112aa1n03x4               g213(.a(new_n306), .b(new_n304), .c(new_n275), .d(new_n302), .o1(new_n309));
  nor002aa1n02x5               g214(.a(new_n308), .b(new_n309), .o1(\s[30] ));
  nano32aa1n02x4               g215(.a(new_n307), .b(new_n295), .c(new_n279), .d(new_n278), .out0(new_n311));
  oaoi03aa1n02x5               g216(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[31] ), .b(\b[30] ), .out0(new_n313));
  aoi112aa1n03x4               g218(.a(new_n313), .b(new_n312), .c(new_n275), .d(new_n311), .o1(new_n314));
  aoai13aa1n03x5               g219(.a(new_n311), .b(new_n285), .c(new_n178), .d(new_n282), .o1(new_n315));
  inv000aa1n02x5               g220(.a(new_n312), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n313), .o1(new_n317));
  tech160nm_fiaoi012aa1n03p5x5 g222(.a(new_n317), .b(new_n315), .c(new_n316), .o1(new_n318));
  nor042aa1n03x5               g223(.a(new_n318), .b(new_n314), .o1(\s[31] ));
  xnrb03aa1n02x5               g224(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g225(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oao003aa1n02x5               g228(.a(new_n118), .b(new_n119), .c(new_n107), .carry(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g230(.a(new_n111), .b(new_n110), .out0(new_n326));
  aoai13aa1n02x5               g231(.a(new_n326), .b(new_n113), .c(new_n324), .d(new_n114), .o1(new_n327));
  aoi112aa1n02x5               g232(.a(new_n326), .b(new_n113), .c(new_n324), .d(new_n114), .o1(new_n328));
  norb02aa1n02x5               g233(.a(new_n327), .b(new_n328), .out0(\s[7] ));
  norb02aa1n02x5               g234(.a(new_n109), .b(new_n108), .out0(new_n330));
  inv000aa1d42x5               g235(.a(new_n110), .o1(new_n331));
  xnbna2aa1n03x5               g236(.a(new_n330), .b(new_n327), .c(new_n331), .out0(\s[8] ));
  xorb03aa1n02x5               g237(.a(new_n123), .b(new_n130), .c(\a[9] ), .out0(\s[9] ));
endmodule


