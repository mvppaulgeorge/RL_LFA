// Benchmark "adder" written by ABC on Thu Jul 18 07:46:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n344, new_n347,
    new_n349, new_n350, new_n352, new_n353, new_n354, new_n355, new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  aoi012aa1n02x5               g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  nand02aa1n06x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  norp02aa1n06x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor042aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n03x5               g009(.a(new_n101), .b(new_n104), .c(new_n103), .d(new_n102), .out0(new_n105));
  aoi012aa1n12x5               g010(.a(new_n102), .b(new_n103), .c(new_n101), .o1(new_n106));
  tech160nm_fioai012aa1n03p5x5 g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  nand42aa1n03x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nanb02aa1n02x5               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  inv000aa1d42x5               g016(.a(\a[5] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[4] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(new_n113), .b(new_n112), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(new_n114), .b(new_n111), .o1(new_n115));
  nor002aa1n04x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand42aa1n02x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nor042aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nona23aa1n02x4               g024(.a(new_n118), .b(new_n117), .c(new_n119), .d(new_n116), .out0(new_n120));
  nor043aa1n02x5               g025(.a(new_n120), .b(new_n115), .c(new_n110), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\a[7] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[6] ), .o1(new_n123));
  aoai13aa1n02x5               g028(.a(new_n117), .b(new_n116), .c(new_n122), .d(new_n123), .o1(new_n124));
  aoai13aa1n02x5               g029(.a(new_n108), .b(new_n109), .c(new_n113), .d(new_n112), .o1(new_n125));
  oai012aa1n02x5               g030(.a(new_n124), .b(new_n120), .c(new_n125), .o1(new_n126));
  nor002aa1n02x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nand42aa1n03x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n126), .c(new_n107), .d(new_n121), .o1(new_n130));
  oai012aa1n02x5               g035(.a(new_n130), .b(\b[8] ), .c(\a[9] ), .o1(new_n131));
  xorb03aa1n02x5               g036(.a(new_n131), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  inv000aa1d42x5               g037(.a(\b[9] ), .o1(new_n133));
  nanb02aa1n02x5               g038(.a(\a[10] ), .b(new_n133), .out0(new_n134));
  nand42aa1n04x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  inv000aa1n02x5               g040(.a(new_n97), .o1(new_n136));
  aob012aa1n02x5               g041(.a(new_n136), .b(new_n98), .c(new_n99), .out0(new_n137));
  norb02aa1n02x5               g042(.a(new_n101), .b(new_n102), .out0(new_n138));
  norb02aa1n02x7               g043(.a(new_n104), .b(new_n103), .out0(new_n139));
  nanp03aa1n02x5               g044(.a(new_n137), .b(new_n138), .c(new_n139), .o1(new_n140));
  nano23aa1n03x7               g045(.a(new_n119), .b(new_n116), .c(new_n117), .d(new_n118), .out0(new_n141));
  nona22aa1n02x4               g046(.a(new_n141), .b(new_n110), .c(new_n115), .out0(new_n142));
  oaoi03aa1n02x5               g047(.a(\a[6] ), .b(\b[5] ), .c(new_n114), .o1(new_n143));
  aobi12aa1n06x5               g048(.a(new_n124), .b(new_n141), .c(new_n143), .out0(new_n144));
  aoai13aa1n12x5               g049(.a(new_n144), .b(new_n142), .c(new_n140), .d(new_n106), .o1(new_n145));
  aoai13aa1n06x5               g050(.a(new_n135), .b(new_n127), .c(new_n145), .d(new_n129), .o1(new_n146));
  nand42aa1n02x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  nor022aa1n16x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nanb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n146), .c(new_n134), .out0(\s[11] ));
  norp02aa1n02x5               g056(.a(\b[9] ), .b(\a[10] ), .o1(new_n152));
  aoai13aa1n02x5               g057(.a(new_n150), .b(new_n152), .c(new_n131), .d(new_n135), .o1(new_n153));
  nor002aa1n06x5               g058(.a(\b[11] ), .b(\a[12] ), .o1(new_n154));
  nand42aa1d28x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  inv000aa1n02x5               g061(.a(new_n148), .o1(new_n157));
  oaib12aa1n18x5               g062(.a(new_n157), .b(new_n154), .c(new_n155), .out0(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n02x5               g064(.a(new_n157), .b(new_n149), .c(new_n146), .d(new_n134), .o1(new_n160));
  aoi022aa1n02x5               g065(.a(new_n160), .b(new_n156), .c(new_n153), .d(new_n159), .o1(\s[12] ));
  norb03aa1n03x5               g066(.a(new_n128), .b(new_n152), .c(new_n127), .out0(new_n162));
  nano22aa1n03x7               g067(.a(new_n148), .b(new_n135), .c(new_n147), .out0(new_n163));
  nanp03aa1d12x5               g068(.a(new_n158), .b(new_n163), .c(new_n162), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n126), .c(new_n107), .d(new_n121), .o1(new_n166));
  oai012aa1n02x5               g071(.a(new_n155), .b(new_n154), .c(new_n148), .o1(new_n167));
  oai112aa1n02x5               g072(.a(new_n134), .b(new_n135), .c(\b[8] ), .d(\a[9] ), .o1(new_n168));
  nand23aa1n04x5               g073(.a(new_n158), .b(new_n163), .c(new_n168), .o1(new_n169));
  nand22aa1n06x5               g074(.a(new_n169), .b(new_n167), .o1(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  nand42aa1n03x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  nor022aa1n16x5               g077(.a(\b[12] ), .b(\a[13] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n166), .c(new_n171), .out0(\s[13] ));
  inv000aa1d42x5               g080(.a(new_n173), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n174), .b(new_n170), .c(new_n145), .d(new_n165), .o1(new_n177));
  nor002aa1n02x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  nand42aa1n03x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n177), .c(new_n176), .out0(\s[14] ));
  nona23aa1n02x4               g086(.a(new_n172), .b(new_n179), .c(new_n178), .d(new_n173), .out0(new_n182));
  oai012aa1n02x5               g087(.a(new_n179), .b(new_n178), .c(new_n173), .o1(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n182), .c(new_n166), .d(new_n171), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  xorc02aa1n12x5               g090(.a(\a[15] ), .b(\b[14] ), .out0(new_n186));
  nanp02aa1n02x5               g091(.a(new_n184), .b(new_n186), .o1(new_n187));
  xorc02aa1n02x5               g092(.a(\a[16] ), .b(\b[15] ), .out0(new_n188));
  nor042aa1n03x5               g093(.a(\b[14] ), .b(\a[15] ), .o1(new_n189));
  norp02aa1n02x5               g094(.a(new_n188), .b(new_n189), .o1(new_n190));
  nano23aa1n03x5               g095(.a(new_n178), .b(new_n173), .c(new_n179), .d(new_n172), .out0(new_n191));
  aoai13aa1n02x5               g096(.a(new_n191), .b(new_n170), .c(new_n145), .d(new_n165), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n189), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n186), .o1(new_n194));
  aoai13aa1n02x5               g099(.a(new_n193), .b(new_n194), .c(new_n192), .d(new_n183), .o1(new_n195));
  aoi022aa1n02x5               g100(.a(new_n195), .b(new_n188), .c(new_n187), .d(new_n190), .o1(\s[16] ));
  nand23aa1n03x5               g101(.a(new_n191), .b(new_n186), .c(new_n188), .o1(new_n197));
  nor042aa1n12x5               g102(.a(new_n197), .b(new_n164), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n126), .c(new_n107), .d(new_n121), .o1(new_n199));
  xnrc02aa1n02x5               g104(.a(\b[15] ), .b(\a[16] ), .out0(new_n200));
  norb03aa1n02x5               g105(.a(new_n186), .b(new_n182), .c(new_n200), .out0(new_n201));
  oaoi03aa1n02x5               g106(.a(\a[16] ), .b(\b[15] ), .c(new_n193), .o1(new_n202));
  oaoi03aa1n02x5               g107(.a(\a[14] ), .b(\b[13] ), .c(new_n176), .o1(new_n203));
  nanp03aa1n02x5               g108(.a(new_n203), .b(new_n186), .c(new_n188), .o1(new_n204));
  nanb02aa1n02x5               g109(.a(new_n202), .b(new_n204), .out0(new_n205));
  aoi012aa1n09x5               g110(.a(new_n205), .b(new_n170), .c(new_n201), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[17] ), .b(\b[16] ), .out0(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n199), .c(new_n206), .out0(\s[17] ));
  inv000aa1d42x5               g113(.a(\a[17] ), .o1(new_n209));
  inv000aa1d42x5               g114(.a(\b[16] ), .o1(new_n210));
  nanp02aa1n02x5               g115(.a(new_n210), .b(new_n209), .o1(new_n211));
  aoi013aa1n02x4               g116(.a(new_n202), .b(new_n203), .c(new_n186), .d(new_n188), .o1(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n197), .c(new_n167), .d(new_n169), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n207), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n214));
  xorc02aa1n02x5               g119(.a(\a[18] ), .b(\b[17] ), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n214), .c(new_n211), .out0(\s[18] ));
  inv000aa1d42x5               g121(.a(\a[18] ), .o1(new_n217));
  xroi22aa1d06x4               g122(.a(new_n209), .b(\b[16] ), .c(new_n217), .d(\b[17] ), .out0(new_n218));
  aoai13aa1n04x5               g123(.a(new_n218), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n219));
  oaih22aa1d12x5               g124(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n220));
  oaib12aa1n06x5               g125(.a(new_n220), .b(new_n217), .c(\b[17] ), .out0(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[18] ), .b(\a[19] ), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n219), .c(new_n221), .out0(\s[19] ));
  xnrc02aa1n02x5               g129(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n09x5               g130(.a(new_n199), .b(new_n206), .o1(new_n226));
  oaoi03aa1n02x5               g131(.a(\a[18] ), .b(\b[17] ), .c(new_n211), .o1(new_n227));
  aoai13aa1n03x5               g132(.a(new_n223), .b(new_n227), .c(new_n226), .d(new_n218), .o1(new_n228));
  xorc02aa1n02x5               g133(.a(\a[20] ), .b(\b[19] ), .out0(new_n229));
  nor042aa1n03x5               g134(.a(\b[18] ), .b(\a[19] ), .o1(new_n230));
  norp02aa1n02x5               g135(.a(new_n229), .b(new_n230), .o1(new_n231));
  inv000aa1n02x5               g136(.a(new_n230), .o1(new_n232));
  aoai13aa1n02x5               g137(.a(new_n232), .b(new_n222), .c(new_n219), .d(new_n221), .o1(new_n233));
  aoi022aa1n03x5               g138(.a(new_n233), .b(new_n229), .c(new_n228), .d(new_n231), .o1(\s[20] ));
  tech160nm_fixnrc02aa1n04x5   g139(.a(\b[19] ), .b(\a[20] ), .out0(new_n235));
  nona22aa1n09x5               g140(.a(new_n218), .b(new_n222), .c(new_n235), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n238));
  oao003aa1n02x5               g143(.a(\a[20] ), .b(\b[19] ), .c(new_n232), .carry(new_n239));
  oai013aa1d12x5               g144(.a(new_n239), .b(new_n222), .c(new_n235), .d(new_n221), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  nand42aa1n02x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  nor042aa1n06x5               g147(.a(\b[20] ), .b(\a[21] ), .o1(new_n243));
  norb02aa1n02x5               g148(.a(new_n242), .b(new_n243), .out0(new_n244));
  xnbna2aa1n03x5               g149(.a(new_n244), .b(new_n238), .c(new_n241), .out0(\s[21] ));
  aoai13aa1n06x5               g150(.a(new_n244), .b(new_n240), .c(new_n226), .d(new_n237), .o1(new_n246));
  nor042aa1n02x5               g151(.a(\b[21] ), .b(\a[22] ), .o1(new_n247));
  nand42aa1n03x5               g152(.a(\b[21] ), .b(\a[22] ), .o1(new_n248));
  norb02aa1n02x5               g153(.a(new_n248), .b(new_n247), .out0(new_n249));
  inv000aa1d42x5               g154(.a(\a[21] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[20] ), .o1(new_n251));
  aboi22aa1n03x5               g156(.a(new_n247), .b(new_n248), .c(new_n250), .d(new_n251), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n243), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n244), .o1(new_n254));
  aoai13aa1n02x5               g159(.a(new_n253), .b(new_n254), .c(new_n238), .d(new_n241), .o1(new_n255));
  aoi022aa1n03x5               g160(.a(new_n255), .b(new_n249), .c(new_n246), .d(new_n252), .o1(\s[22] ));
  nano23aa1d15x5               g161(.a(new_n247), .b(new_n243), .c(new_n248), .d(new_n242), .out0(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  norp02aa1n02x5               g163(.a(new_n236), .b(new_n258), .o1(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n260));
  tech160nm_fioaoi03aa1n03p5x5 g165(.a(\a[22] ), .b(\b[21] ), .c(new_n253), .o1(new_n261));
  aoi012aa1d18x5               g166(.a(new_n261), .b(new_n240), .c(new_n257), .o1(new_n262));
  nor042aa1n04x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  nanb02aa1n02x5               g169(.a(new_n263), .b(new_n264), .out0(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n260), .c(new_n262), .out0(\s[23] ));
  inv000aa1d42x5               g172(.a(new_n262), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n266), .b(new_n268), .c(new_n226), .d(new_n259), .o1(new_n269));
  norp02aa1n02x5               g174(.a(\b[23] ), .b(\a[24] ), .o1(new_n270));
  nanp02aa1n02x5               g175(.a(\b[23] ), .b(\a[24] ), .o1(new_n271));
  norb02aa1n02x5               g176(.a(new_n271), .b(new_n270), .out0(new_n272));
  aoib12aa1n02x5               g177(.a(new_n263), .b(new_n271), .c(new_n270), .out0(new_n273));
  inv000aa1d42x5               g178(.a(new_n263), .o1(new_n274));
  aoai13aa1n02x5               g179(.a(new_n274), .b(new_n265), .c(new_n260), .d(new_n262), .o1(new_n275));
  aoi022aa1n03x5               g180(.a(new_n275), .b(new_n272), .c(new_n269), .d(new_n273), .o1(\s[24] ));
  nano23aa1n06x5               g181(.a(new_n263), .b(new_n270), .c(new_n271), .d(new_n264), .out0(new_n277));
  nand22aa1n03x5               g182(.a(new_n277), .b(new_n257), .o1(new_n278));
  nor002aa1n02x5               g183(.a(new_n236), .b(new_n278), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n279), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n280));
  nanb03aa1n02x5               g185(.a(new_n222), .b(new_n227), .c(new_n229), .out0(new_n281));
  aoi012aa1n02x5               g186(.a(new_n270), .b(new_n263), .c(new_n271), .o1(new_n282));
  aobi12aa1n06x5               g187(.a(new_n282), .b(new_n277), .c(new_n261), .out0(new_n283));
  aoai13aa1n06x5               g188(.a(new_n283), .b(new_n278), .c(new_n281), .d(new_n239), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n284), .c(new_n226), .d(new_n279), .o1(new_n286));
  inv000aa1n02x5               g191(.a(new_n283), .o1(new_n287));
  aoi113aa1n02x5               g192(.a(new_n287), .b(new_n285), .c(new_n240), .d(new_n257), .e(new_n277), .o1(new_n288));
  aobi12aa1n03x7               g193(.a(new_n286), .b(new_n288), .c(new_n280), .out0(\s[25] ));
  xorc02aa1n02x5               g194(.a(\a[26] ), .b(\b[25] ), .out0(new_n290));
  nor042aa1n03x5               g195(.a(\b[24] ), .b(\a[25] ), .o1(new_n291));
  norp02aa1n02x5               g196(.a(new_n290), .b(new_n291), .o1(new_n292));
  aoib12aa1n06x5               g197(.a(new_n287), .b(new_n240), .c(new_n278), .out0(new_n293));
  inv000aa1d42x5               g198(.a(new_n291), .o1(new_n294));
  inv000aa1d42x5               g199(.a(new_n285), .o1(new_n295));
  aoai13aa1n02x7               g200(.a(new_n294), .b(new_n295), .c(new_n280), .d(new_n293), .o1(new_n296));
  aoi022aa1n02x7               g201(.a(new_n296), .b(new_n290), .c(new_n286), .d(new_n292), .o1(\s[26] ));
  and002aa1n12x5               g202(.a(new_n290), .b(new_n285), .o(new_n298));
  nano32aa1n03x7               g203(.a(new_n236), .b(new_n298), .c(new_n257), .d(new_n277), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n213), .c(new_n145), .d(new_n198), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[26] ), .b(\b[25] ), .c(new_n294), .carry(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  tech160nm_fiaoi012aa1n05x5   g207(.a(new_n302), .b(new_n284), .c(new_n298), .o1(new_n303));
  xorc02aa1n12x5               g208(.a(\a[27] ), .b(\b[26] ), .out0(new_n304));
  xnbna2aa1n03x5               g209(.a(new_n304), .b(new_n300), .c(new_n303), .out0(\s[27] ));
  inv000aa1d42x5               g210(.a(new_n298), .o1(new_n306));
  oai012aa1n06x5               g211(.a(new_n301), .b(new_n293), .c(new_n306), .o1(new_n307));
  aoai13aa1n03x5               g212(.a(new_n304), .b(new_n307), .c(new_n226), .d(new_n299), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[28] ), .b(\b[27] ), .out0(new_n309));
  norp02aa1n02x5               g214(.a(\b[26] ), .b(\a[27] ), .o1(new_n310));
  norp02aa1n02x5               g215(.a(new_n309), .b(new_n310), .o1(new_n311));
  inv000aa1n03x5               g216(.a(new_n310), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n304), .o1(new_n313));
  aoai13aa1n02x5               g218(.a(new_n312), .b(new_n313), .c(new_n300), .d(new_n303), .o1(new_n314));
  aoi022aa1n03x5               g219(.a(new_n314), .b(new_n309), .c(new_n308), .d(new_n311), .o1(\s[28] ));
  and002aa1n02x5               g220(.a(new_n309), .b(new_n304), .o(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n307), .c(new_n226), .d(new_n299), .o1(new_n317));
  inv000aa1d42x5               g222(.a(new_n316), .o1(new_n318));
  oao003aa1n02x5               g223(.a(\a[28] ), .b(\b[27] ), .c(new_n312), .carry(new_n319));
  aoai13aa1n02x5               g224(.a(new_n319), .b(new_n318), .c(new_n300), .d(new_n303), .o1(new_n320));
  xorc02aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .out0(new_n321));
  norb02aa1n02x5               g226(.a(new_n319), .b(new_n321), .out0(new_n322));
  aoi022aa1n03x5               g227(.a(new_n320), .b(new_n321), .c(new_n317), .d(new_n322), .o1(\s[29] ));
  xorb03aa1n02x5               g228(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g229(.a(new_n313), .b(new_n309), .c(new_n321), .out0(new_n325));
  aoai13aa1n02x5               g230(.a(new_n325), .b(new_n307), .c(new_n226), .d(new_n299), .o1(new_n326));
  inv000aa1d42x5               g231(.a(new_n325), .o1(new_n327));
  oao003aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .c(new_n319), .carry(new_n328));
  aoai13aa1n02x5               g233(.a(new_n328), .b(new_n327), .c(new_n300), .d(new_n303), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .out0(new_n330));
  norb02aa1n02x5               g235(.a(new_n328), .b(new_n330), .out0(new_n331));
  aoi022aa1n03x5               g236(.a(new_n329), .b(new_n330), .c(new_n326), .d(new_n331), .o1(\s[30] ));
  nano32aa1d15x5               g237(.a(new_n313), .b(new_n330), .c(new_n309), .d(new_n321), .out0(new_n333));
  aoai13aa1n03x5               g238(.a(new_n333), .b(new_n307), .c(new_n226), .d(new_n299), .o1(new_n334));
  xorc02aa1n02x5               g239(.a(\a[31] ), .b(\b[30] ), .out0(new_n335));
  and002aa1n02x5               g240(.a(\b[29] ), .b(\a[30] ), .o(new_n336));
  oabi12aa1n02x5               g241(.a(new_n335), .b(\a[30] ), .c(\b[29] ), .out0(new_n337));
  oab012aa1n02x4               g242(.a(new_n337), .b(new_n328), .c(new_n336), .out0(new_n338));
  inv000aa1d42x5               g243(.a(new_n333), .o1(new_n339));
  oao003aa1n02x5               g244(.a(\a[30] ), .b(\b[29] ), .c(new_n328), .carry(new_n340));
  aoai13aa1n02x5               g245(.a(new_n340), .b(new_n339), .c(new_n300), .d(new_n303), .o1(new_n341));
  aoi022aa1n03x5               g246(.a(new_n341), .b(new_n335), .c(new_n334), .d(new_n338), .o1(\s[31] ));
  xnrb03aa1n02x5               g247(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi112aa1n02x5               g248(.a(new_n103), .b(new_n138), .c(new_n137), .d(new_n104), .o1(new_n344));
  aoib12aa1n02x5               g249(.a(new_n344), .b(new_n107), .c(new_n102), .out0(\s[4] ));
  xorb03aa1n02x5               g250(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n02x5               g251(.a(new_n114), .b(new_n115), .c(new_n140), .d(new_n106), .o1(new_n347));
  xorb03aa1n02x5               g252(.a(new_n347), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g253(.a(new_n118), .b(new_n119), .out0(new_n349));
  nanb02aa1n02x5               g254(.a(new_n110), .b(new_n347), .out0(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n349), .b(new_n350), .c(new_n125), .out0(\s[7] ));
  norb02aa1n02x5               g256(.a(new_n117), .b(new_n116), .out0(new_n352));
  aob012aa1n02x5               g257(.a(new_n349), .b(new_n350), .c(new_n125), .out0(new_n353));
  aoib12aa1n02x5               g258(.a(new_n143), .b(new_n347), .c(new_n110), .out0(new_n354));
  oaoi03aa1n02x5               g259(.a(\a[7] ), .b(\b[6] ), .c(new_n354), .o1(new_n355));
  aboi22aa1n03x5               g260(.a(new_n116), .b(new_n117), .c(new_n122), .d(new_n123), .out0(new_n356));
  aoi022aa1n02x5               g261(.a(new_n355), .b(new_n352), .c(new_n353), .d(new_n356), .o1(\s[8] ));
  xorb03aa1n02x5               g262(.a(new_n145), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


