// Benchmark "adder" written by ABC on Thu Jul 18 11:52:31 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n335, new_n337, new_n338,
    new_n339, new_n341, new_n342, new_n343, new_n344, new_n345, new_n347,
    new_n348, new_n350, new_n351, new_n353, new_n354;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  oaih22aa1n04x5               g003(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n99));
  xnrc02aa1n12x5               g004(.a(\b[2] ), .b(\a[3] ), .out0(new_n100));
  tech160nm_finand02aa1n03p5x5 g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand02aa1d16x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  nor042aa1n06x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oaih12aa1n06x5               g008(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n104));
  oabi12aa1n18x5               g009(.a(new_n99), .b(new_n100), .c(new_n104), .out0(new_n105));
  nand42aa1n02x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nor002aa1d32x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  aoi012aa1n06x5               g012(.a(new_n107), .b(\a[5] ), .c(\b[4] ), .o1(new_n108));
  nor002aa1d24x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  aoi012aa1n06x5               g014(.a(new_n109), .b(\a[4] ), .c(\b[3] ), .o1(new_n110));
  nand22aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  norp02aa1n24x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nanp02aa1n12x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n113), .b(new_n111), .c(new_n114), .d(new_n112), .out0(new_n115));
  nano32aa1n03x7               g020(.a(new_n115), .b(new_n110), .c(new_n108), .d(new_n106), .out0(new_n116));
  inv000aa1d42x5               g021(.a(new_n107), .o1(new_n117));
  inv000aa1d42x5               g022(.a(new_n109), .o1(new_n118));
  oai012aa1n12x5               g023(.a(new_n113), .b(new_n114), .c(new_n112), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n111), .b(new_n106), .o1(new_n120));
  aoai13aa1n09x5               g025(.a(new_n117), .b(new_n120), .c(new_n119), .d(new_n118), .o1(new_n121));
  xnrc02aa1n12x5               g026(.a(\b[8] ), .b(\a[9] ), .out0(new_n122));
  inv000aa1d42x5               g027(.a(new_n122), .o1(new_n123));
  aoai13aa1n06x5               g028(.a(new_n123), .b(new_n121), .c(new_n116), .d(new_n105), .o1(new_n124));
  nor002aa1d32x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nand02aa1d20x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nanb02aa1n12x5               g031(.a(new_n125), .b(new_n126), .out0(new_n127));
  inv000aa1d42x5               g032(.a(new_n127), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n124), .c(new_n98), .out0(\s[10] ));
  nand22aa1n03x5               g034(.a(new_n124), .b(new_n98), .o1(new_n130));
  oaoi03aa1n02x5               g035(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n131));
  nor042aa1n09x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nand02aa1n08x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n133), .b(new_n132), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n134), .b(new_n131), .c(new_n130), .d(new_n128), .o1(new_n135));
  aoi112aa1n02x5               g040(.a(new_n134), .b(new_n131), .c(new_n130), .d(new_n128), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(\s[11] ));
  nor002aa1d32x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand02aa1d28x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  inv000aa1d42x5               g045(.a(new_n138), .o1(new_n141));
  aoi012aa1n02x5               g046(.a(new_n132), .b(new_n141), .c(new_n139), .o1(new_n142));
  tech160nm_fioai012aa1n03p5x5 g047(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .o1(new_n143));
  aoi022aa1n02x5               g048(.a(new_n143), .b(new_n140), .c(new_n135), .d(new_n142), .o1(\s[12] ));
  nona23aa1n09x5               g049(.a(new_n139), .b(new_n133), .c(new_n132), .d(new_n138), .out0(new_n145));
  nor043aa1n06x5               g050(.a(new_n145), .b(new_n127), .c(new_n122), .o1(new_n146));
  aoai13aa1n06x5               g051(.a(new_n146), .b(new_n121), .c(new_n116), .d(new_n105), .o1(new_n147));
  nanb03aa1n12x5               g052(.a(new_n138), .b(new_n139), .c(new_n133), .out0(new_n148));
  oai122aa1n12x5               g053(.a(new_n126), .b(new_n125), .c(new_n97), .d(\b[10] ), .e(\a[11] ), .o1(new_n149));
  aoi012aa1d18x5               g054(.a(new_n138), .b(new_n132), .c(new_n139), .o1(new_n150));
  oai012aa1d24x5               g055(.a(new_n150), .b(new_n149), .c(new_n148), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand42aa1n08x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  xnbna2aa1n03x5               g060(.a(new_n155), .b(new_n147), .c(new_n152), .out0(\s[13] ));
  inv000aa1n06x5               g061(.a(new_n153), .o1(new_n157));
  nanp02aa1n02x5               g062(.a(new_n147), .b(new_n152), .o1(new_n158));
  nanp02aa1n02x5               g063(.a(new_n158), .b(new_n155), .o1(new_n159));
  nor002aa1n04x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n08x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n159), .c(new_n157), .out0(\s[14] ));
  nano23aa1d15x5               g068(.a(new_n153), .b(new_n160), .c(new_n161), .d(new_n154), .out0(new_n164));
  oaoi03aa1n09x5               g069(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n165));
  norp02aa1n24x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nanp02aa1n04x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanb02aa1n02x5               g072(.a(new_n166), .b(new_n167), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n165), .c(new_n158), .d(new_n164), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n169), .b(new_n165), .c(new_n158), .d(new_n164), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(\s[15] ));
  nor002aa1d32x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand02aa1n06x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  aoib12aa1n02x5               g080(.a(new_n166), .b(new_n174), .c(new_n173), .out0(new_n176));
  tech160nm_fioai012aa1n03p5x5 g081(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .o1(new_n177));
  aboi22aa1n03x5               g082(.a(new_n175), .b(new_n177), .c(new_n170), .d(new_n176), .out0(\s[16] ));
  nanp02aa1n04x5               g083(.a(new_n116), .b(new_n105), .o1(new_n179));
  inv040aa1n03x5               g084(.a(new_n121), .o1(new_n180));
  nona23aa1n02x4               g085(.a(new_n161), .b(new_n154), .c(new_n153), .d(new_n160), .out0(new_n181));
  nona23aa1d16x5               g086(.a(new_n174), .b(new_n167), .c(new_n166), .d(new_n173), .out0(new_n182));
  nona22aa1n09x5               g087(.a(new_n146), .b(new_n181), .c(new_n182), .out0(new_n183));
  aoi012aa1d18x5               g088(.a(new_n183), .b(new_n179), .c(new_n180), .o1(new_n184));
  inv000aa1n02x5               g089(.a(new_n165), .o1(new_n185));
  nano22aa1n03x7               g090(.a(new_n138), .b(new_n133), .c(new_n139), .out0(new_n186));
  oai012aa1n02x7               g091(.a(new_n126), .b(\b[10] ), .c(\a[11] ), .o1(new_n187));
  oab012aa1n04x5               g092(.a(new_n187), .b(new_n97), .c(new_n125), .out0(new_n188));
  inv000aa1n02x5               g093(.a(new_n150), .o1(new_n189));
  aoai13aa1n12x5               g094(.a(new_n164), .b(new_n189), .c(new_n188), .d(new_n186), .o1(new_n190));
  tech160nm_fiaoi012aa1n03p5x5 g095(.a(new_n173), .b(new_n166), .c(new_n174), .o1(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n182), .c(new_n190), .d(new_n185), .o1(new_n192));
  nor042aa1d18x5               g097(.a(\b[16] ), .b(\a[17] ), .o1(new_n193));
  nand42aa1n03x5               g098(.a(\b[16] ), .b(\a[17] ), .o1(new_n194));
  norb02aa1n06x4               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  tech160nm_fioai012aa1n03p5x5 g100(.a(new_n195), .b(new_n192), .c(new_n184), .o1(new_n196));
  inv000aa1d42x5               g101(.a(new_n182), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n165), .c(new_n151), .d(new_n164), .o1(new_n198));
  nano23aa1n02x4               g103(.a(new_n195), .b(new_n184), .c(new_n198), .d(new_n191), .out0(new_n199));
  norb02aa1n02x5               g104(.a(new_n196), .b(new_n199), .out0(\s[17] ));
  inv000aa1n06x5               g105(.a(new_n193), .o1(new_n201));
  nor042aa1d18x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand42aa1n10x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norb02aa1n06x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n196), .c(new_n201), .out0(\s[18] ));
  nano23aa1n02x4               g110(.a(new_n193), .b(new_n202), .c(new_n203), .d(new_n194), .out0(new_n206));
  tech160nm_fioai012aa1n03p5x5 g111(.a(new_n206), .b(new_n192), .c(new_n184), .o1(new_n207));
  oaoi03aa1n02x5               g112(.a(\a[18] ), .b(\b[17] ), .c(new_n201), .o1(new_n208));
  inv000aa1n02x5               g113(.a(new_n208), .o1(new_n209));
  nor002aa1d24x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nand02aa1d16x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  norb02aa1n06x4               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  xnbna2aa1n03x5               g117(.a(new_n212), .b(new_n207), .c(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g118(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoi012aa1n06x5               g119(.a(new_n121), .b(new_n116), .c(new_n105), .o1(new_n215));
  oai112aa1n06x5               g120(.a(new_n198), .b(new_n191), .c(new_n215), .d(new_n183), .o1(new_n216));
  aoai13aa1n03x5               g121(.a(new_n212), .b(new_n208), .c(new_n216), .d(new_n206), .o1(new_n217));
  nor002aa1d32x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  nand02aa1d28x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  norb02aa1n03x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  inv000aa1d42x5               g125(.a(\a[19] ), .o1(new_n221));
  inv000aa1d42x5               g126(.a(\b[18] ), .o1(new_n222));
  aboi22aa1n03x5               g127(.a(new_n218), .b(new_n219), .c(new_n221), .d(new_n222), .out0(new_n223));
  inv040aa1n03x5               g128(.a(new_n210), .o1(new_n224));
  inv000aa1n03x5               g129(.a(new_n212), .o1(new_n225));
  aoai13aa1n02x7               g130(.a(new_n224), .b(new_n225), .c(new_n207), .d(new_n209), .o1(new_n226));
  aoi022aa1n03x5               g131(.a(new_n226), .b(new_n220), .c(new_n217), .d(new_n223), .o1(\s[20] ));
  nano32aa1n03x7               g132(.a(new_n225), .b(new_n195), .c(new_n220), .d(new_n204), .out0(new_n228));
  tech160nm_fioai012aa1n03p5x5 g133(.a(new_n228), .b(new_n192), .c(new_n184), .o1(new_n229));
  nanb03aa1n12x5               g134(.a(new_n218), .b(new_n219), .c(new_n211), .out0(new_n230));
  oai112aa1n06x5               g135(.a(new_n224), .b(new_n203), .c(new_n202), .d(new_n193), .o1(new_n231));
  aoi012aa1n06x5               g136(.a(new_n218), .b(new_n210), .c(new_n219), .o1(new_n232));
  oai012aa1d24x5               g137(.a(new_n232), .b(new_n231), .c(new_n230), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  xnbna2aa1n03x5               g141(.a(new_n236), .b(new_n229), .c(new_n234), .out0(\s[21] ));
  aoai13aa1n03x5               g142(.a(new_n236), .b(new_n233), .c(new_n216), .d(new_n228), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[21] ), .b(\a[22] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nor042aa1n09x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n239), .b(new_n241), .out0(new_n242));
  inv000aa1n06x5               g147(.a(new_n241), .o1(new_n243));
  aoai13aa1n02x7               g148(.a(new_n243), .b(new_n235), .c(new_n229), .d(new_n234), .o1(new_n244));
  aoi022aa1n03x5               g149(.a(new_n244), .b(new_n240), .c(new_n238), .d(new_n242), .o1(\s[22] ));
  nor042aa1n06x5               g150(.a(new_n239), .b(new_n235), .o1(new_n246));
  and002aa1n02x5               g151(.a(new_n228), .b(new_n246), .o(new_n247));
  oaih12aa1n02x5               g152(.a(new_n247), .b(new_n192), .c(new_n184), .o1(new_n248));
  oao003aa1n12x5               g153(.a(\a[22] ), .b(\b[21] ), .c(new_n243), .carry(new_n249));
  inv000aa1n02x5               g154(.a(new_n249), .o1(new_n250));
  tech160nm_fiaoi012aa1n04x5   g155(.a(new_n250), .b(new_n233), .c(new_n246), .o1(new_n251));
  inv000aa1n02x5               g156(.a(new_n251), .o1(new_n252));
  xorc02aa1n12x5               g157(.a(\a[23] ), .b(\b[22] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n252), .c(new_n216), .d(new_n247), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n253), .b(new_n250), .c(new_n233), .d(new_n246), .o1(new_n255));
  aobi12aa1n03x7               g160(.a(new_n254), .b(new_n255), .c(new_n248), .out0(\s[23] ));
  xorc02aa1n03x5               g161(.a(\a[24] ), .b(\b[23] ), .out0(new_n257));
  nor042aa1n09x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  norp02aa1n02x5               g163(.a(new_n257), .b(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n258), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n253), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n260), .b(new_n261), .c(new_n248), .d(new_n251), .o1(new_n262));
  aoi022aa1n02x7               g167(.a(new_n262), .b(new_n257), .c(new_n254), .d(new_n259), .o1(\s[24] ));
  inv000aa1n02x5               g168(.a(new_n228), .o1(new_n264));
  and002aa1n06x5               g169(.a(new_n257), .b(new_n253), .o(new_n265));
  nano22aa1n03x5               g170(.a(new_n264), .b(new_n246), .c(new_n265), .out0(new_n266));
  oaih12aa1n02x5               g171(.a(new_n266), .b(new_n192), .c(new_n184), .o1(new_n267));
  nano22aa1n02x4               g172(.a(new_n218), .b(new_n211), .c(new_n219), .out0(new_n268));
  tech160nm_fioai012aa1n03p5x5 g173(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .o1(new_n269));
  oab012aa1n03x5               g174(.a(new_n269), .b(new_n193), .c(new_n202), .out0(new_n270));
  inv000aa1n02x5               g175(.a(new_n232), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n246), .b(new_n271), .c(new_n270), .d(new_n268), .o1(new_n272));
  inv020aa1n04x5               g177(.a(new_n265), .o1(new_n273));
  oao003aa1n02x5               g178(.a(\a[24] ), .b(\b[23] ), .c(new_n260), .carry(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n273), .c(new_n272), .d(new_n249), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n216), .d(new_n266), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n265), .b(new_n250), .c(new_n233), .d(new_n246), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n276), .o1(new_n279));
  and003aa1n02x5               g184(.a(new_n278), .b(new_n279), .c(new_n274), .o(new_n280));
  aobi12aa1n03x7               g185(.a(new_n277), .b(new_n280), .c(new_n267), .out0(\s[25] ));
  tech160nm_fixorc02aa1n04x5   g186(.a(\a[26] ), .b(\b[25] ), .out0(new_n282));
  nor042aa1n06x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  norp02aa1n02x5               g188(.a(new_n282), .b(new_n283), .o1(new_n284));
  inv000aa1n02x5               g189(.a(new_n275), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n283), .o1(new_n286));
  aoai13aa1n02x7               g191(.a(new_n286), .b(new_n279), .c(new_n267), .d(new_n285), .o1(new_n287));
  aoi022aa1n02x7               g192(.a(new_n287), .b(new_n282), .c(new_n277), .d(new_n284), .o1(\s[26] ));
  and002aa1n12x5               g193(.a(new_n282), .b(new_n276), .o(new_n289));
  nano32aa1d15x5               g194(.a(new_n264), .b(new_n289), .c(new_n246), .d(new_n265), .out0(new_n290));
  oai012aa1n12x5               g195(.a(new_n290), .b(new_n192), .c(new_n184), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n289), .o1(new_n292));
  oao003aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .c(new_n286), .carry(new_n293));
  aoai13aa1n04x5               g198(.a(new_n293), .b(new_n292), .c(new_n278), .d(new_n274), .o1(new_n294));
  xorc02aa1n12x5               g199(.a(\a[27] ), .b(\b[26] ), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n216), .d(new_n290), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n293), .o1(new_n297));
  aoi112aa1n03x4               g202(.a(new_n295), .b(new_n297), .c(new_n275), .d(new_n289), .o1(new_n298));
  aobi12aa1n02x7               g203(.a(new_n296), .b(new_n298), .c(new_n291), .out0(\s[27] ));
  tech160nm_fixorc02aa1n03p5x5 g204(.a(\a[28] ), .b(\b[27] ), .out0(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  norp02aa1n02x5               g206(.a(new_n300), .b(new_n301), .o1(new_n302));
  tech160nm_fiaoi012aa1n05x5   g207(.a(new_n297), .b(new_n275), .c(new_n289), .o1(new_n303));
  inv000aa1n03x5               g208(.a(new_n301), .o1(new_n304));
  inv000aa1n02x5               g209(.a(new_n295), .o1(new_n305));
  aoai13aa1n02x7               g210(.a(new_n304), .b(new_n305), .c(new_n303), .d(new_n291), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n306), .b(new_n300), .c(new_n296), .d(new_n302), .o1(\s[28] ));
  and002aa1n02x5               g212(.a(new_n300), .b(new_n295), .o(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n294), .c(new_n216), .d(new_n290), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n308), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[28] ), .b(\b[27] ), .c(new_n304), .carry(new_n311));
  aoai13aa1n02x7               g216(.a(new_n311), .b(new_n310), .c(new_n303), .d(new_n291), .o1(new_n312));
  tech160nm_fixorc02aa1n03p5x5 g217(.a(\a[29] ), .b(\b[28] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n311), .b(new_n313), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[29] ));
  xorb03aa1n02x5               g220(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g221(.a(new_n305), .b(new_n300), .c(new_n313), .out0(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n294), .c(new_n216), .d(new_n290), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .carry(new_n320));
  aoai13aa1n04x5               g225(.a(new_n320), .b(new_n319), .c(new_n303), .d(new_n291), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n320), .b(new_n322), .out0(new_n323));
  aoi022aa1n02x7               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[30] ));
  xorc02aa1n02x5               g229(.a(\a[31] ), .b(\b[30] ), .out0(new_n325));
  nano32aa1n06x5               g230(.a(new_n305), .b(new_n322), .c(new_n300), .d(new_n313), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n294), .c(new_n216), .d(new_n290), .o1(new_n327));
  inv000aa1d42x5               g232(.a(new_n326), .o1(new_n328));
  oao003aa1n02x5               g233(.a(\a[30] ), .b(\b[29] ), .c(new_n320), .carry(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n328), .c(new_n303), .d(new_n291), .o1(new_n330));
  and002aa1n02x5               g235(.a(\b[29] ), .b(\a[30] ), .o(new_n331));
  oabi12aa1n02x5               g236(.a(new_n325), .b(\a[30] ), .c(\b[29] ), .out0(new_n332));
  oab012aa1n02x4               g237(.a(new_n332), .b(new_n320), .c(new_n331), .out0(new_n333));
  aoi022aa1n03x5               g238(.a(new_n330), .b(new_n325), .c(new_n327), .d(new_n333), .o1(\s[31] ));
  inv000aa1d42x5               g239(.a(\a[3] ), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n104), .b(\b[2] ), .c(new_n335), .out0(\s[3] ));
  norp02aa1n02x5               g241(.a(new_n100), .b(new_n104), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[4] ), .b(\b[3] ), .out0(new_n338));
  aoib12aa1n02x5               g243(.a(new_n338), .b(new_n335), .c(\b[2] ), .out0(new_n339));
  aboi22aa1n03x5               g244(.a(new_n337), .b(new_n339), .c(new_n105), .d(new_n338), .out0(\s[4] ));
  and002aa1n02x5               g245(.a(\b[4] ), .b(\a[5] ), .o(new_n341));
  and002aa1n02x5               g246(.a(\b[3] ), .b(\a[4] ), .o(new_n342));
  nona32aa1n03x5               g247(.a(new_n105), .b(new_n114), .c(new_n342), .d(new_n341), .out0(new_n343));
  xnrc02aa1n02x5               g248(.a(\b[4] ), .b(\a[5] ), .out0(new_n344));
  oabi12aa1n02x5               g249(.a(new_n342), .b(new_n337), .c(new_n99), .out0(new_n345));
  aobi12aa1n02x5               g250(.a(new_n343), .b(new_n345), .c(new_n344), .out0(\s[5] ));
  inv000aa1d42x5               g251(.a(new_n114), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n113), .b(new_n112), .out0(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n348), .b(new_n343), .c(new_n347), .out0(\s[6] ));
  nanb02aa1n02x5               g254(.a(new_n112), .b(new_n113), .out0(new_n350));
  aoai13aa1n03x5               g255(.a(new_n119), .b(new_n350), .c(new_n343), .d(new_n347), .o1(new_n351));
  xorb03aa1n02x5               g256(.a(new_n351), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp03aa1n03x5               g257(.a(new_n351), .b(new_n118), .c(new_n111), .o1(new_n353));
  norb02aa1n02x5               g258(.a(new_n106), .b(new_n107), .out0(new_n354));
  xnbna2aa1n03x5               g259(.a(new_n354), .b(new_n353), .c(new_n118), .out0(\s[8] ));
  xnbna2aa1n03x5               g260(.a(new_n123), .b(new_n179), .c(new_n180), .out0(\s[9] ));
endmodule


