// Benchmark "adder" written by ABC on Thu Jul 18 09:25:14 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n338, new_n339, new_n341,
    new_n342, new_n344;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\a[10] ), .b(new_n97), .out0(new_n98));
  nanp02aa1n09x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  nor022aa1n06x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[4] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(new_n103), .b(new_n102), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(new_n104), .b(new_n101), .o1(new_n105));
  inv000aa1d42x5               g010(.a(\a[3] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[2] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(new_n107), .b(new_n106), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(new_n108), .b(new_n109), .o1(new_n110));
  nor002aa1n02x5               g015(.a(\b[1] ), .b(\a[2] ), .o1(new_n111));
  nand42aa1n02x5               g016(.a(\b[1] ), .b(\a[2] ), .o1(new_n112));
  nand02aa1d06x5               g017(.a(\b[0] ), .b(\a[1] ), .o1(new_n113));
  tech160nm_fiaoi012aa1n04x5   g018(.a(new_n111), .b(new_n112), .c(new_n113), .o1(new_n114));
  norp03aa1n02x5               g019(.a(new_n114), .b(new_n105), .c(new_n110), .o1(new_n115));
  nor042aa1n04x5               g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  oaoi03aa1n12x5               g021(.a(new_n102), .b(new_n103), .c(new_n116), .o1(new_n117));
  inv000aa1d42x5               g022(.a(new_n117), .o1(new_n118));
  nanp02aa1n04x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nor042aa1n06x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nanb02aa1n02x5               g025(.a(new_n120), .b(new_n119), .out0(new_n121));
  nor002aa1n16x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  nand42aa1n03x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  nor002aa1n06x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  nand42aa1n03x5               g029(.a(\b[6] ), .b(\a[7] ), .o1(new_n125));
  nona23aa1n02x4               g030(.a(new_n125), .b(new_n123), .c(new_n122), .d(new_n124), .out0(new_n126));
  xnrc02aa1n02x5               g031(.a(\b[4] ), .b(\a[5] ), .out0(new_n127));
  nor043aa1n03x5               g032(.a(new_n126), .b(new_n127), .c(new_n121), .o1(new_n128));
  oai012aa1n02x7               g033(.a(new_n128), .b(new_n115), .c(new_n118), .o1(new_n129));
  nano23aa1n02x4               g034(.a(new_n122), .b(new_n124), .c(new_n125), .d(new_n123), .out0(new_n130));
  nor002aa1n03x5               g035(.a(\b[4] ), .b(\a[5] ), .o1(new_n131));
  nor022aa1n06x5               g036(.a(new_n131), .b(new_n120), .o1(new_n132));
  inv000aa1n02x5               g037(.a(new_n132), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n122), .o1(new_n134));
  aob012aa1n02x5               g039(.a(new_n134), .b(new_n124), .c(new_n123), .out0(new_n135));
  aoi013aa1n02x4               g040(.a(new_n135), .b(new_n130), .c(new_n133), .d(new_n119), .o1(new_n136));
  nanp02aa1n03x5               g041(.a(new_n129), .b(new_n136), .o1(new_n137));
  nand42aa1n03x5               g042(.a(\b[8] ), .b(\a[9] ), .o1(new_n138));
  tech160nm_fiaoi012aa1n05x5   g043(.a(new_n100), .b(new_n137), .c(new_n138), .o1(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n139), .b(new_n98), .c(new_n99), .out0(\s[10] ));
  nor002aa1n02x5               g045(.a(\b[9] ), .b(\a[10] ), .o1(new_n141));
  inv000aa1n02x5               g046(.a(new_n99), .o1(new_n142));
  nona22aa1n02x4               g047(.a(new_n139), .b(new_n142), .c(new_n141), .out0(new_n143));
  nor042aa1n04x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nand42aa1n04x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  norb02aa1n12x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n147), .b(new_n143), .c(new_n99), .out0(\s[11] ));
  nona22aa1n02x4               g053(.a(new_n143), .b(new_n147), .c(new_n142), .out0(new_n149));
  nor002aa1n04x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  nanp02aa1n09x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  norb02aa1n09x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  oaoi13aa1n04x5               g058(.a(new_n153), .b(new_n149), .c(\a[11] ), .d(\b[10] ), .o1(new_n154));
  aoi113aa1n02x5               g059(.a(new_n152), .b(new_n144), .c(new_n143), .d(new_n146), .e(new_n99), .o1(new_n155));
  norp02aa1n02x5               g060(.a(new_n154), .b(new_n155), .o1(\s[12] ));
  nand02aa1n02x5               g061(.a(new_n98), .b(new_n99), .o1(new_n157));
  nanb02aa1n06x5               g062(.a(new_n100), .b(new_n138), .out0(new_n158));
  nano23aa1n03x5               g063(.a(new_n144), .b(new_n150), .c(new_n151), .d(new_n145), .out0(new_n159));
  nona22aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n157), .out0(new_n160));
  norp02aa1n02x5               g065(.a(new_n100), .b(new_n141), .o1(new_n161));
  nona23aa1d18x5               g066(.a(new_n152), .b(new_n146), .c(new_n161), .d(new_n142), .out0(new_n162));
  aoi012aa1n02x5               g067(.a(new_n150), .b(new_n144), .c(new_n151), .o1(new_n163));
  nand02aa1d08x5               g068(.a(new_n162), .b(new_n163), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n160), .c(new_n129), .d(new_n136), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  xorc02aa1n12x5               g072(.a(\a[14] ), .b(\b[13] ), .out0(new_n168));
  norp02aa1n02x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  tech160nm_fixorc02aa1n03p5x5 g074(.a(\a[13] ), .b(\b[12] ), .out0(new_n170));
  aoi012aa1n02x5               g075(.a(new_n169), .b(new_n166), .c(new_n170), .o1(new_n171));
  xnrc02aa1n02x5               g076(.a(new_n171), .b(new_n168), .out0(\s[14] ));
  nor002aa1d32x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  nand42aa1n03x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  oai022aa1d24x5               g080(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n176));
  aob012aa1d15x5               g081(.a(new_n176), .b(\b[13] ), .c(\a[14] ), .out0(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  aoi013aa1n06x4               g083(.a(new_n178), .b(new_n166), .c(new_n170), .d(new_n168), .o1(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n174), .c(new_n175), .out0(\s[15] ));
  nanb02aa1n02x5               g085(.a(new_n173), .b(new_n175), .out0(new_n181));
  nor022aa1n04x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand42aa1n03x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nanb02aa1n02x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  oaoi13aa1n02x5               g089(.a(new_n184), .b(new_n174), .c(new_n179), .d(new_n181), .o1(new_n185));
  norp02aa1n02x5               g090(.a(new_n179), .b(new_n181), .o1(new_n186));
  nano22aa1n02x4               g091(.a(new_n186), .b(new_n174), .c(new_n184), .out0(new_n187));
  norp02aa1n03x5               g092(.a(new_n185), .b(new_n187), .o1(\s[16] ));
  oai013aa1n03x5               g093(.a(new_n117), .b(new_n114), .c(new_n105), .d(new_n110), .o1(new_n189));
  inv000aa1n02x5               g094(.a(new_n119), .o1(new_n190));
  norb02aa1n09x5               g095(.a(new_n123), .b(new_n122), .out0(new_n191));
  norb02aa1n06x4               g096(.a(new_n125), .b(new_n124), .out0(new_n192));
  nona23aa1n03x5               g097(.a(new_n192), .b(new_n191), .c(new_n132), .d(new_n190), .out0(new_n193));
  aoi012aa1n02x5               g098(.a(new_n122), .b(new_n124), .c(new_n123), .o1(new_n194));
  nand02aa1n02x5               g099(.a(new_n193), .b(new_n194), .o1(new_n195));
  nano23aa1n02x4               g100(.a(new_n173), .b(new_n182), .c(new_n183), .d(new_n175), .out0(new_n196));
  nano32aa1n03x7               g101(.a(new_n160), .b(new_n196), .c(new_n170), .d(new_n168), .out0(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n195), .c(new_n189), .d(new_n128), .o1(new_n198));
  nona23aa1n03x5               g103(.a(new_n183), .b(new_n175), .c(new_n173), .d(new_n182), .out0(new_n199));
  nano22aa1n03x7               g104(.a(new_n199), .b(new_n170), .c(new_n168), .out0(new_n200));
  nanp02aa1n02x5               g105(.a(new_n173), .b(new_n183), .o1(new_n201));
  oai122aa1n12x5               g106(.a(new_n201), .b(new_n199), .c(new_n177), .d(\b[15] ), .e(\a[16] ), .o1(new_n202));
  aoi012aa1d24x5               g107(.a(new_n202), .b(new_n164), .c(new_n200), .o1(new_n203));
  xnrc02aa1n02x5               g108(.a(\b[16] ), .b(\a[17] ), .out0(new_n204));
  xobna2aa1n03x5               g109(.a(new_n204), .b(new_n198), .c(new_n203), .out0(\s[17] ));
  inv000aa1d42x5               g110(.a(\a[17] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[16] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  aoai13aa1n02x5               g113(.a(new_n208), .b(new_n204), .c(new_n198), .d(new_n203), .o1(new_n209));
  xorb03aa1n02x5               g114(.a(new_n209), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  norp02aa1n24x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  nor042aa1n04x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  nand42aa1n06x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  aoai13aa1n12x5               g120(.a(new_n215), .b(new_n214), .c(new_n206), .d(new_n207), .o1(new_n216));
  nand22aa1n09x5               g121(.a(new_n198), .b(new_n203), .o1(new_n217));
  nanb02aa1n02x5               g122(.a(new_n214), .b(new_n215), .out0(new_n218));
  nona22aa1n03x5               g123(.a(new_n217), .b(new_n204), .c(new_n218), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n213), .b(new_n219), .c(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g125(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g126(.a(new_n211), .o1(new_n222));
  inv000aa1n02x5               g127(.a(new_n216), .o1(new_n223));
  aoi112aa1n02x5               g128(.a(new_n218), .b(new_n204), .c(new_n198), .d(new_n203), .o1(new_n224));
  oai012aa1n02x5               g129(.a(new_n213), .b(new_n224), .c(new_n223), .o1(new_n225));
  nor002aa1n03x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  nand22aa1n02x5               g131(.a(\b[19] ), .b(\a[20] ), .o1(new_n227));
  nanb02aa1n02x5               g132(.a(new_n226), .b(new_n227), .out0(new_n228));
  aoi012aa1n02x5               g133(.a(new_n228), .b(new_n225), .c(new_n222), .o1(new_n229));
  aobi12aa1n03x5               g134(.a(new_n213), .b(new_n219), .c(new_n216), .out0(new_n230));
  nano22aa1n03x7               g135(.a(new_n230), .b(new_n222), .c(new_n228), .out0(new_n231));
  norp02aa1n02x5               g136(.a(new_n229), .b(new_n231), .o1(\s[20] ));
  nano23aa1n02x4               g137(.a(new_n211), .b(new_n226), .c(new_n227), .d(new_n212), .out0(new_n233));
  nona22aa1n02x4               g138(.a(new_n233), .b(new_n204), .c(new_n218), .out0(new_n234));
  nona23aa1n03x5               g139(.a(new_n227), .b(new_n212), .c(new_n211), .d(new_n226), .out0(new_n235));
  tech160nm_fiaoi012aa1n03p5x5 g140(.a(new_n226), .b(new_n211), .c(new_n227), .o1(new_n236));
  oai012aa1n09x5               g141(.a(new_n236), .b(new_n235), .c(new_n216), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n234), .c(new_n198), .d(new_n203), .o1(new_n239));
  xorb03aa1n02x5               g144(.a(new_n239), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  xorc02aa1n02x5               g146(.a(\a[21] ), .b(\b[20] ), .out0(new_n242));
  xorc02aa1n02x5               g147(.a(\a[22] ), .b(\b[21] ), .out0(new_n243));
  aoai13aa1n02x5               g148(.a(new_n243), .b(new_n241), .c(new_n239), .d(new_n242), .o1(new_n244));
  aoi112aa1n02x5               g149(.a(new_n241), .b(new_n243), .c(new_n239), .d(new_n242), .o1(new_n245));
  norb02aa1n03x4               g150(.a(new_n244), .b(new_n245), .out0(\s[22] ));
  inv000aa1d42x5               g151(.a(\a[21] ), .o1(new_n247));
  inv040aa1d32x5               g152(.a(\a[22] ), .o1(new_n248));
  xroi22aa1d06x4               g153(.a(new_n247), .b(\b[20] ), .c(new_n248), .d(\b[21] ), .out0(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  nona22aa1n06x5               g155(.a(new_n217), .b(new_n234), .c(new_n250), .out0(new_n251));
  inv000aa1n02x5               g156(.a(new_n236), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n249), .b(new_n252), .c(new_n233), .d(new_n223), .o1(new_n253));
  inv000aa1d42x5               g158(.a(\b[21] ), .o1(new_n254));
  oaoi03aa1n09x5               g159(.a(new_n248), .b(new_n254), .c(new_n241), .o1(new_n255));
  nanp02aa1n02x5               g160(.a(new_n253), .b(new_n255), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  xnrc02aa1n12x5               g162(.a(\b[22] ), .b(\a[23] ), .out0(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n251), .c(new_n257), .out0(\s[23] ));
  nor042aa1n03x5               g165(.a(\b[22] ), .b(\a[23] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aoi112aa1n02x5               g167(.a(new_n250), .b(new_n234), .c(new_n198), .d(new_n203), .o1(new_n263));
  oaih12aa1n02x5               g168(.a(new_n259), .b(new_n263), .c(new_n256), .o1(new_n264));
  xnrc02aa1n02x5               g169(.a(\b[23] ), .b(\a[24] ), .out0(new_n265));
  aoi012aa1n02x5               g170(.a(new_n265), .b(new_n264), .c(new_n262), .o1(new_n266));
  tech160nm_fiaoi012aa1n05x5   g171(.a(new_n258), .b(new_n251), .c(new_n257), .o1(new_n267));
  nano22aa1n03x7               g172(.a(new_n267), .b(new_n262), .c(new_n265), .out0(new_n268));
  norp02aa1n02x5               g173(.a(new_n266), .b(new_n268), .o1(\s[24] ));
  techfinor002aa1n02p5x5       g174(.a(new_n265), .b(new_n258), .o1(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  nona32aa1n02x4               g176(.a(new_n217), .b(new_n271), .c(new_n250), .d(new_n234), .out0(new_n272));
  oao003aa1n02x5               g177(.a(\a[24] ), .b(\b[23] ), .c(new_n262), .carry(new_n273));
  aoai13aa1n04x5               g178(.a(new_n273), .b(new_n271), .c(new_n253), .d(new_n255), .o1(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  xnrc02aa1n12x5               g180(.a(\b[24] ), .b(\a[25] ), .out0(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  xnbna2aa1n03x5               g182(.a(new_n277), .b(new_n272), .c(new_n275), .out0(\s[25] ));
  nor042aa1n03x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(new_n249), .b(new_n270), .o1(new_n281));
  aoi112aa1n02x5               g186(.a(new_n281), .b(new_n234), .c(new_n198), .d(new_n203), .o1(new_n282));
  oaih12aa1n02x5               g187(.a(new_n277), .b(new_n282), .c(new_n274), .o1(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[25] ), .b(\a[26] ), .out0(new_n284));
  aoi012aa1n02x5               g189(.a(new_n284), .b(new_n283), .c(new_n280), .o1(new_n285));
  aoi012aa1n03x5               g190(.a(new_n276), .b(new_n272), .c(new_n275), .o1(new_n286));
  nano22aa1n03x5               g191(.a(new_n286), .b(new_n280), .c(new_n284), .out0(new_n287));
  norp02aa1n02x5               g192(.a(new_n285), .b(new_n287), .o1(\s[26] ));
  xorc02aa1n02x5               g193(.a(\a[27] ), .b(\b[26] ), .out0(new_n289));
  nor002aa1n02x5               g194(.a(new_n284), .b(new_n276), .o1(new_n290));
  inv000aa1n02x5               g195(.a(new_n290), .o1(new_n291));
  nona32aa1n09x5               g196(.a(new_n217), .b(new_n291), .c(new_n281), .d(new_n234), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[26] ), .b(\b[25] ), .c(new_n280), .carry(new_n293));
  aobi12aa1n09x5               g198(.a(new_n293), .b(new_n274), .c(new_n290), .out0(new_n294));
  xnbna2aa1n06x5               g199(.a(new_n289), .b(new_n294), .c(new_n292), .out0(\s[27] ));
  norp02aa1n02x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  inv040aa1n03x5               g201(.a(new_n296), .o1(new_n297));
  nanp03aa1n02x5               g202(.a(new_n249), .b(new_n270), .c(new_n290), .o1(new_n298));
  aoi112aa1n03x5               g203(.a(new_n298), .b(new_n234), .c(new_n198), .d(new_n203), .o1(new_n299));
  inv000aa1n02x5               g204(.a(new_n255), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n270), .b(new_n300), .c(new_n237), .d(new_n249), .o1(new_n301));
  aoai13aa1n04x5               g206(.a(new_n293), .b(new_n291), .c(new_n301), .d(new_n273), .o1(new_n302));
  oaih12aa1n02x5               g207(.a(new_n289), .b(new_n299), .c(new_n302), .o1(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[27] ), .b(\a[28] ), .out0(new_n304));
  tech160nm_fiaoi012aa1n02p5x5 g209(.a(new_n304), .b(new_n303), .c(new_n297), .o1(new_n305));
  aobi12aa1n06x5               g210(.a(new_n289), .b(new_n294), .c(new_n292), .out0(new_n306));
  nano22aa1n03x5               g211(.a(new_n306), .b(new_n297), .c(new_n304), .out0(new_n307));
  norp02aa1n03x5               g212(.a(new_n305), .b(new_n307), .o1(\s[28] ));
  xnrc02aa1n02x5               g213(.a(\b[28] ), .b(\a[29] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n289), .b(new_n304), .out0(new_n310));
  oai012aa1n02x5               g215(.a(new_n310), .b(new_n299), .c(new_n302), .o1(new_n311));
  oao003aa1n02x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n297), .carry(new_n312));
  aoi012aa1n02x5               g217(.a(new_n309), .b(new_n311), .c(new_n312), .o1(new_n313));
  aobi12aa1n06x5               g218(.a(new_n310), .b(new_n294), .c(new_n292), .out0(new_n314));
  nano22aa1n03x5               g219(.a(new_n314), .b(new_n309), .c(new_n312), .out0(new_n315));
  norp02aa1n03x5               g220(.a(new_n313), .b(new_n315), .o1(\s[29] ));
  xorb03aa1n02x5               g221(.a(new_n113), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .out0(new_n318));
  norb03aa1n02x5               g223(.a(new_n289), .b(new_n309), .c(new_n304), .out0(new_n319));
  oai012aa1n02x5               g224(.a(new_n319), .b(new_n299), .c(new_n302), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .carry(new_n321));
  tech160nm_fiaoi012aa1n02p5x5 g226(.a(new_n318), .b(new_n320), .c(new_n321), .o1(new_n322));
  aobi12aa1n06x5               g227(.a(new_n319), .b(new_n294), .c(new_n292), .out0(new_n323));
  nano22aa1n03x5               g228(.a(new_n323), .b(new_n318), .c(new_n321), .out0(new_n324));
  norp02aa1n03x5               g229(.a(new_n322), .b(new_n324), .o1(\s[30] ));
  norb02aa1n02x5               g230(.a(new_n319), .b(new_n318), .out0(new_n326));
  aobi12aa1n06x5               g231(.a(new_n326), .b(new_n294), .c(new_n292), .out0(new_n327));
  oao003aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n328));
  xnrc02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  nano22aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n329), .out0(new_n330));
  oai012aa1n02x5               g235(.a(new_n326), .b(new_n299), .c(new_n302), .o1(new_n331));
  aoi012aa1n02x5               g236(.a(new_n329), .b(new_n331), .c(new_n328), .o1(new_n332));
  norp02aa1n03x5               g237(.a(new_n332), .b(new_n330), .o1(\s[31] ));
  xnbna2aa1n03x5               g238(.a(new_n114), .b(new_n108), .c(new_n109), .out0(\s[3] ));
  oaoi03aa1n02x5               g239(.a(\a[3] ), .b(\b[2] ), .c(new_n114), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g241(.a(new_n189), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oabi12aa1n02x5               g242(.a(new_n127), .b(new_n115), .c(new_n118), .out0(new_n338));
  oai012aa1n02x5               g243(.a(new_n338), .b(\b[4] ), .c(\a[5] ), .o1(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g245(.a(new_n192), .b(new_n120), .c(new_n339), .d(new_n119), .o1(new_n341));
  aoi112aa1n02x5               g246(.a(new_n192), .b(new_n120), .c(new_n339), .d(new_n119), .o1(new_n342));
  norb02aa1n02x5               g247(.a(new_n341), .b(new_n342), .out0(\s[7] ));
  orn002aa1n02x5               g248(.a(\a[7] ), .b(\b[6] ), .o(new_n344));
  xnbna2aa1n03x5               g249(.a(new_n191), .b(new_n341), .c(new_n344), .out0(\s[8] ));
  xobna2aa1n03x5               g250(.a(new_n158), .b(new_n129), .c(new_n136), .out0(\s[9] ));
endmodule


