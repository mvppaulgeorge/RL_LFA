// Benchmark "adder" written by ABC on Thu Jul 18 03:55:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n181,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n297, new_n300, new_n301, new_n302, new_n304, new_n305, new_n306,
    new_n308;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n16x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nor002aa1d32x5               g002(.a(\b[6] ), .b(\a[7] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  tech160nm_fiaoi012aa1n03p5x5 g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nona23aa1d18x5               g006(.a(new_n99), .b(new_n101), .c(new_n98), .d(new_n97), .out0(new_n102));
  nanp02aa1n04x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  norp02aa1n04x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nor042aa1n02x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  oai012aa1n03x5               g010(.a(new_n103), .b(new_n105), .c(new_n104), .o1(new_n106));
  oaih12aa1n06x5               g011(.a(new_n100), .b(new_n102), .c(new_n106), .o1(new_n107));
  nor022aa1n16x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nand42aa1n04x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  nor022aa1n16x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nona23aa1d18x5               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  nand22aa1n03x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand02aa1d08x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nor042aa1n03x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  oai012aa1n06x5               g020(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n116));
  tech160nm_fioai012aa1n03p5x5 g021(.a(new_n109), .b(new_n110), .c(new_n108), .o1(new_n117));
  oaih12aa1n12x5               g022(.a(new_n117), .b(new_n112), .c(new_n116), .o1(new_n118));
  nanb02aa1n06x5               g023(.a(new_n104), .b(new_n103), .out0(new_n119));
  tech160nm_fixnrc02aa1n04x5   g024(.a(\b[4] ), .b(\a[5] ), .out0(new_n120));
  nor043aa1n09x5               g025(.a(new_n102), .b(new_n119), .c(new_n120), .o1(new_n121));
  aoi012aa1n02x5               g026(.a(new_n107), .b(new_n118), .c(new_n121), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[9] ), .b(\b[8] ), .c(new_n122), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor022aa1n08x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  aoi112aa1n09x5               g030(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n126));
  norp02aa1n02x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nand42aa1n20x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nand42aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nano23aa1n06x5               g034(.a(new_n127), .b(new_n125), .c(new_n129), .d(new_n128), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n107), .c(new_n118), .d(new_n121), .o1(new_n131));
  nona22aa1n02x4               g036(.a(new_n131), .b(new_n126), .c(new_n125), .out0(new_n132));
  xorb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand22aa1n12x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n134), .b(new_n132), .c(new_n135), .o1(new_n136));
  nor042aa1n09x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nand02aa1d06x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  norb02aa1n12x5               g043(.a(new_n138), .b(new_n137), .out0(new_n139));
  xnrc02aa1n02x5               g044(.a(new_n136), .b(new_n139), .out0(\s[12] ));
  norb02aa1n12x5               g045(.a(new_n135), .b(new_n134), .out0(new_n141));
  nano32aa1n02x4               g046(.a(new_n137), .b(new_n130), .c(new_n141), .d(new_n138), .out0(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n107), .c(new_n118), .d(new_n121), .o1(new_n143));
  aoi112aa1n09x5               g048(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n144));
  oai112aa1n06x5               g049(.a(new_n139), .b(new_n141), .c(new_n126), .d(new_n125), .o1(new_n145));
  nona22aa1d18x5               g050(.a(new_n145), .b(new_n144), .c(new_n137), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  nanp02aa1n02x5               g052(.a(new_n143), .b(new_n147), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor022aa1n08x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nanp02aa1n09x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  aoi012aa1n02x5               g056(.a(new_n150), .b(new_n148), .c(new_n151), .o1(new_n152));
  xnrb03aa1n02x5               g057(.a(new_n152), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor022aa1n08x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nanp02aa1n04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nona23aa1n02x5               g060(.a(new_n155), .b(new_n151), .c(new_n150), .d(new_n154), .out0(new_n156));
  aoi012aa1n02x7               g061(.a(new_n154), .b(new_n150), .c(new_n155), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n156), .c(new_n143), .d(new_n147), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n03x5               g064(.a(\b[14] ), .b(\a[15] ), .o1(new_n160));
  nand42aa1n16x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nor042aa1n12x5               g066(.a(\b[15] ), .b(\a[16] ), .o1(new_n162));
  nand02aa1d08x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nanb02aa1n12x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n160), .c(new_n158), .d(new_n161), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n165), .b(new_n160), .c(new_n158), .d(new_n161), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  nano23aa1n03x7               g073(.a(new_n150), .b(new_n154), .c(new_n155), .d(new_n151), .out0(new_n169));
  nano23aa1n06x5               g074(.a(new_n160), .b(new_n162), .c(new_n163), .d(new_n161), .out0(new_n170));
  nand02aa1n02x5               g075(.a(new_n170), .b(new_n169), .o1(new_n171));
  nano32aa1n03x7               g076(.a(new_n171), .b(new_n130), .c(new_n139), .d(new_n141), .out0(new_n172));
  aoai13aa1n12x5               g077(.a(new_n172), .b(new_n107), .c(new_n118), .d(new_n121), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n160), .b(new_n161), .out0(new_n174));
  nor043aa1n02x5               g079(.a(new_n156), .b(new_n164), .c(new_n174), .o1(new_n175));
  aoi112aa1n02x5               g080(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n176));
  obai22aa1n03x5               g081(.a(new_n170), .b(new_n157), .c(\a[16] ), .d(\b[15] ), .out0(new_n177));
  aoi112aa1n09x5               g082(.a(new_n177), .b(new_n176), .c(new_n146), .d(new_n175), .o1(new_n178));
  xorc02aa1n02x5               g083(.a(\a[17] ), .b(\b[16] ), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n178), .c(new_n173), .out0(\s[17] ));
  inv040aa1d32x5               g085(.a(\a[18] ), .o1(new_n181));
  nand22aa1n09x5               g086(.a(new_n178), .b(new_n173), .o1(new_n182));
  norp02aa1n02x5               g087(.a(\b[16] ), .b(\a[17] ), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n183), .b(new_n182), .c(new_n179), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[17] ), .c(new_n181), .out0(\s[18] ));
  inv000aa1d42x5               g090(.a(\a[17] ), .o1(new_n186));
  xroi22aa1d06x4               g091(.a(new_n186), .b(\b[16] ), .c(new_n181), .d(\b[17] ), .out0(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\b[17] ), .o1(new_n189));
  oao003aa1n02x5               g094(.a(new_n181), .b(new_n189), .c(new_n183), .carry(new_n190));
  inv000aa1d42x5               g095(.a(new_n190), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n188), .c(new_n178), .d(new_n173), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g098(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n04x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand02aa1d06x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nor042aa1n09x5               g101(.a(\b[19] ), .b(\a[20] ), .o1(new_n197));
  nand02aa1d06x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  norb02aa1n12x5               g103(.a(new_n198), .b(new_n197), .out0(new_n199));
  aoi112aa1n02x5               g104(.a(new_n195), .b(new_n199), .c(new_n192), .d(new_n196), .o1(new_n200));
  aoai13aa1n02x5               g105(.a(new_n199), .b(new_n195), .c(new_n192), .d(new_n196), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(\s[20] ));
  nano23aa1n09x5               g107(.a(new_n195), .b(new_n197), .c(new_n198), .d(new_n196), .out0(new_n203));
  nand02aa1d04x5               g108(.a(new_n187), .b(new_n203), .o1(new_n204));
  aoi112aa1n02x5               g109(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n205));
  nor002aa1n02x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  aoi112aa1n03x5               g111(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n207));
  norb02aa1n06x4               g112(.a(new_n196), .b(new_n195), .out0(new_n208));
  oai112aa1n06x5               g113(.a(new_n208), .b(new_n199), .c(new_n207), .d(new_n206), .o1(new_n209));
  nona22aa1d18x5               g114(.a(new_n209), .b(new_n205), .c(new_n197), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n204), .c(new_n178), .d(new_n173), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n06x5               g118(.a(\b[20] ), .b(\a[21] ), .o1(new_n214));
  nanp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  nor002aa1n06x5               g120(.a(\b[21] ), .b(\a[22] ), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(\b[21] ), .b(\a[22] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  aoi112aa1n02x5               g123(.a(new_n214), .b(new_n218), .c(new_n212), .d(new_n215), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n218), .b(new_n214), .c(new_n212), .d(new_n215), .o1(new_n220));
  norb02aa1n02x7               g125(.a(new_n220), .b(new_n219), .out0(\s[22] ));
  nona23aa1n06x5               g126(.a(new_n217), .b(new_n215), .c(new_n214), .d(new_n216), .out0(new_n222));
  inv030aa1n03x5               g127(.a(new_n222), .o1(new_n223));
  tech160nm_fiao0012aa1n02p5x5 g128(.a(new_n216), .b(new_n214), .c(new_n217), .o(new_n224));
  aoi012aa1n02x5               g129(.a(new_n224), .b(new_n210), .c(new_n223), .o1(new_n225));
  nand23aa1n06x5               g130(.a(new_n187), .b(new_n223), .c(new_n203), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n225), .b(new_n226), .c(new_n178), .d(new_n173), .o1(new_n227));
  xorb03aa1n02x5               g132(.a(new_n227), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g133(.a(\b[22] ), .b(\a[23] ), .o1(new_n229));
  xorc02aa1n02x5               g134(.a(\a[23] ), .b(\b[22] ), .out0(new_n230));
  xorc02aa1n02x5               g135(.a(\a[24] ), .b(\b[23] ), .out0(new_n231));
  aoi112aa1n02x7               g136(.a(new_n229), .b(new_n231), .c(new_n227), .d(new_n230), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n231), .b(new_n229), .c(new_n227), .d(new_n230), .o1(new_n233));
  norb02aa1n02x7               g138(.a(new_n233), .b(new_n232), .out0(\s[24] ));
  and002aa1n02x5               g139(.a(new_n231), .b(new_n230), .o(new_n235));
  nanb03aa1n06x5               g140(.a(new_n204), .b(new_n235), .c(new_n223), .out0(new_n236));
  norp02aa1n02x5               g141(.a(\b[23] ), .b(\a[24] ), .o1(new_n237));
  aoi112aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n238));
  nand03aa1n02x5               g143(.a(new_n224), .b(new_n230), .c(new_n231), .o1(new_n239));
  nona22aa1n06x5               g144(.a(new_n239), .b(new_n238), .c(new_n237), .out0(new_n240));
  nano22aa1n03x7               g145(.a(new_n222), .b(new_n230), .c(new_n231), .out0(new_n241));
  aoi012aa1n02x5               g146(.a(new_n240), .b(new_n210), .c(new_n241), .o1(new_n242));
  aoai13aa1n04x5               g147(.a(new_n242), .b(new_n236), .c(new_n178), .d(new_n173), .o1(new_n243));
  xorb03aa1n02x5               g148(.a(new_n243), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g149(.a(\b[24] ), .b(\a[25] ), .o1(new_n245));
  xorc02aa1n02x5               g150(.a(\a[25] ), .b(\b[24] ), .out0(new_n246));
  xorc02aa1n02x5               g151(.a(\a[26] ), .b(\b[25] ), .out0(new_n247));
  aoi112aa1n02x7               g152(.a(new_n245), .b(new_n247), .c(new_n243), .d(new_n246), .o1(new_n248));
  aoai13aa1n03x5               g153(.a(new_n247), .b(new_n245), .c(new_n243), .d(new_n246), .o1(new_n249));
  norb02aa1n03x4               g154(.a(new_n249), .b(new_n248), .out0(\s[26] ));
  and002aa1n02x5               g155(.a(new_n247), .b(new_n246), .o(new_n251));
  nano22aa1n12x5               g156(.a(new_n226), .b(new_n251), .c(new_n235), .out0(new_n252));
  norp02aa1n02x5               g157(.a(\b[25] ), .b(\a[26] ), .o1(new_n253));
  aoi112aa1n02x5               g158(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n254));
  aoai13aa1n04x5               g159(.a(new_n251), .b(new_n240), .c(new_n210), .d(new_n241), .o1(new_n255));
  nona22aa1d18x5               g160(.a(new_n255), .b(new_n254), .c(new_n253), .out0(new_n256));
  xorc02aa1n02x5               g161(.a(\a[27] ), .b(\b[26] ), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n256), .c(new_n182), .d(new_n252), .o1(new_n258));
  aoi112aa1n02x5               g163(.a(new_n256), .b(new_n257), .c(new_n182), .d(new_n252), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n258), .b(new_n259), .out0(\s[27] ));
  nor042aa1n03x5               g165(.a(\b[26] ), .b(\a[27] ), .o1(new_n261));
  xorc02aa1n12x5               g166(.a(\a[28] ), .b(\b[27] ), .out0(new_n262));
  nona22aa1n02x5               g167(.a(new_n258), .b(new_n262), .c(new_n261), .out0(new_n263));
  inv000aa1n03x5               g168(.a(new_n261), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n262), .o1(new_n265));
  tech160nm_fiaoi012aa1n02p5x5 g170(.a(new_n265), .b(new_n258), .c(new_n264), .o1(new_n266));
  norb02aa1n03x4               g171(.a(new_n263), .b(new_n266), .out0(\s[28] ));
  and002aa1n02x5               g172(.a(new_n262), .b(new_n257), .o(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n256), .c(new_n182), .d(new_n252), .o1(new_n269));
  oaoi03aa1n02x5               g174(.a(\a[28] ), .b(\b[27] ), .c(new_n264), .o1(new_n270));
  inv000aa1n03x5               g175(.a(new_n270), .o1(new_n271));
  xorc02aa1n02x5               g176(.a(\a[29] ), .b(\b[28] ), .out0(new_n272));
  inv000aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  tech160nm_fiaoi012aa1n05x5   g178(.a(new_n273), .b(new_n269), .c(new_n271), .o1(new_n274));
  nona22aa1n02x5               g179(.a(new_n269), .b(new_n270), .c(new_n272), .out0(new_n275));
  norb02aa1n03x4               g180(.a(new_n275), .b(new_n274), .out0(\s[29] ));
  xorb03aa1n02x5               g181(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g182(.a(new_n273), .b(new_n257), .c(new_n262), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n256), .c(new_n182), .d(new_n252), .o1(new_n279));
  oao003aa1n09x5               g184(.a(\a[29] ), .b(\b[28] ), .c(new_n271), .carry(new_n280));
  xorc02aa1n02x5               g185(.a(\a[30] ), .b(\b[29] ), .out0(new_n281));
  inv000aa1d42x5               g186(.a(new_n281), .o1(new_n282));
  tech160nm_fiaoi012aa1n05x5   g187(.a(new_n282), .b(new_n279), .c(new_n280), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n280), .o1(new_n284));
  nona22aa1n02x5               g189(.a(new_n279), .b(new_n284), .c(new_n281), .out0(new_n285));
  norb02aa1n03x4               g190(.a(new_n285), .b(new_n283), .out0(\s[30] ));
  xnrc02aa1n02x5               g191(.a(\b[30] ), .b(\a[31] ), .out0(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  nano32aa1n03x7               g193(.a(new_n282), .b(new_n272), .c(new_n262), .d(new_n257), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n256), .c(new_n182), .d(new_n252), .o1(new_n290));
  oaoi03aa1n02x5               g195(.a(\a[30] ), .b(\b[29] ), .c(new_n280), .o1(new_n291));
  nona22aa1n02x5               g196(.a(new_n290), .b(new_n291), .c(new_n288), .out0(new_n292));
  inv000aa1n02x5               g197(.a(new_n291), .o1(new_n293));
  tech160nm_fiaoi012aa1n02p5x5 g198(.a(new_n287), .b(new_n290), .c(new_n293), .o1(new_n294));
  norb02aa1n03x4               g199(.a(new_n292), .b(new_n294), .out0(\s[31] ));
  xnrb03aa1n02x5               g200(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g201(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n297));
  xorb03aa1n02x5               g202(.a(new_n297), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g203(.a(new_n118), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi13aa1n02x5               g204(.a(new_n120), .b(new_n117), .c(new_n112), .d(new_n116), .o1(new_n300));
  oai012aa1n02x5               g205(.a(new_n119), .b(new_n300), .c(new_n105), .o1(new_n301));
  nor043aa1n03x5               g206(.a(new_n300), .b(new_n119), .c(new_n105), .o1(new_n302));
  nanb02aa1n02x5               g207(.a(new_n302), .b(new_n301), .out0(\s[6] ));
  norb02aa1n02x5               g208(.a(new_n101), .b(new_n98), .out0(new_n304));
  nano22aa1n02x4               g209(.a(new_n302), .b(new_n304), .c(new_n103), .out0(new_n305));
  aoib12aa1n02x5               g210(.a(new_n304), .b(new_n103), .c(new_n302), .out0(new_n306));
  norp02aa1n02x5               g211(.a(new_n306), .b(new_n305), .o1(\s[7] ));
  norp02aa1n02x5               g212(.a(new_n305), .b(new_n98), .o1(new_n308));
  xnrb03aa1n03x5               g213(.a(new_n308), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g214(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


