// Benchmark "adder" written by ABC on Wed Jul 17 22:32:47 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n175, new_n176, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n305, new_n307, new_n310, new_n312, new_n314;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n04x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  nand42aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nor042aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  oai112aa1n03x5               g010(.a(new_n105), .b(new_n103), .c(new_n104), .d(new_n102), .o1(new_n106));
  oa0022aa1n02x5               g011(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n107));
  aoi022aa1n06x5               g012(.a(new_n106), .b(new_n107), .c(\b[3] ), .d(\a[4] ), .o1(new_n108));
  nand42aa1n16x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nor022aa1n08x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nanb03aa1n06x5               g016(.a(new_n110), .b(new_n111), .c(new_n109), .out0(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .out0(new_n113));
  orn002aa1n03x5               g018(.a(\a[5] ), .b(\b[4] ), .o(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  oai112aa1n03x5               g020(.a(new_n114), .b(new_n115), .c(\b[7] ), .d(\a[8] ), .o1(new_n116));
  norp03aa1n06x5               g021(.a(new_n116), .b(new_n112), .c(new_n113), .o1(new_n117));
  orn002aa1n02x5               g022(.a(\a[8] ), .b(\b[7] ), .o(new_n118));
  nanp02aa1n02x5               g023(.a(new_n110), .b(new_n109), .o1(new_n119));
  inv000aa1d42x5               g024(.a(new_n109), .o1(new_n120));
  norb02aa1n06x4               g025(.a(new_n111), .b(new_n110), .out0(new_n121));
  and002aa1n02x5               g026(.a(\b[5] ), .b(\a[6] ), .o(new_n122));
  oai022aa1n02x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  nona23aa1n02x4               g028(.a(new_n121), .b(new_n123), .c(new_n122), .d(new_n120), .out0(new_n124));
  nanp03aa1n03x5               g029(.a(new_n124), .b(new_n118), .c(new_n119), .o1(new_n125));
  nanp02aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n100), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n108), .d(new_n117), .o1(new_n128));
  xobna2aa1n03x5               g033(.a(new_n99), .b(new_n128), .c(new_n101), .out0(\s[10] ));
  nor042aa1n06x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nanp02aa1n04x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  nona22aa1n02x4               g037(.a(new_n128), .b(new_n100), .c(new_n97), .out0(new_n133));
  xobna2aa1n03x5               g038(.a(new_n132), .b(new_n133), .c(new_n98), .out0(\s[11] ));
  nor042aa1d18x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nand02aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  aoi013aa1n02x4               g042(.a(new_n130), .b(new_n133), .c(new_n132), .d(new_n98), .o1(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n136), .c(new_n137), .out0(\s[12] ));
  aoi012aa1n06x5               g044(.a(new_n125), .b(new_n108), .c(new_n117), .o1(new_n140));
  nano22aa1n12x5               g045(.a(new_n135), .b(new_n131), .c(new_n137), .out0(new_n141));
  nona23aa1n02x4               g046(.a(new_n141), .b(new_n127), .c(new_n99), .d(new_n130), .out0(new_n142));
  nanb03aa1n12x5               g047(.a(new_n135), .b(new_n137), .c(new_n131), .out0(new_n143));
  inv000aa1d42x5               g048(.a(new_n130), .o1(new_n144));
  oai112aa1n04x5               g049(.a(new_n144), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n145));
  aob012aa1n03x5               g050(.a(new_n136), .b(new_n130), .c(new_n137), .out0(new_n146));
  oabi12aa1n06x5               g051(.a(new_n146), .b(new_n145), .c(new_n143), .out0(new_n147));
  oabi12aa1n06x5               g052(.a(new_n147), .b(new_n140), .c(new_n142), .out0(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  inv040aa1d32x5               g054(.a(\a[14] ), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\a[13] ), .o1(new_n151));
  nanb02aa1n12x5               g056(.a(\b[12] ), .b(new_n151), .out0(new_n152));
  xorc02aa1n02x5               g057(.a(\a[13] ), .b(\b[12] ), .out0(new_n153));
  aobi12aa1n02x5               g058(.a(new_n152), .b(new_n148), .c(new_n153), .out0(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(new_n150), .out0(\s[14] ));
  xroi22aa1d06x4               g060(.a(new_n151), .b(\b[12] ), .c(new_n150), .d(\b[13] ), .out0(new_n156));
  oaoi03aa1n02x5               g061(.a(\a[14] ), .b(\b[13] ), .c(new_n152), .o1(new_n157));
  xorc02aa1n12x5               g062(.a(\a[15] ), .b(\b[14] ), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n157), .c(new_n148), .d(new_n156), .o1(new_n159));
  aoi112aa1n02x5               g064(.a(new_n158), .b(new_n157), .c(new_n148), .d(new_n156), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(\s[15] ));
  xorc02aa1n12x5               g066(.a(\a[16] ), .b(\b[15] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  oai112aa1n02x5               g068(.a(new_n159), .b(new_n163), .c(\b[14] ), .d(\a[15] ), .o1(new_n164));
  oaoi13aa1n06x5               g069(.a(new_n163), .b(new_n159), .c(\a[15] ), .d(\b[14] ), .o1(new_n165));
  norb02aa1n03x4               g070(.a(new_n164), .b(new_n165), .out0(\s[16] ));
  nand02aa1d04x5               g071(.a(new_n162), .b(new_n158), .o1(new_n167));
  nano32aa1n03x7               g072(.a(new_n143), .b(new_n144), .c(new_n101), .d(new_n126), .out0(new_n168));
  nona23aa1n09x5               g073(.a(new_n156), .b(new_n168), .c(new_n167), .d(new_n99), .out0(new_n169));
  tech160nm_fiaoi012aa1n02p5x5 g074(.a(new_n157), .b(new_n147), .c(new_n156), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n171));
  oab012aa1n02x4               g076(.a(new_n171), .b(\a[16] ), .c(\b[15] ), .out0(new_n172));
  oai122aa1n03x5               g077(.a(new_n172), .b(new_n140), .c(new_n169), .d(new_n170), .e(new_n167), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nand42aa1n02x5               g079(.a(new_n108), .b(new_n117), .o1(new_n175));
  norb03aa1n02x5               g080(.a(new_n123), .b(new_n112), .c(new_n122), .out0(new_n176));
  nano22aa1n03x7               g081(.a(new_n176), .b(new_n118), .c(new_n119), .out0(new_n177));
  aoi012aa1n12x5               g082(.a(new_n169), .b(new_n175), .c(new_n177), .o1(new_n178));
  inv030aa1n02x5               g083(.a(new_n157), .o1(new_n179));
  tech160nm_fioai012aa1n03p5x5 g084(.a(new_n98), .b(\b[10] ), .c(\a[11] ), .o1(new_n180));
  oab012aa1n04x5               g085(.a(new_n180), .b(new_n97), .c(new_n100), .out0(new_n181));
  aoai13aa1n04x5               g086(.a(new_n156), .b(new_n146), .c(new_n181), .d(new_n141), .o1(new_n182));
  aoai13aa1n12x5               g087(.a(new_n172), .b(new_n167), .c(new_n182), .d(new_n179), .o1(new_n183));
  nor042aa1n06x5               g088(.a(new_n183), .b(new_n178), .o1(new_n184));
  oaoi03aa1n03x5               g089(.a(\a[17] ), .b(\b[16] ), .c(new_n184), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv000aa1d42x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\a[18] ), .o1(new_n188));
  xroi22aa1d06x4               g093(.a(new_n187), .b(\b[16] ), .c(new_n188), .d(\b[17] ), .out0(new_n189));
  oai012aa1n06x5               g094(.a(new_n189), .b(new_n183), .c(new_n178), .o1(new_n190));
  inv000aa1d42x5               g095(.a(\b[17] ), .o1(new_n191));
  oai022aa1d24x5               g096(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n192));
  oaib12aa1n18x5               g097(.a(new_n192), .b(new_n191), .c(\a[18] ), .out0(new_n193));
  nor002aa1d32x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  nand42aa1n16x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nanb02aa1n02x5               g100(.a(new_n194), .b(new_n195), .out0(new_n196));
  xobna2aa1n03x5               g101(.a(new_n196), .b(new_n190), .c(new_n193), .out0(\s[19] ));
  xnrc02aa1n02x5               g102(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g103(.a(new_n194), .o1(new_n199));
  tech160nm_fiaoi012aa1n04x5   g104(.a(new_n196), .b(new_n190), .c(new_n193), .o1(new_n200));
  nor002aa1d32x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand42aa1n16x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nanb02aa1n02x5               g107(.a(new_n201), .b(new_n202), .out0(new_n203));
  nano22aa1n02x4               g108(.a(new_n200), .b(new_n199), .c(new_n203), .out0(new_n204));
  inv030aa1n06x5               g109(.a(new_n193), .o1(new_n205));
  oaoi13aa1n03x5               g110(.a(new_n205), .b(new_n189), .c(new_n183), .d(new_n178), .o1(new_n206));
  oaoi13aa1n02x7               g111(.a(new_n203), .b(new_n199), .c(new_n206), .d(new_n196), .o1(new_n207));
  norp02aa1n03x5               g112(.a(new_n207), .b(new_n204), .o1(\s[20] ));
  nona23aa1d18x5               g113(.a(new_n202), .b(new_n195), .c(new_n194), .d(new_n201), .out0(new_n209));
  norb02aa1n12x5               g114(.a(new_n189), .b(new_n209), .out0(new_n210));
  aoi012aa1n12x5               g115(.a(new_n201), .b(new_n194), .c(new_n202), .o1(new_n211));
  oai012aa1n18x5               g116(.a(new_n211), .b(new_n209), .c(new_n193), .o1(new_n212));
  oaoi13aa1n06x5               g117(.a(new_n212), .b(new_n210), .c(new_n183), .d(new_n178), .o1(new_n213));
  xnrb03aa1n03x5               g118(.a(new_n213), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  inv000aa1n02x5               g120(.a(new_n215), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n210), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n212), .o1(new_n218));
  xnrc02aa1n12x5               g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  oaoi13aa1n09x5               g124(.a(new_n219), .b(new_n218), .c(new_n184), .d(new_n217), .o1(new_n220));
  tech160nm_fixnrc02aa1n04x5   g125(.a(\b[21] ), .b(\a[22] ), .out0(new_n221));
  nano22aa1n03x5               g126(.a(new_n220), .b(new_n216), .c(new_n221), .out0(new_n222));
  oaoi13aa1n02x5               g127(.a(new_n221), .b(new_n216), .c(new_n213), .d(new_n219), .o1(new_n223));
  norp02aa1n03x5               g128(.a(new_n223), .b(new_n222), .o1(\s[22] ));
  nano23aa1d15x5               g129(.a(new_n194), .b(new_n201), .c(new_n202), .d(new_n195), .out0(new_n225));
  nor042aa1n04x5               g130(.a(new_n221), .b(new_n219), .o1(new_n226));
  nand23aa1n06x5               g131(.a(new_n189), .b(new_n226), .c(new_n225), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  inv030aa1n04x5               g133(.a(new_n211), .o1(new_n229));
  aoai13aa1n12x5               g134(.a(new_n226), .b(new_n229), .c(new_n225), .d(new_n205), .o1(new_n230));
  oao003aa1n12x5               g135(.a(\a[22] ), .b(\b[21] ), .c(new_n216), .carry(new_n231));
  nand22aa1n03x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  oaoi13aa1n06x5               g137(.a(new_n232), .b(new_n228), .c(new_n183), .d(new_n178), .o1(new_n233));
  xnrb03aa1n03x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n232), .o1(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[22] ), .b(\a[23] ), .out0(new_n238));
  oaoi13aa1n09x5               g143(.a(new_n238), .b(new_n237), .c(new_n184), .d(new_n227), .o1(new_n239));
  tech160nm_fixnrc02aa1n04x5   g144(.a(\b[23] ), .b(\a[24] ), .out0(new_n240));
  nano22aa1n03x5               g145(.a(new_n239), .b(new_n236), .c(new_n240), .out0(new_n241));
  oaoi13aa1n02x5               g146(.a(new_n240), .b(new_n236), .c(new_n233), .d(new_n238), .o1(new_n242));
  norp02aa1n03x5               g147(.a(new_n242), .b(new_n241), .o1(\s[24] ));
  norp02aa1n02x5               g148(.a(new_n240), .b(new_n238), .o1(new_n244));
  inv000aa1n03x5               g149(.a(new_n244), .o1(new_n245));
  nano32aa1n02x4               g150(.a(new_n245), .b(new_n189), .c(new_n226), .d(new_n225), .out0(new_n246));
  oai012aa1n06x5               g151(.a(new_n246), .b(new_n183), .c(new_n178), .o1(new_n247));
  oao003aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .c(new_n236), .carry(new_n248));
  aoai13aa1n12x5               g153(.a(new_n248), .b(new_n245), .c(new_n230), .d(new_n231), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n249), .o1(new_n250));
  tech160nm_fixnrc02aa1n05x5   g155(.a(\b[24] ), .b(\a[25] ), .out0(new_n251));
  xobna2aa1n03x5               g156(.a(new_n251), .b(new_n247), .c(new_n250), .out0(\s[25] ));
  nor042aa1n03x5               g157(.a(\b[24] ), .b(\a[25] ), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  aoi012aa1n03x5               g159(.a(new_n251), .b(new_n247), .c(new_n250), .o1(new_n255));
  tech160nm_fixnrc02aa1n05x5   g160(.a(\b[25] ), .b(\a[26] ), .out0(new_n256));
  nano22aa1n03x5               g161(.a(new_n255), .b(new_n254), .c(new_n256), .out0(new_n257));
  oaoi13aa1n03x5               g162(.a(new_n249), .b(new_n246), .c(new_n183), .d(new_n178), .o1(new_n258));
  oaoi13aa1n03x5               g163(.a(new_n256), .b(new_n254), .c(new_n258), .d(new_n251), .o1(new_n259));
  norp02aa1n03x5               g164(.a(new_n259), .b(new_n257), .o1(\s[26] ));
  nor042aa1n03x5               g165(.a(new_n256), .b(new_n251), .o1(new_n261));
  nano22aa1n03x7               g166(.a(new_n227), .b(new_n244), .c(new_n261), .out0(new_n262));
  oai012aa1n12x5               g167(.a(new_n262), .b(new_n183), .c(new_n178), .o1(new_n263));
  oao003aa1n02x5               g168(.a(\a[26] ), .b(\b[25] ), .c(new_n254), .carry(new_n264));
  aobi12aa1n12x5               g169(.a(new_n264), .b(new_n249), .c(new_n261), .out0(new_n265));
  xorc02aa1n02x5               g170(.a(\a[27] ), .b(\b[26] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n265), .c(new_n263), .out0(\s[27] ));
  norp02aa1n02x5               g172(.a(\b[26] ), .b(\a[27] ), .o1(new_n268));
  inv040aa1n03x5               g173(.a(new_n268), .o1(new_n269));
  aobi12aa1n03x5               g174(.a(new_n266), .b(new_n265), .c(new_n263), .out0(new_n270));
  xnrc02aa1n02x5               g175(.a(\b[27] ), .b(\a[28] ), .out0(new_n271));
  nano22aa1n03x5               g176(.a(new_n270), .b(new_n269), .c(new_n271), .out0(new_n272));
  inv000aa1d42x5               g177(.a(new_n231), .o1(new_n273));
  aoai13aa1n04x5               g178(.a(new_n244), .b(new_n273), .c(new_n212), .d(new_n226), .o1(new_n274));
  inv000aa1d42x5               g179(.a(new_n261), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n264), .b(new_n275), .c(new_n274), .d(new_n248), .o1(new_n276));
  aoai13aa1n03x5               g181(.a(new_n266), .b(new_n276), .c(new_n173), .d(new_n262), .o1(new_n277));
  tech160nm_fiaoi012aa1n02p5x5 g182(.a(new_n271), .b(new_n277), .c(new_n269), .o1(new_n278));
  norp02aa1n03x5               g183(.a(new_n278), .b(new_n272), .o1(\s[28] ));
  norb02aa1n02x5               g184(.a(new_n266), .b(new_n271), .out0(new_n280));
  aoai13aa1n02x5               g185(.a(new_n280), .b(new_n276), .c(new_n173), .d(new_n262), .o1(new_n281));
  oao003aa1n02x5               g186(.a(\a[28] ), .b(\b[27] ), .c(new_n269), .carry(new_n282));
  xnrc02aa1n02x5               g187(.a(\b[28] ), .b(\a[29] ), .out0(new_n283));
  tech160nm_fiaoi012aa1n02p5x5 g188(.a(new_n283), .b(new_n281), .c(new_n282), .o1(new_n284));
  aobi12aa1n02x7               g189(.a(new_n280), .b(new_n265), .c(new_n263), .out0(new_n285));
  nano22aa1n03x5               g190(.a(new_n285), .b(new_n282), .c(new_n283), .out0(new_n286));
  norp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[29] ));
  xorb03aa1n02x5               g192(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g193(.a(new_n266), .b(new_n283), .c(new_n271), .out0(new_n289));
  aoai13aa1n02x5               g194(.a(new_n289), .b(new_n276), .c(new_n173), .d(new_n262), .o1(new_n290));
  oao003aa1n02x5               g195(.a(\a[29] ), .b(\b[28] ), .c(new_n282), .carry(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[29] ), .b(\a[30] ), .out0(new_n292));
  tech160nm_fiaoi012aa1n02p5x5 g197(.a(new_n292), .b(new_n290), .c(new_n291), .o1(new_n293));
  aobi12aa1n03x5               g198(.a(new_n289), .b(new_n265), .c(new_n263), .out0(new_n294));
  nano22aa1n03x5               g199(.a(new_n294), .b(new_n291), .c(new_n292), .out0(new_n295));
  norp02aa1n03x5               g200(.a(new_n293), .b(new_n295), .o1(\s[30] ));
  xnrc02aa1n02x5               g201(.a(\b[30] ), .b(\a[31] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n289), .b(new_n292), .out0(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n276), .c(new_n173), .d(new_n262), .o1(new_n299));
  oao003aa1n02x5               g204(.a(\a[30] ), .b(\b[29] ), .c(new_n291), .carry(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n297), .b(new_n299), .c(new_n300), .o1(new_n301));
  aobi12aa1n02x7               g206(.a(new_n298), .b(new_n265), .c(new_n263), .out0(new_n302));
  nano22aa1n03x5               g207(.a(new_n302), .b(new_n297), .c(new_n300), .out0(new_n303));
  norp02aa1n03x5               g208(.a(new_n301), .b(new_n303), .o1(\s[31] ));
  oai012aa1n02x5               g209(.a(new_n103), .b(new_n104), .c(new_n102), .o1(new_n305));
  xnrb03aa1n02x5               g210(.a(new_n305), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g211(.a(\a[3] ), .b(\b[2] ), .c(new_n305), .o1(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g213(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaib12aa1n02x5               g214(.a(new_n115), .b(new_n108), .c(new_n114), .out0(new_n310));
  xnrb03aa1n02x5               g215(.a(new_n310), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oao003aa1n02x5               g216(.a(\a[6] ), .b(\b[5] ), .c(new_n310), .carry(new_n312));
  xnrc02aa1n02x5               g217(.a(new_n312), .b(new_n121), .out0(\s[7] ));
  oaoi03aa1n02x5               g218(.a(\a[7] ), .b(\b[6] ), .c(new_n312), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g220(.a(new_n127), .b(new_n177), .c(new_n175), .out0(\s[9] ));
endmodule


