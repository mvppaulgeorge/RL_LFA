// Benchmark "adder" written by ABC on Thu Jul 18 03:37:45 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n310, new_n312, new_n313, new_n314, new_n316, new_n317, new_n319,
    new_n321, new_n322, new_n323, new_n325, new_n326, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n06x5               g001(.a(\b[2] ), .b(\a[3] ), .out0(new_n97));
  nand42aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n09x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nor042aa1n04x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oai012aa1n06x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  oa0022aa1n02x5               g006(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n102));
  oai012aa1n06x5               g007(.a(new_n102), .b(new_n97), .c(new_n101), .o1(new_n103));
  nand02aa1n08x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand02aa1n08x5               g009(.a(\b[4] ), .b(\a[5] ), .o1(new_n105));
  orn002aa1n24x5               g010(.a(\a[5] ), .b(\b[4] ), .o(new_n106));
  nanp03aa1d24x5               g011(.a(new_n106), .b(new_n104), .c(new_n105), .o1(new_n107));
  norp02aa1n06x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  tech160nm_fiaoi012aa1n05x5   g013(.a(new_n108), .b(\a[6] ), .c(\b[5] ), .o1(new_n109));
  orn002aa1n24x5               g014(.a(\a[6] ), .b(\b[5] ), .o(new_n110));
  nor002aa1n16x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand02aa1d06x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanp02aa1n09x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanb03aa1n03x5               g018(.a(new_n111), .b(new_n113), .c(new_n112), .out0(new_n114));
  nano23aa1n06x5               g019(.a(new_n107), .b(new_n114), .c(new_n109), .d(new_n110), .out0(new_n115));
  nano22aa1n03x7               g020(.a(new_n111), .b(new_n112), .c(new_n113), .out0(new_n116));
  inv030aa1n02x5               g021(.a(new_n111), .o1(new_n117));
  oaoi03aa1n03x5               g022(.a(\a[8] ), .b(\b[7] ), .c(new_n117), .o1(new_n118));
  oai022aa1n06x5               g023(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n119));
  aoi013aa1n06x4               g024(.a(new_n118), .b(new_n116), .c(new_n109), .d(new_n119), .o1(new_n120));
  aobi12aa1n03x7               g025(.a(new_n120), .b(new_n115), .c(new_n103), .out0(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .c(new_n121), .o1(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1d18x5               g028(.a(\b[8] ), .b(\a[9] ), .o1(new_n124));
  nand02aa1n03x5               g029(.a(new_n115), .b(new_n103), .o1(new_n125));
  nanp02aa1n02x5               g030(.a(new_n125), .b(new_n120), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[9] ), .b(\b[8] ), .out0(new_n127));
  xorc02aa1n12x5               g032(.a(\a[10] ), .b(\b[9] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n124), .c(new_n126), .d(new_n127), .o1(new_n129));
  inv040aa1n08x5               g034(.a(new_n124), .o1(new_n130));
  oaoi03aa1n12x5               g035(.a(\a[10] ), .b(\b[9] ), .c(new_n130), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand02aa1n08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n15x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  xnbna2aa1n03x5               g040(.a(new_n135), .b(new_n129), .c(new_n132), .out0(\s[11] ));
  aoai13aa1n02x5               g041(.a(new_n135), .b(new_n131), .c(new_n122), .d(new_n128), .o1(new_n137));
  inv000aa1n02x5               g042(.a(new_n133), .o1(new_n138));
  inv000aa1d42x5               g043(.a(new_n135), .o1(new_n139));
  aoai13aa1n02x5               g044(.a(new_n138), .b(new_n139), .c(new_n129), .d(new_n132), .o1(new_n140));
  nor022aa1n12x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  nanp02aa1n06x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  norb02aa1n02x5               g047(.a(new_n142), .b(new_n141), .out0(new_n143));
  aoib12aa1n02x5               g048(.a(new_n133), .b(new_n142), .c(new_n141), .out0(new_n144));
  aoi022aa1n02x5               g049(.a(new_n140), .b(new_n143), .c(new_n137), .d(new_n144), .o1(\s[12] ));
  nona23aa1d18x5               g050(.a(new_n142), .b(new_n134), .c(new_n133), .d(new_n141), .out0(new_n146));
  nano22aa1d15x5               g051(.a(new_n146), .b(new_n127), .c(new_n128), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  nano23aa1n09x5               g053(.a(new_n133), .b(new_n141), .c(new_n142), .d(new_n134), .out0(new_n149));
  tech160nm_fioaoi03aa1n03p5x5 g054(.a(\a[12] ), .b(\b[11] ), .c(new_n138), .o1(new_n150));
  aoi012aa1n02x5               g055(.a(new_n150), .b(new_n149), .c(new_n131), .o1(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n148), .c(new_n125), .d(new_n120), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  inv000aa1n06x5               g059(.a(new_n154), .o1(new_n155));
  tech160nm_finand02aa1n03p5x5 g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n154), .out0(new_n157));
  nanp02aa1n02x5               g062(.a(new_n152), .b(new_n157), .o1(new_n158));
  xorc02aa1n02x5               g063(.a(\a[14] ), .b(\b[13] ), .out0(new_n159));
  xnbna2aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n155), .out0(\s[14] ));
  xnrc02aa1n02x5               g065(.a(\b[13] ), .b(\a[14] ), .out0(new_n161));
  nano22aa1n03x7               g066(.a(new_n161), .b(new_n155), .c(new_n156), .out0(new_n162));
  tech160nm_fioaoi03aa1n03p5x5 g067(.a(\a[14] ), .b(\b[13] ), .c(new_n155), .o1(new_n163));
  xorc02aa1n12x5               g068(.a(\a[15] ), .b(\b[14] ), .out0(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n163), .c(new_n152), .d(new_n162), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n164), .b(new_n163), .c(new_n152), .d(new_n162), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(\s[15] ));
  tech160nm_fioai012aa1n03p5x5 g072(.a(new_n165), .b(\b[14] ), .c(\a[15] ), .o1(new_n168));
  tech160nm_fixorc02aa1n05x5   g073(.a(\a[16] ), .b(\b[15] ), .out0(new_n169));
  oabi12aa1n02x5               g074(.a(new_n169), .b(\a[15] ), .c(\b[14] ), .out0(new_n170));
  aboi22aa1n03x5               g075(.a(new_n170), .b(new_n165), .c(new_n168), .d(new_n169), .out0(\s[16] ));
  nand02aa1n02x5               g076(.a(new_n159), .b(new_n157), .o1(new_n172));
  nand22aa1n03x5               g077(.a(new_n169), .b(new_n164), .o1(new_n173));
  nona22aa1n06x5               g078(.a(new_n147), .b(new_n172), .c(new_n173), .out0(new_n174));
  inv000aa1n02x5               g079(.a(new_n163), .o1(new_n175));
  aoai13aa1n06x5               g080(.a(new_n162), .b(new_n150), .c(new_n149), .d(new_n131), .o1(new_n176));
  ao0012aa1n03x7               g081(.a(new_n173), .b(new_n176), .c(new_n175), .o(new_n177));
  aoi112aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n178));
  oab012aa1n02x4               g083(.a(new_n178), .b(\a[16] ), .c(\b[15] ), .out0(new_n179));
  oai112aa1n06x5               g084(.a(new_n177), .b(new_n179), .c(new_n121), .d(new_n174), .o1(new_n180));
  xorb03aa1n03x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d30x5               g086(.a(\a[17] ), .o1(new_n182));
  nanb02aa1n12x5               g087(.a(\b[16] ), .b(new_n182), .out0(new_n183));
  aoi012aa1n09x5               g088(.a(new_n174), .b(new_n125), .c(new_n120), .o1(new_n184));
  aoai13aa1n09x5               g089(.a(new_n179), .b(new_n173), .c(new_n176), .d(new_n175), .o1(new_n185));
  xorc02aa1n02x5               g090(.a(\a[17] ), .b(\b[16] ), .out0(new_n186));
  oai012aa1n03x5               g091(.a(new_n186), .b(new_n185), .c(new_n184), .o1(new_n187));
  tech160nm_fixorc02aa1n02p5x5 g092(.a(\a[18] ), .b(\b[17] ), .out0(new_n188));
  xnbna2aa1n03x5               g093(.a(new_n188), .b(new_n187), .c(new_n183), .out0(\s[18] ));
  inv000aa1d42x5               g094(.a(\a[18] ), .o1(new_n190));
  xroi22aa1d04x5               g095(.a(new_n182), .b(\b[16] ), .c(new_n190), .d(\b[17] ), .out0(new_n191));
  tech160nm_fioai012aa1n05x5   g096(.a(new_n191), .b(new_n185), .c(new_n184), .o1(new_n192));
  oai022aa1n04x5               g097(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n193));
  oaib12aa1n09x5               g098(.a(new_n193), .b(new_n190), .c(\b[17] ), .out0(new_n194));
  nor002aa1d32x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nand42aa1n20x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  norb02aa1n02x5               g101(.a(new_n196), .b(new_n195), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n192), .c(new_n194), .out0(\s[19] ));
  xnrc02aa1n02x5               g103(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n12x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n183), .o1(new_n200));
  aoai13aa1n03x5               g105(.a(new_n197), .b(new_n200), .c(new_n180), .d(new_n191), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n195), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n197), .o1(new_n203));
  aoai13aa1n02x5               g108(.a(new_n202), .b(new_n203), .c(new_n192), .d(new_n194), .o1(new_n204));
  nor002aa1n20x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nand42aa1d28x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  aoib12aa1n02x5               g112(.a(new_n195), .b(new_n206), .c(new_n205), .out0(new_n208));
  aoi022aa1n03x5               g113(.a(new_n204), .b(new_n207), .c(new_n201), .d(new_n208), .o1(\s[20] ));
  nona23aa1d18x5               g114(.a(new_n206), .b(new_n196), .c(new_n195), .d(new_n205), .out0(new_n210));
  nano22aa1n09x5               g115(.a(new_n210), .b(new_n186), .c(new_n188), .out0(new_n211));
  tech160nm_fioai012aa1n05x5   g116(.a(new_n211), .b(new_n185), .c(new_n184), .o1(new_n212));
  aoi012aa1d24x5               g117(.a(new_n205), .b(new_n195), .c(new_n206), .o1(new_n213));
  oai012aa1d24x5               g118(.a(new_n213), .b(new_n210), .c(new_n194), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  xorc02aa1n02x5               g120(.a(\a[21] ), .b(\b[20] ), .out0(new_n216));
  xnbna2aa1n03x5               g121(.a(new_n216), .b(new_n212), .c(new_n215), .out0(\s[21] ));
  aoai13aa1n06x5               g122(.a(new_n216), .b(new_n214), .c(new_n180), .d(new_n211), .o1(new_n218));
  nor002aa1d32x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n216), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n220), .b(new_n221), .c(new_n212), .d(new_n215), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[22] ), .b(\b[21] ), .out0(new_n223));
  norp02aa1n02x5               g128(.a(new_n223), .b(new_n219), .o1(new_n224));
  aoi022aa1n03x5               g129(.a(new_n222), .b(new_n223), .c(new_n218), .d(new_n224), .o1(\s[22] ));
  nano23aa1n09x5               g130(.a(new_n195), .b(new_n205), .c(new_n206), .d(new_n196), .out0(new_n226));
  nand42aa1n02x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  nano22aa1n09x5               g133(.a(new_n228), .b(new_n220), .c(new_n227), .out0(new_n229));
  and003aa1n02x5               g134(.a(new_n191), .b(new_n229), .c(new_n226), .o(new_n230));
  oai012aa1n03x5               g135(.a(new_n230), .b(new_n185), .c(new_n184), .o1(new_n231));
  oao003aa1n12x5               g136(.a(\a[22] ), .b(\b[21] ), .c(new_n220), .carry(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoi012aa1n09x5               g138(.a(new_n233), .b(new_n214), .c(new_n229), .o1(new_n234));
  xorc02aa1n12x5               g139(.a(\a[23] ), .b(\b[22] ), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n231), .c(new_n234), .out0(\s[23] ));
  inv000aa1d42x5               g141(.a(new_n234), .o1(new_n237));
  aoai13aa1n02x7               g142(.a(new_n235), .b(new_n237), .c(new_n180), .d(new_n230), .o1(new_n238));
  nor042aa1n06x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n235), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n241), .c(new_n231), .d(new_n234), .o1(new_n242));
  tech160nm_fixorc02aa1n02p5x5 g147(.a(\a[24] ), .b(\b[23] ), .out0(new_n243));
  norp02aa1n02x5               g148(.a(new_n243), .b(new_n239), .o1(new_n244));
  aoi022aa1n03x5               g149(.a(new_n242), .b(new_n243), .c(new_n238), .d(new_n244), .o1(\s[24] ));
  and002aa1n12x5               g150(.a(new_n243), .b(new_n235), .o(new_n246));
  inv040aa1n08x5               g151(.a(new_n246), .o1(new_n247));
  nano32aa1n02x4               g152(.a(new_n247), .b(new_n191), .c(new_n226), .d(new_n229), .out0(new_n248));
  oai012aa1n03x5               g153(.a(new_n248), .b(new_n185), .c(new_n184), .o1(new_n249));
  inv020aa1n03x5               g154(.a(new_n213), .o1(new_n250));
  aoai13aa1n04x5               g155(.a(new_n229), .b(new_n250), .c(new_n226), .d(new_n200), .o1(new_n251));
  oao003aa1n02x5               g156(.a(\a[24] ), .b(\b[23] ), .c(new_n240), .carry(new_n252));
  aoai13aa1n12x5               g157(.a(new_n252), .b(new_n247), .c(new_n251), .d(new_n232), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  xnbna2aa1n03x5               g160(.a(new_n255), .b(new_n249), .c(new_n254), .out0(\s[25] ));
  aoai13aa1n02x7               g161(.a(new_n255), .b(new_n253), .c(new_n180), .d(new_n248), .o1(new_n257));
  nor042aa1n03x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n255), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n259), .b(new_n260), .c(new_n249), .d(new_n254), .o1(new_n261));
  xorc02aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .out0(new_n262));
  norp02aa1n02x5               g167(.a(new_n262), .b(new_n258), .o1(new_n263));
  aoi022aa1n03x5               g168(.a(new_n261), .b(new_n262), .c(new_n257), .d(new_n263), .o1(\s[26] ));
  and002aa1n03x5               g169(.a(new_n262), .b(new_n255), .o(new_n265));
  inv000aa1n02x5               g170(.a(new_n265), .o1(new_n266));
  nano32aa1n03x7               g171(.a(new_n266), .b(new_n211), .c(new_n229), .d(new_n246), .out0(new_n267));
  oai012aa1n12x5               g172(.a(new_n267), .b(new_n185), .c(new_n184), .o1(new_n268));
  oao003aa1n02x5               g173(.a(\a[26] ), .b(\b[25] ), .c(new_n259), .carry(new_n269));
  aobi12aa1n12x5               g174(.a(new_n269), .b(new_n253), .c(new_n265), .out0(new_n270));
  xorc02aa1n12x5               g175(.a(\a[27] ), .b(\b[26] ), .out0(new_n271));
  xnbna2aa1n06x5               g176(.a(new_n271), .b(new_n270), .c(new_n268), .out0(\s[27] ));
  aoai13aa1n03x5               g177(.a(new_n246), .b(new_n233), .c(new_n214), .d(new_n229), .o1(new_n273));
  aoai13aa1n04x5               g178(.a(new_n269), .b(new_n266), .c(new_n273), .d(new_n252), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n271), .b(new_n274), .c(new_n180), .d(new_n267), .o1(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  inv000aa1n03x5               g181(.a(new_n276), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n271), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n277), .b(new_n278), .c(new_n270), .d(new_n268), .o1(new_n279));
  tech160nm_fixorc02aa1n03p5x5 g184(.a(\a[28] ), .b(\b[27] ), .out0(new_n280));
  norp02aa1n02x5               g185(.a(new_n280), .b(new_n276), .o1(new_n281));
  aoi022aa1n03x5               g186(.a(new_n279), .b(new_n280), .c(new_n275), .d(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g187(.a(new_n280), .b(new_n271), .o(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n274), .c(new_n180), .d(new_n267), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n283), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[28] ), .b(\b[27] ), .c(new_n277), .carry(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n270), .d(new_n268), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[29] ), .b(\b[28] ), .out0(new_n288));
  norb02aa1n02x5               g193(.a(new_n286), .b(new_n288), .out0(new_n289));
  aoi022aa1n03x5               g194(.a(new_n287), .b(new_n288), .c(new_n284), .d(new_n289), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g196(.a(new_n278), .b(new_n280), .c(new_n288), .out0(new_n292));
  aoai13aa1n02x5               g197(.a(new_n292), .b(new_n274), .c(new_n180), .d(new_n267), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n292), .o1(new_n294));
  oao003aa1n02x5               g199(.a(\a[29] ), .b(\b[28] ), .c(new_n286), .carry(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n270), .d(new_n268), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[30] ), .b(\b[29] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n295), .b(new_n297), .out0(new_n298));
  aoi022aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n293), .d(new_n298), .o1(\s[30] ));
  xorc02aa1n02x5               g204(.a(\a[31] ), .b(\b[30] ), .out0(new_n300));
  nano32aa1n03x7               g205(.a(new_n278), .b(new_n297), .c(new_n280), .d(new_n288), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n274), .c(new_n180), .d(new_n267), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n301), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[30] ), .b(\b[29] ), .c(new_n295), .carry(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n303), .c(new_n270), .d(new_n268), .o1(new_n305));
  and002aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .o(new_n306));
  oabi12aa1n02x5               g211(.a(new_n300), .b(\a[30] ), .c(\b[29] ), .out0(new_n307));
  oab012aa1n02x4               g212(.a(new_n307), .b(new_n295), .c(new_n306), .out0(new_n308));
  aoi022aa1n03x5               g213(.a(new_n305), .b(new_n300), .c(new_n302), .d(new_n308), .o1(\s[31] ));
  inv000aa1d42x5               g214(.a(\a[3] ), .o1(new_n310));
  xorb03aa1n02x5               g215(.a(new_n101), .b(\b[2] ), .c(new_n310), .out0(\s[3] ));
  orn002aa1n02x5               g216(.a(new_n97), .b(new_n101), .o(new_n312));
  xorc02aa1n02x5               g217(.a(\a[4] ), .b(\b[3] ), .out0(new_n313));
  aoib12aa1n02x5               g218(.a(new_n313), .b(new_n310), .c(\b[2] ), .out0(new_n314));
  aoi022aa1n02x5               g219(.a(new_n312), .b(new_n314), .c(new_n103), .d(new_n313), .o1(\s[4] ));
  inv000aa1d42x5               g220(.a(new_n107), .o1(new_n316));
  aoi022aa1n02x5               g221(.a(new_n103), .b(new_n104), .c(new_n106), .d(new_n105), .o1(new_n317));
  aoi012aa1n02x5               g222(.a(new_n317), .b(new_n103), .c(new_n316), .o1(\s[5] ));
  aob012aa1n02x5               g223(.a(new_n106), .b(new_n103), .c(new_n316), .out0(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb02aa1n02x5               g225(.a(new_n111), .b(new_n112), .out0(new_n321));
  xorc02aa1n02x5               g226(.a(\a[6] ), .b(\b[5] ), .out0(new_n322));
  nanp02aa1n02x5               g227(.a(new_n319), .b(new_n322), .o1(new_n323));
  xobna2aa1n03x5               g228(.a(new_n321), .b(new_n323), .c(new_n110), .out0(\s[7] ));
  nanp02aa1n02x5               g229(.a(new_n323), .b(new_n110), .o1(new_n325));
  nanb02aa1n02x5               g230(.a(new_n321), .b(new_n325), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n113), .b(new_n108), .out0(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n327), .b(new_n326), .c(new_n117), .out0(\s[8] ));
  xnbna2aa1n03x5               g233(.a(new_n127), .b(new_n125), .c(new_n120), .out0(\s[9] ));
endmodule


