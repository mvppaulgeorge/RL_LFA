// Benchmark "adder" written by ABC on Wed Jul 17 22:21:38 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n321, new_n323, new_n326,
    new_n328, new_n329, new_n330, new_n331, new_n333, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d24x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n03x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  orn002aa1n02x5               g004(.a(\a[9] ), .b(\b[8] ), .o(new_n100));
  nor002aa1d24x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  nand02aa1n08x5               g006(.a(\b[5] ), .b(\a[6] ), .o1(new_n102));
  nor022aa1n16x5               g007(.a(\b[4] ), .b(\a[5] ), .o1(new_n103));
  nand42aa1n03x5               g008(.a(\b[4] ), .b(\a[5] ), .o1(new_n104));
  nona23aa1n09x5               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  nor042aa1d18x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand02aa1n10x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nanb02aa1n02x5               g012(.a(new_n106), .b(new_n107), .out0(new_n108));
  nor002aa1d32x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanp02aa1n12x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb02aa1n02x5               g015(.a(new_n109), .b(new_n110), .out0(new_n111));
  nor043aa1n03x5               g016(.a(new_n105), .b(new_n108), .c(new_n111), .o1(new_n112));
  oa0022aa1n06x5               g017(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n113));
  nand22aa1n12x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nand42aa1n20x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nor042aa1n06x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nanp02aa1n04x5               g021(.a(\b[2] ), .b(\a[3] ), .o1(new_n117));
  oai112aa1n06x5               g022(.a(new_n117), .b(new_n115), .c(new_n116), .d(new_n114), .o1(new_n118));
  aoi022aa1n06x5               g023(.a(new_n118), .b(new_n113), .c(\a[4] ), .d(\b[3] ), .o1(new_n119));
  nanb03aa1n12x5               g024(.a(new_n109), .b(new_n110), .c(new_n107), .out0(new_n120));
  inv040aa1n02x5               g025(.a(new_n106), .o1(new_n121));
  oai112aa1n06x5               g026(.a(new_n121), .b(new_n102), .c(new_n103), .d(new_n101), .o1(new_n122));
  tech160nm_fiaoi012aa1n03p5x5 g027(.a(new_n106), .b(new_n109), .c(new_n107), .o1(new_n123));
  oai012aa1n12x5               g028(.a(new_n123), .b(new_n122), .c(new_n120), .o1(new_n124));
  xnrc02aa1n12x5               g029(.a(\b[8] ), .b(\a[9] ), .out0(new_n125));
  inv000aa1d42x5               g030(.a(new_n125), .o1(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n124), .c(new_n112), .d(new_n119), .o1(new_n127));
  xobna2aa1n03x5               g032(.a(new_n99), .b(new_n127), .c(new_n100), .out0(\s[10] ));
  nor042aa1n06x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nand22aa1n04x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  nor002aa1d32x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  nona22aa1n03x5               g037(.a(new_n127), .b(new_n132), .c(new_n97), .out0(new_n133));
  xobna2aa1n03x5               g038(.a(new_n131), .b(new_n133), .c(new_n98), .out0(\s[11] ));
  nor002aa1d32x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  inv000aa1d42x5               g040(.a(new_n135), .o1(new_n136));
  nand22aa1n12x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  aoi013aa1n03x5               g042(.a(new_n129), .b(new_n133), .c(new_n130), .d(new_n98), .o1(new_n138));
  xnbna2aa1n03x5               g043(.a(new_n138), .b(new_n136), .c(new_n137), .out0(\s[12] ));
  nona23aa1n09x5               g044(.a(new_n137), .b(new_n130), .c(new_n129), .d(new_n135), .out0(new_n140));
  nor043aa1n06x5               g045(.a(new_n140), .b(new_n125), .c(new_n99), .o1(new_n141));
  aoai13aa1n06x5               g046(.a(new_n141), .b(new_n124), .c(new_n112), .d(new_n119), .o1(new_n142));
  nanb03aa1n02x5               g047(.a(new_n135), .b(new_n137), .c(new_n130), .out0(new_n143));
  oai122aa1n02x7               g048(.a(new_n98), .b(new_n97), .c(new_n132), .d(\b[10] ), .e(\a[11] ), .o1(new_n144));
  tech160nm_fiaoi012aa1n05x5   g049(.a(new_n135), .b(new_n129), .c(new_n137), .o1(new_n145));
  oai012aa1n02x7               g050(.a(new_n145), .b(new_n144), .c(new_n143), .o1(new_n146));
  inv000aa1n02x5               g051(.a(new_n146), .o1(new_n147));
  nor042aa1n06x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  nand22aa1n12x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n142), .c(new_n147), .out0(\s[13] ));
  nanp02aa1n02x5               g056(.a(new_n142), .b(new_n147), .o1(new_n152));
  aoi012aa1n02x5               g057(.a(new_n148), .b(new_n152), .c(new_n149), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n04x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nanp02aa1n09x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nona23aa1n03x5               g061(.a(new_n156), .b(new_n149), .c(new_n148), .d(new_n155), .out0(new_n157));
  tech160nm_fiaoi012aa1n03p5x5 g062(.a(new_n155), .b(new_n148), .c(new_n156), .o1(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n157), .c(new_n142), .d(new_n147), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nand02aa1n06x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nor022aa1n16x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nand42aa1n04x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  aoai13aa1n02x5               g070(.a(new_n165), .b(new_n161), .c(new_n159), .d(new_n162), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n161), .b(new_n165), .c(new_n159), .d(new_n162), .o1(new_n167));
  nanb02aa1n03x5               g072(.a(new_n167), .b(new_n166), .out0(\s[16] ));
  inv000aa1d42x5               g073(.a(\a[17] ), .o1(new_n169));
  nano23aa1n03x7               g074(.a(new_n106), .b(new_n109), .c(new_n110), .d(new_n107), .out0(new_n170));
  and002aa1n02x5               g075(.a(\b[3] ), .b(\a[4] ), .o(new_n171));
  nand42aa1n02x5               g076(.a(new_n118), .b(new_n113), .o1(new_n172));
  nona23aa1d18x5               g077(.a(new_n172), .b(new_n170), .c(new_n105), .d(new_n171), .out0(new_n173));
  inv030aa1n08x5               g078(.a(new_n124), .o1(new_n174));
  nona23aa1d24x5               g079(.a(new_n164), .b(new_n162), .c(new_n161), .d(new_n163), .out0(new_n175));
  nona22aa1n09x5               g080(.a(new_n141), .b(new_n157), .c(new_n175), .out0(new_n176));
  aoi012aa1d24x5               g081(.a(new_n176), .b(new_n173), .c(new_n174), .o1(new_n177));
  nano22aa1n03x7               g082(.a(new_n135), .b(new_n130), .c(new_n137), .out0(new_n178));
  oai012aa1n04x7               g083(.a(new_n98), .b(\b[10] ), .c(\a[11] ), .o1(new_n179));
  oab012aa1n06x5               g084(.a(new_n179), .b(new_n97), .c(new_n132), .out0(new_n180));
  inv020aa1n04x5               g085(.a(new_n145), .o1(new_n181));
  nano23aa1n06x5               g086(.a(new_n148), .b(new_n155), .c(new_n156), .d(new_n149), .out0(new_n182));
  aoai13aa1n12x5               g087(.a(new_n182), .b(new_n181), .c(new_n180), .d(new_n178), .o1(new_n183));
  tech160nm_fiaoi012aa1n03p5x5 g088(.a(new_n163), .b(new_n161), .c(new_n164), .o1(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n175), .c(new_n183), .d(new_n158), .o1(new_n185));
  norp02aa1n06x5               g090(.a(new_n185), .b(new_n177), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(new_n169), .out0(\s[17] ));
  oaoi03aa1n03x5               g092(.a(\a[17] ), .b(\b[16] ), .c(new_n186), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor002aa1d24x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  nor002aa1n16x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nand22aa1n09x5               g097(.a(\b[17] ), .b(\a[18] ), .o1(new_n193));
  nano23aa1n06x5               g098(.a(new_n190), .b(new_n192), .c(new_n193), .d(new_n191), .out0(new_n194));
  oai012aa1n06x5               g099(.a(new_n194), .b(new_n185), .c(new_n177), .o1(new_n195));
  oa0012aa1n02x5               g100(.a(new_n193), .b(new_n192), .c(new_n190), .o(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  nor042aa1n09x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand42aa1n04x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n06x4               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n200), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g106(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n03p5x5 g107(.a(new_n195), .b(new_n197), .o1(new_n203));
  nor042aa1n06x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand22aa1n12x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  aoai13aa1n03x5               g111(.a(new_n206), .b(new_n198), .c(new_n203), .d(new_n199), .o1(new_n207));
  aoi012aa1n06x5               g112(.a(new_n124), .b(new_n112), .c(new_n119), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n175), .o1(new_n209));
  aob012aa1n03x5               g114(.a(new_n209), .b(new_n183), .c(new_n158), .out0(new_n210));
  oai112aa1n06x5               g115(.a(new_n210), .b(new_n184), .c(new_n208), .d(new_n176), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n200), .b(new_n196), .c(new_n211), .d(new_n194), .o1(new_n212));
  nona22aa1n02x5               g117(.a(new_n212), .b(new_n206), .c(new_n198), .out0(new_n213));
  nanp02aa1n03x5               g118(.a(new_n207), .b(new_n213), .o1(\s[20] ));
  nano22aa1n03x7               g119(.a(new_n206), .b(new_n194), .c(new_n200), .out0(new_n215));
  oai012aa1n06x5               g120(.a(new_n215), .b(new_n185), .c(new_n177), .o1(new_n216));
  nanb03aa1n12x5               g121(.a(new_n204), .b(new_n205), .c(new_n199), .out0(new_n217));
  oai122aa1n12x5               g122(.a(new_n193), .b(new_n192), .c(new_n190), .d(\b[18] ), .e(\a[19] ), .o1(new_n218));
  aoi012aa1n06x5               g123(.a(new_n204), .b(new_n198), .c(new_n205), .o1(new_n219));
  oai012aa1d24x5               g124(.a(new_n219), .b(new_n218), .c(new_n217), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[20] ), .b(\a[21] ), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n216), .c(new_n221), .out0(\s[21] ));
  nand42aa1n02x5               g129(.a(new_n216), .b(new_n221), .o1(new_n225));
  nor042aa1n03x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[21] ), .b(\a[22] ), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n226), .c(new_n225), .d(new_n223), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n223), .b(new_n220), .c(new_n211), .d(new_n215), .o1(new_n229));
  nona22aa1n02x5               g134(.a(new_n229), .b(new_n227), .c(new_n226), .out0(new_n230));
  nanp02aa1n03x5               g135(.a(new_n228), .b(new_n230), .o1(\s[22] ));
  nor042aa1n06x5               g136(.a(new_n227), .b(new_n222), .o1(new_n232));
  nano32aa1n02x5               g137(.a(new_n206), .b(new_n232), .c(new_n194), .d(new_n200), .out0(new_n233));
  oai012aa1n06x5               g138(.a(new_n233), .b(new_n185), .c(new_n177), .o1(new_n234));
  inv000aa1d42x5               g139(.a(\a[22] ), .o1(new_n235));
  inv000aa1d42x5               g140(.a(\b[21] ), .o1(new_n236));
  oaoi03aa1n12x5               g141(.a(new_n235), .b(new_n236), .c(new_n226), .o1(new_n237));
  inv000aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1d18x5               g143(.a(new_n238), .b(new_n220), .c(new_n232), .o1(new_n239));
  xorc02aa1n12x5               g144(.a(\a[23] ), .b(\b[22] ), .out0(new_n240));
  xnbna2aa1n03x5               g145(.a(new_n240), .b(new_n234), .c(new_n239), .out0(\s[23] ));
  tech160nm_finand02aa1n03p5x5 g146(.a(new_n234), .b(new_n239), .o1(new_n242));
  norp02aa1n02x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  xnrc02aa1n12x5               g148(.a(\b[23] ), .b(\a[24] ), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n243), .c(new_n242), .d(new_n240), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n239), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n240), .b(new_n246), .c(new_n211), .d(new_n233), .o1(new_n247));
  nona22aa1n02x5               g152(.a(new_n247), .b(new_n244), .c(new_n243), .out0(new_n248));
  nanp02aa1n03x5               g153(.a(new_n245), .b(new_n248), .o1(\s[24] ));
  inv020aa1n03x5               g154(.a(new_n215), .o1(new_n250));
  norb02aa1n03x5               g155(.a(new_n240), .b(new_n244), .out0(new_n251));
  nano22aa1n03x7               g156(.a(new_n250), .b(new_n232), .c(new_n251), .out0(new_n252));
  oai012aa1n06x5               g157(.a(new_n252), .b(new_n185), .c(new_n177), .o1(new_n253));
  nano22aa1n03x5               g158(.a(new_n204), .b(new_n199), .c(new_n205), .out0(new_n254));
  oai012aa1n02x5               g159(.a(new_n193), .b(\b[18] ), .c(\a[19] ), .o1(new_n255));
  oab012aa1n02x4               g160(.a(new_n255), .b(new_n190), .c(new_n192), .out0(new_n256));
  inv000aa1n02x5               g161(.a(new_n219), .o1(new_n257));
  aoai13aa1n06x5               g162(.a(new_n232), .b(new_n257), .c(new_n256), .d(new_n254), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n251), .o1(new_n259));
  orn002aa1n02x5               g164(.a(\a[23] ), .b(\b[22] ), .o(new_n260));
  oao003aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .c(new_n260), .carry(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n259), .c(new_n258), .d(new_n237), .o1(new_n262));
  inv040aa1n03x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n12x5               g168(.a(\a[25] ), .b(\b[24] ), .out0(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n253), .c(new_n263), .out0(\s[25] ));
  nand42aa1n03x5               g170(.a(new_n253), .b(new_n263), .o1(new_n266));
  norp02aa1n02x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  tech160nm_fixnrc02aa1n05x5   g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n266), .d(new_n264), .o1(new_n269));
  aoai13aa1n03x5               g174(.a(new_n264), .b(new_n262), .c(new_n211), .d(new_n252), .o1(new_n270));
  nona22aa1n03x5               g175(.a(new_n270), .b(new_n268), .c(new_n267), .out0(new_n271));
  nanp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[26] ));
  norb02aa1n06x5               g177(.a(new_n264), .b(new_n268), .out0(new_n273));
  nano32aa1n06x5               g178(.a(new_n250), .b(new_n273), .c(new_n232), .d(new_n251), .out0(new_n274));
  tech160nm_fioai012aa1n04x5   g179(.a(new_n274), .b(new_n185), .c(new_n177), .o1(new_n275));
  inv000aa1d42x5               g180(.a(\a[26] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(\b[25] ), .o1(new_n277));
  oaoi03aa1n09x5               g182(.a(new_n276), .b(new_n277), .c(new_n267), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  aoi012aa1n09x5               g184(.a(new_n279), .b(new_n262), .c(new_n273), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[27] ), .b(\b[26] ), .out0(new_n281));
  xnbna2aa1n03x5               g186(.a(new_n281), .b(new_n280), .c(new_n275), .out0(\s[27] ));
  inv000aa1n02x5               g187(.a(new_n274), .o1(new_n283));
  oai012aa1n06x5               g188(.a(new_n280), .b(new_n186), .c(new_n283), .o1(new_n284));
  norp02aa1n02x5               g189(.a(\b[26] ), .b(\a[27] ), .o1(new_n285));
  nor002aa1n03x5               g190(.a(\b[27] ), .b(\a[28] ), .o1(new_n286));
  nand02aa1d24x5               g191(.a(\b[27] ), .b(\a[28] ), .o1(new_n287));
  norb02aa1n06x4               g192(.a(new_n287), .b(new_n286), .out0(new_n288));
  inv000aa1n06x5               g193(.a(new_n288), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n285), .c(new_n284), .d(new_n281), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n251), .b(new_n238), .c(new_n220), .d(new_n232), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n273), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n278), .b(new_n292), .c(new_n291), .d(new_n261), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n281), .b(new_n293), .c(new_n211), .d(new_n274), .o1(new_n294));
  nona22aa1n02x4               g199(.a(new_n294), .b(new_n289), .c(new_n285), .out0(new_n295));
  nanp02aa1n03x5               g200(.a(new_n290), .b(new_n295), .o1(\s[28] ));
  norb02aa1n09x5               g201(.a(new_n281), .b(new_n289), .out0(new_n297));
  aoai13aa1n02x5               g202(.a(new_n297), .b(new_n293), .c(new_n211), .d(new_n274), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n297), .o1(new_n299));
  oai012aa1n02x5               g204(.a(new_n287), .b(new_n286), .c(new_n285), .o1(new_n300));
  aoai13aa1n02x7               g205(.a(new_n300), .b(new_n299), .c(new_n280), .d(new_n275), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[29] ), .b(\b[28] ), .out0(new_n302));
  norb02aa1n02x5               g207(.a(new_n300), .b(new_n302), .out0(new_n303));
  aoi022aa1n03x5               g208(.a(new_n301), .b(new_n302), .c(new_n298), .d(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g210(.a(new_n281), .b(new_n302), .c(new_n288), .o(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n293), .c(new_n211), .d(new_n274), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n306), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n300), .carry(new_n309));
  aoai13aa1n02x7               g214(.a(new_n309), .b(new_n308), .c(new_n280), .d(new_n275), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[30] ), .b(\b[29] ), .out0(new_n311));
  norb02aa1n02x5               g216(.a(new_n309), .b(new_n311), .out0(new_n312));
  aoi022aa1n03x5               g217(.a(new_n310), .b(new_n311), .c(new_n307), .d(new_n312), .o1(\s[30] ));
  nand23aa1n03x5               g218(.a(new_n297), .b(new_n302), .c(new_n311), .o1(new_n314));
  nanb02aa1n03x5               g219(.a(new_n314), .b(new_n284), .out0(new_n315));
  xorc02aa1n02x5               g220(.a(\a[31] ), .b(\b[30] ), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[30] ), .b(\b[29] ), .c(new_n309), .carry(new_n317));
  norb02aa1n02x5               g222(.a(new_n317), .b(new_n316), .out0(new_n318));
  aoai13aa1n02x7               g223(.a(new_n317), .b(new_n314), .c(new_n280), .d(new_n275), .o1(new_n319));
  aoi022aa1n03x5               g224(.a(new_n319), .b(new_n316), .c(new_n315), .d(new_n318), .o1(\s[31] ));
  oai012aa1n02x5               g225(.a(new_n115), .b(new_n116), .c(new_n114), .o1(new_n321));
  xnrb03aa1n02x5               g226(.a(new_n321), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g227(.a(\a[3] ), .b(\b[2] ), .c(new_n321), .o1(new_n323));
  xorb03aa1n02x5               g228(.a(new_n323), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g229(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai012aa1n03x5               g230(.a(new_n104), .b(new_n119), .c(new_n103), .o1(new_n326));
  xnrb03aa1n02x5               g231(.a(new_n326), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaib12aa1n02x5               g232(.a(new_n102), .b(new_n101), .c(new_n326), .out0(new_n328));
  inv000aa1d42x5               g233(.a(new_n109), .o1(new_n329));
  nano22aa1n03x7               g234(.a(new_n101), .b(new_n326), .c(new_n102), .out0(new_n330));
  nano32aa1n03x7               g235(.a(new_n330), .b(new_n110), .c(new_n329), .d(new_n102), .out0(new_n331));
  aoi012aa1n02x5               g236(.a(new_n331), .b(new_n111), .c(new_n328), .o1(\s[7] ));
  oai012aa1n02x5               g237(.a(new_n108), .b(new_n331), .c(new_n109), .o1(new_n333));
  nano32aa1n02x4               g238(.a(new_n331), .b(new_n329), .c(new_n107), .d(new_n121), .out0(new_n334));
  nanb02aa1n03x5               g239(.a(new_n334), .b(new_n333), .out0(\s[8] ));
  xnbna2aa1n03x5               g240(.a(new_n126), .b(new_n173), .c(new_n174), .out0(\s[9] ));
endmodule


