// Benchmark "adder" written by ABC on Thu Jul 18 05:29:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n323, new_n324,
    new_n326, new_n328, new_n330, new_n331, new_n332, new_n334;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  orn002aa1n03x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nand02aa1n08x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand02aa1d16x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aob012aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  nor042aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n06x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nor042aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nand42aa1n06x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  norb02aa1n06x4               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  nand23aa1n06x5               g013(.a(new_n102), .b(new_n105), .c(new_n108), .o1(new_n109));
  tech160nm_fiaoi012aa1n05x5   g014(.a(new_n103), .b(new_n106), .c(new_n104), .o1(new_n110));
  nor002aa1n03x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand42aa1n16x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand42aa1n16x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nano23aa1n09x5               g019(.a(new_n111), .b(new_n113), .c(new_n114), .d(new_n112), .out0(new_n115));
  nor002aa1n12x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nand22aa1n12x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor042aa1d18x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nand22aa1n12x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano23aa1n06x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nand22aa1n03x5               g025(.a(new_n120), .b(new_n115), .o1(new_n121));
  ao0012aa1n03x7               g026(.a(new_n116), .b(new_n118), .c(new_n117), .o(new_n122));
  inv000aa1n02x5               g027(.a(new_n113), .o1(new_n123));
  oaoi03aa1n06x5               g028(.a(\a[8] ), .b(\b[7] ), .c(new_n123), .o1(new_n124));
  aoi012aa1n06x5               g029(.a(new_n124), .b(new_n115), .c(new_n122), .o1(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n126));
  nor002aa1n12x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nand42aa1n04x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  aoai13aa1n06x5               g034(.a(new_n129), .b(new_n97), .c(new_n126), .d(new_n98), .o1(new_n130));
  aoi112aa1n02x5               g035(.a(new_n129), .b(new_n97), .c(new_n126), .d(new_n98), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n130), .b(new_n131), .out0(\s[10] ));
  tech160nm_fioai012aa1n05x5   g037(.a(new_n128), .b(new_n127), .c(new_n97), .o1(new_n133));
  nor002aa1n20x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1n16x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n12x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n136), .b(new_n130), .c(new_n133), .out0(\s[11] ));
  inv000aa1d42x5               g042(.a(new_n134), .o1(new_n138));
  aob012aa1n02x5               g043(.a(new_n136), .b(new_n130), .c(new_n133), .out0(new_n139));
  norp02aa1n04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1n10x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n03x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  inv000aa1d42x5               g047(.a(new_n136), .o1(new_n143));
  norb03aa1n02x5               g048(.a(new_n141), .b(new_n134), .c(new_n140), .out0(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n143), .c(new_n130), .d(new_n133), .o1(new_n145));
  aoai13aa1n02x5               g050(.a(new_n145), .b(new_n142), .c(new_n139), .d(new_n138), .o1(\s[12] ));
  nano23aa1n03x7               g051(.a(new_n97), .b(new_n127), .c(new_n128), .d(new_n98), .out0(new_n147));
  and003aa1n02x5               g052(.a(new_n147), .b(new_n142), .c(new_n136), .o(new_n148));
  nano22aa1n03x7               g053(.a(new_n140), .b(new_n135), .c(new_n141), .out0(new_n149));
  nanb03aa1n06x5               g054(.a(new_n133), .b(new_n149), .c(new_n138), .out0(new_n150));
  oai012aa1n02x5               g055(.a(new_n141), .b(new_n140), .c(new_n134), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n150), .b(new_n151), .o1(new_n152));
  tech160nm_fiao0012aa1n02p5x5 g057(.a(new_n152), .b(new_n126), .c(new_n148), .o(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  nand02aa1n03x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nanb03aa1n02x5               g061(.a(new_n155), .b(new_n153), .c(new_n156), .out0(new_n157));
  nor042aa1n04x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand02aa1d08x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  aoib12aa1n02x5               g064(.a(new_n155), .b(new_n159), .c(new_n158), .out0(new_n160));
  nano23aa1n06x5               g065(.a(new_n155), .b(new_n158), .c(new_n159), .d(new_n156), .out0(new_n161));
  aoai13aa1n06x5               g066(.a(new_n161), .b(new_n152), .c(new_n126), .d(new_n148), .o1(new_n162));
  aoi012aa1n12x5               g067(.a(new_n158), .b(new_n155), .c(new_n159), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n158), .b(new_n162), .c(new_n163), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n164), .b(new_n157), .c(new_n160), .o1(\s[14] ));
  nor042aa1n12x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nand22aa1n04x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n162), .c(new_n163), .out0(\s[15] ));
  inv000aa1d42x5               g074(.a(new_n166), .o1(new_n170));
  inv000aa1n02x5               g075(.a(new_n168), .o1(new_n171));
  aoai13aa1n03x5               g076(.a(new_n170), .b(new_n171), .c(new_n162), .d(new_n163), .o1(new_n172));
  nor002aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand02aa1d08x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  nanb02aa1n02x5               g079(.a(new_n173), .b(new_n174), .out0(new_n175));
  norb03aa1n02x5               g080(.a(new_n174), .b(new_n166), .c(new_n173), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n171), .c(new_n162), .d(new_n163), .o1(new_n177));
  aob012aa1n03x5               g082(.a(new_n177), .b(new_n172), .c(new_n175), .out0(\s[16] ));
  nano23aa1n06x5               g083(.a(new_n166), .b(new_n173), .c(new_n174), .d(new_n167), .out0(new_n179));
  nand02aa1n03x5               g084(.a(new_n179), .b(new_n161), .o1(new_n180));
  nano32aa1n03x7               g085(.a(new_n180), .b(new_n147), .c(new_n142), .d(new_n136), .out0(new_n181));
  nanp02aa1n06x5               g086(.a(new_n126), .b(new_n181), .o1(new_n182));
  inv000aa1n06x5               g087(.a(new_n163), .o1(new_n183));
  oai012aa1n02x5               g088(.a(new_n174), .b(new_n173), .c(new_n166), .o1(new_n184));
  aobi12aa1n06x5               g089(.a(new_n184), .b(new_n179), .c(new_n183), .out0(new_n185));
  aoai13aa1n04x5               g090(.a(new_n185), .b(new_n180), .c(new_n150), .d(new_n151), .o1(new_n186));
  inv030aa1n03x5               g091(.a(new_n186), .o1(new_n187));
  nand02aa1d10x5               g092(.a(new_n182), .b(new_n187), .o1(new_n188));
  nor042aa1n04x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  nand42aa1n03x5               g094(.a(\b[16] ), .b(\a[17] ), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n190), .b(new_n189), .out0(new_n191));
  aob012aa1n02x5               g096(.a(new_n179), .b(new_n162), .c(new_n163), .out0(new_n192));
  oaoi13aa1n02x5               g097(.a(new_n191), .b(new_n174), .c(new_n166), .d(new_n173), .o1(new_n193));
  aoi022aa1n02x5               g098(.a(new_n192), .b(new_n193), .c(new_n191), .d(new_n188), .o1(\s[17] ));
  nor042aa1n04x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nanp02aa1n06x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  obai22aa1n02x7               g101(.a(new_n196), .b(new_n195), .c(\a[17] ), .d(\b[16] ), .out0(new_n197));
  aoi012aa1n02x5               g102(.a(new_n197), .b(new_n188), .c(new_n191), .o1(new_n198));
  nano23aa1n06x5               g103(.a(new_n189), .b(new_n195), .c(new_n196), .d(new_n190), .out0(new_n199));
  aoai13aa1n02x5               g104(.a(new_n199), .b(new_n186), .c(new_n126), .d(new_n181), .o1(new_n200));
  aoi012aa1n06x5               g105(.a(new_n195), .b(new_n189), .c(new_n196), .o1(new_n201));
  aoi012aa1n02x5               g106(.a(new_n195), .b(new_n200), .c(new_n201), .o1(new_n202));
  norp02aa1n02x5               g107(.a(new_n202), .b(new_n198), .o1(\s[18] ));
  nor042aa1n06x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nand42aa1n08x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  norb02aa1n06x5               g110(.a(new_n205), .b(new_n204), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n200), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n06x5               g113(.a(new_n204), .o1(new_n209));
  inv020aa1n08x5               g114(.a(new_n201), .o1(new_n210));
  aoai13aa1n06x5               g115(.a(new_n206), .b(new_n210), .c(new_n188), .d(new_n199), .o1(new_n211));
  nor002aa1n06x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nand42aa1n16x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  norb02aa1n06x5               g118(.a(new_n213), .b(new_n212), .out0(new_n214));
  norb03aa1n02x5               g119(.a(new_n213), .b(new_n204), .c(new_n212), .out0(new_n215));
  nanp02aa1n03x5               g120(.a(new_n211), .b(new_n215), .o1(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n214), .c(new_n211), .d(new_n209), .o1(\s[20] ));
  nano23aa1n06x5               g122(.a(new_n204), .b(new_n212), .c(new_n213), .d(new_n205), .out0(new_n218));
  and002aa1n02x5               g123(.a(new_n218), .b(new_n199), .o(new_n219));
  aoi112aa1n06x5               g124(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n220));
  oai112aa1n04x5               g125(.a(new_n206), .b(new_n214), .c(new_n220), .d(new_n195), .o1(new_n221));
  oaoi03aa1n03x5               g126(.a(\a[20] ), .b(\b[19] ), .c(new_n209), .o1(new_n222));
  inv030aa1n02x5               g127(.a(new_n222), .o1(new_n223));
  nanp02aa1n02x5               g128(.a(new_n221), .b(new_n223), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n224), .c(new_n188), .d(new_n219), .o1(new_n226));
  aoi112aa1n02x7               g131(.a(new_n225), .b(new_n224), .c(new_n188), .d(new_n219), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n226), .b(new_n227), .out0(\s[21] ));
  nor002aa1d32x5               g133(.a(\b[20] ), .b(\a[21] ), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[22] ), .b(\b[21] ), .out0(new_n231));
  nand42aa1n16x5               g136(.a(\b[21] ), .b(\a[22] ), .o1(new_n232));
  oai022aa1n02x5               g137(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n233));
  norb02aa1n02x5               g138(.a(new_n232), .b(new_n233), .out0(new_n234));
  nanp02aa1n03x5               g139(.a(new_n226), .b(new_n234), .o1(new_n235));
  aoai13aa1n03x5               g140(.a(new_n235), .b(new_n231), .c(new_n230), .d(new_n226), .o1(\s[22] ));
  nand42aa1n16x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  nor042aa1n03x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  nano23aa1n03x7               g143(.a(new_n229), .b(new_n238), .c(new_n232), .d(new_n237), .out0(new_n239));
  inv030aa1n02x5               g144(.a(new_n239), .o1(new_n240));
  nano22aa1n02x4               g145(.a(new_n240), .b(new_n199), .c(new_n218), .out0(new_n241));
  tech160nm_fioai012aa1n03p5x5 g146(.a(new_n232), .b(new_n238), .c(new_n229), .o1(new_n242));
  aoai13aa1n12x5               g147(.a(new_n242), .b(new_n240), .c(new_n221), .d(new_n223), .o1(new_n243));
  tech160nm_fixorc02aa1n02p5x5 g148(.a(\a[23] ), .b(\b[22] ), .out0(new_n244));
  aoai13aa1n06x5               g149(.a(new_n244), .b(new_n243), .c(new_n188), .d(new_n241), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n244), .b(new_n243), .c(new_n188), .d(new_n241), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n245), .b(new_n246), .out0(\s[23] ));
  nor042aa1n03x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  inv040aa1n03x5               g153(.a(new_n248), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[24] ), .b(\b[23] ), .out0(new_n250));
  oai022aa1n02x5               g155(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n251));
  aoi012aa1n02x5               g156(.a(new_n251), .b(\a[24] ), .c(\b[23] ), .o1(new_n252));
  nand42aa1n02x5               g157(.a(new_n245), .b(new_n252), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n250), .c(new_n249), .d(new_n245), .o1(\s[24] ));
  xnrc02aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .out0(new_n255));
  norb02aa1n03x5               g160(.a(new_n250), .b(new_n255), .out0(new_n256));
  inv000aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  nano23aa1n02x4               g162(.a(new_n257), .b(new_n240), .c(new_n218), .d(new_n199), .out0(new_n258));
  aoai13aa1n03x5               g163(.a(new_n239), .b(new_n222), .c(new_n218), .d(new_n210), .o1(new_n259));
  oaoi03aa1n02x5               g164(.a(\a[24] ), .b(\b[23] ), .c(new_n249), .o1(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  aoai13aa1n04x5               g166(.a(new_n261), .b(new_n257), .c(new_n259), .d(new_n242), .o1(new_n262));
  xorc02aa1n12x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n188), .d(new_n258), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n262), .c(new_n188), .d(new_n258), .o1(new_n265));
  norb02aa1n03x4               g170(.a(new_n264), .b(new_n265), .out0(\s[25] ));
  norp02aa1n02x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  tech160nm_fixorc02aa1n03p5x5 g173(.a(\a[26] ), .b(\b[25] ), .out0(new_n269));
  oai022aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n270));
  aoi012aa1n02x5               g175(.a(new_n270), .b(\a[26] ), .c(\b[25] ), .o1(new_n271));
  nanp02aa1n03x5               g176(.a(new_n264), .b(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n269), .c(new_n268), .d(new_n264), .o1(\s[26] ));
  nand03aa1n02x5               g178(.a(new_n239), .b(new_n244), .c(new_n250), .o1(new_n274));
  and002aa1n02x7               g179(.a(new_n269), .b(new_n263), .o(new_n275));
  nano32aa1n03x7               g180(.a(new_n274), .b(new_n275), .c(new_n199), .d(new_n218), .out0(new_n276));
  aoai13aa1n09x5               g181(.a(new_n276), .b(new_n186), .c(new_n126), .d(new_n181), .o1(new_n277));
  aoai13aa1n04x5               g182(.a(new_n275), .b(new_n260), .c(new_n243), .d(new_n256), .o1(new_n278));
  aob012aa1n02x5               g183(.a(new_n270), .b(\b[25] ), .c(\a[26] ), .out0(new_n279));
  nand23aa1n06x5               g184(.a(new_n277), .b(new_n278), .c(new_n279), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[27] ), .b(\b[26] ), .out0(new_n281));
  inv000aa1d42x5               g186(.a(new_n281), .o1(new_n282));
  and003aa1n02x5               g187(.a(new_n278), .b(new_n282), .c(new_n279), .o(new_n283));
  aoi022aa1n02x5               g188(.a(new_n283), .b(new_n277), .c(new_n280), .d(new_n281), .o1(\s[27] ));
  inv000aa1d42x5               g189(.a(\a[27] ), .o1(new_n285));
  nanb02aa1n02x5               g190(.a(\b[26] ), .b(new_n285), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n280), .b(new_n281), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .out0(new_n288));
  aobi12aa1n06x5               g193(.a(new_n279), .b(new_n262), .c(new_n275), .out0(new_n289));
  oai022aa1n02x5               g194(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(\a[28] ), .c(\b[27] ), .o1(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n282), .c(new_n289), .d(new_n277), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n292), .b(new_n288), .c(new_n287), .d(new_n286), .o1(\s[28] ));
  inv000aa1d42x5               g198(.a(\b[27] ), .o1(new_n294));
  xroi22aa1d04x5               g199(.a(new_n294), .b(\a[28] ), .c(new_n285), .d(\b[26] ), .out0(new_n295));
  inv000aa1d42x5               g200(.a(new_n295), .o1(new_n296));
  oaoi03aa1n02x5               g201(.a(\a[28] ), .b(\b[27] ), .c(new_n286), .o1(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[28] ), .b(\a[29] ), .out0(new_n298));
  norp02aa1n02x5               g203(.a(new_n297), .b(new_n298), .o1(new_n299));
  aoai13aa1n02x5               g204(.a(new_n299), .b(new_n296), .c(new_n289), .d(new_n277), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n298), .b(new_n297), .c(new_n280), .d(new_n295), .o1(new_n301));
  nanp02aa1n03x5               g206(.a(new_n301), .b(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g207(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n12x5               g208(.a(new_n298), .b(new_n281), .c(new_n288), .out0(new_n304));
  aob012aa1n02x5               g209(.a(new_n297), .b(\b[28] ), .c(\a[29] ), .out0(new_n305));
  oai012aa1n02x5               g210(.a(new_n305), .b(\b[28] ), .c(\a[29] ), .o1(new_n306));
  tech160nm_fixorc02aa1n03p5x5 g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n306), .c(new_n280), .d(new_n304), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n304), .o1(new_n310));
  norp02aa1n02x5               g215(.a(new_n306), .b(new_n308), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n310), .c(new_n289), .d(new_n277), .o1(new_n312));
  nanp02aa1n03x5               g217(.a(new_n309), .b(new_n312), .o1(\s[30] ));
  nano32aa1n03x7               g218(.a(new_n298), .b(new_n307), .c(new_n281), .d(new_n288), .out0(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  xnrc02aa1n02x5               g220(.a(\b[30] ), .b(\a[31] ), .out0(new_n316));
  aoi012aa1n02x5               g221(.a(new_n311), .b(\a[30] ), .c(\b[29] ), .o1(new_n317));
  norp02aa1n02x5               g222(.a(new_n317), .b(new_n316), .o1(new_n318));
  aoai13aa1n03x5               g223(.a(new_n318), .b(new_n315), .c(new_n289), .d(new_n277), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n316), .b(new_n317), .c(new_n280), .d(new_n314), .o1(new_n320));
  nanp02aa1n03x5               g225(.a(new_n320), .b(new_n319), .o1(\s[31] ));
  xorb03aa1n02x5               g226(.a(new_n102), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g227(.a(new_n109), .b(new_n110), .o1(new_n323));
  oaoi13aa1n02x5               g228(.a(new_n105), .b(new_n107), .c(new_n102), .d(new_n106), .o1(new_n324));
  aoib12aa1n02x5               g229(.a(new_n324), .b(new_n323), .c(new_n103), .out0(\s[4] ));
  norb02aa1n02x5               g230(.a(new_n119), .b(new_n118), .out0(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n326), .b(new_n109), .c(new_n110), .out0(\s[5] ));
  aoi012aa1n02x5               g232(.a(new_n118), .b(new_n323), .c(new_n119), .o1(new_n328));
  xnrb03aa1n02x5               g233(.a(new_n328), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g234(.a(new_n114), .b(new_n113), .out0(new_n330));
  aoai13aa1n02x5               g235(.a(new_n330), .b(new_n122), .c(new_n323), .d(new_n120), .o1(new_n331));
  aoi112aa1n02x5               g236(.a(new_n330), .b(new_n122), .c(new_n323), .d(new_n120), .o1(new_n332));
  norb02aa1n02x5               g237(.a(new_n331), .b(new_n332), .out0(\s[7] ));
  norb02aa1n02x5               g238(.a(new_n112), .b(new_n111), .out0(new_n334));
  xnbna2aa1n03x5               g239(.a(new_n334), .b(new_n331), .c(new_n123), .out0(\s[8] ));
  xorb03aa1n02x5               g240(.a(new_n126), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


