// Benchmark "adder" written by ABC on Wed Jul 17 20:42:02 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n320, new_n322, new_n323, new_n325,
    new_n327, new_n329, new_n331, new_n332, new_n333;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nand42aa1n08x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  norb02aa1n12x5               g005(.a(new_n100), .b(new_n99), .out0(new_n101));
  nand42aa1n16x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nor002aa1n20x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand42aa1n08x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nano22aa1n03x7               g009(.a(new_n103), .b(new_n102), .c(new_n104), .out0(new_n105));
  nand22aa1n12x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nor042aa1n06x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nona22aa1n09x5               g012(.a(new_n102), .b(new_n107), .c(new_n106), .out0(new_n108));
  nanp03aa1n06x5               g013(.a(new_n105), .b(new_n108), .c(new_n101), .o1(new_n109));
  tech160nm_fioai012aa1n04x5   g014(.a(new_n100), .b(new_n103), .c(new_n99), .o1(new_n110));
  nand02aa1d24x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor022aa1n16x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nand02aa1n08x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nano23aa1n03x7               g019(.a(new_n113), .b(new_n112), .c(new_n114), .d(new_n111), .out0(new_n115));
  nor002aa1n06x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand02aa1d12x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor002aa1n12x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nanp02aa1n12x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano23aa1n09x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nand02aa1n02x5               g025(.a(new_n120), .b(new_n115), .o1(new_n121));
  oa0012aa1n03x5               g026(.a(new_n117), .b(new_n118), .c(new_n116), .o(new_n122));
  oa0012aa1n03x5               g027(.a(new_n111), .b(new_n112), .c(new_n113), .o(new_n123));
  aoi012aa1n06x5               g028(.a(new_n122), .b(new_n120), .c(new_n123), .o1(new_n124));
  aoai13aa1n06x5               g029(.a(new_n124), .b(new_n121), .c(new_n109), .d(new_n110), .o1(new_n125));
  xnrc02aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  nanb02aa1n02x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  xnrc02aa1n12x5               g032(.a(\b[9] ), .b(\a[10] ), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  inv000aa1d42x5               g034(.a(\a[10] ), .o1(new_n130));
  inv000aa1d42x5               g035(.a(\b[9] ), .o1(new_n131));
  aoi012aa1n02x5               g036(.a(new_n97), .b(new_n130), .c(new_n131), .o1(new_n132));
  oai112aa1n02x5               g037(.a(new_n127), .b(new_n132), .c(new_n131), .d(new_n130), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n133), .b(new_n129), .c(new_n98), .d(new_n127), .o1(\s[10] ));
  norp02aa1n02x5               g039(.a(new_n128), .b(new_n126), .o1(new_n135));
  oaoi03aa1n09x5               g040(.a(new_n130), .b(new_n131), .c(new_n97), .o1(new_n136));
  aob012aa1n02x5               g041(.a(new_n136), .b(new_n125), .c(new_n135), .out0(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1d32x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  inv040aa1n03x5               g044(.a(new_n139), .o1(new_n140));
  nanp02aa1n06x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  and003aa1n02x5               g046(.a(new_n137), .b(new_n141), .c(new_n140), .o(new_n142));
  nor002aa1d32x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1n04x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  aoai13aa1n02x5               g050(.a(new_n145), .b(new_n139), .c(new_n137), .d(new_n141), .o1(new_n146));
  nona22aa1n02x4               g051(.a(new_n144), .b(new_n143), .c(new_n139), .out0(new_n147));
  oai012aa1n02x5               g052(.a(new_n146), .b(new_n142), .c(new_n147), .o1(\s[12] ));
  nano23aa1n06x5               g053(.a(new_n139), .b(new_n143), .c(new_n144), .d(new_n141), .out0(new_n149));
  nona22aa1n09x5               g054(.a(new_n149), .b(new_n128), .c(new_n126), .out0(new_n150));
  nona23aa1n09x5               g055(.a(new_n144), .b(new_n141), .c(new_n139), .d(new_n143), .out0(new_n151));
  oaoi03aa1n09x5               g056(.a(\a[12] ), .b(\b[11] ), .c(new_n140), .o1(new_n152));
  oabi12aa1n06x5               g057(.a(new_n152), .b(new_n151), .c(new_n136), .out0(new_n153));
  aoib12aa1n02x5               g058(.a(new_n153), .b(new_n125), .c(new_n150), .out0(new_n154));
  xnrb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .c(new_n154), .o1(new_n156));
  xnrc02aa1n12x5               g061(.a(\b[13] ), .b(\a[14] ), .out0(new_n157));
  tech160nm_fixnrc02aa1n05x5   g062(.a(\b[12] ), .b(\a[13] ), .out0(new_n158));
  nanp02aa1n02x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  oai022aa1n02x5               g064(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n160));
  nanb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  oabi12aa1n02x5               g066(.a(new_n161), .b(new_n154), .c(new_n158), .out0(new_n162));
  aob012aa1n02x5               g067(.a(new_n162), .b(new_n156), .c(new_n157), .out0(\s[14] ));
  nor042aa1n02x5               g068(.a(new_n157), .b(new_n158), .o1(new_n164));
  aoi022aa1n06x5               g069(.a(new_n153), .b(new_n164), .c(new_n159), .d(new_n160), .o1(new_n165));
  nona32aa1n02x4               g070(.a(new_n125), .b(new_n157), .c(new_n158), .d(new_n150), .out0(new_n166));
  xorc02aa1n02x5               g071(.a(\a[15] ), .b(\b[14] ), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n166), .c(new_n165), .out0(\s[15] ));
  nor022aa1n08x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  inv000aa1n06x5               g074(.a(new_n169), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(new_n166), .b(new_n165), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(new_n171), .b(new_n167), .o1(new_n172));
  xorc02aa1n02x5               g077(.a(\a[16] ), .b(\b[15] ), .out0(new_n173));
  and002aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .o(new_n174));
  oai022aa1n02x5               g079(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n175));
  nona22aa1n02x4               g080(.a(new_n172), .b(new_n174), .c(new_n175), .out0(new_n176));
  aoai13aa1n02x5               g081(.a(new_n176), .b(new_n173), .c(new_n170), .d(new_n172), .o1(\s[16] ));
  inv000aa1d42x5               g082(.a(\a[17] ), .o1(new_n178));
  nand42aa1n03x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  xnrc02aa1n12x5               g084(.a(\b[15] ), .b(\a[16] ), .out0(new_n180));
  nano22aa1n12x5               g085(.a(new_n180), .b(new_n170), .c(new_n179), .out0(new_n181));
  nano22aa1n06x5               g086(.a(new_n150), .b(new_n164), .c(new_n181), .out0(new_n182));
  oaoi03aa1n02x5               g087(.a(\a[16] ), .b(\b[15] ), .c(new_n170), .o1(new_n183));
  oaoi03aa1n02x5               g088(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n184));
  aoai13aa1n03x5               g089(.a(new_n164), .b(new_n152), .c(new_n149), .d(new_n184), .o1(new_n185));
  nanp02aa1n02x5               g090(.a(new_n160), .b(new_n159), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n181), .o1(new_n187));
  aoi012aa1n02x5               g092(.a(new_n187), .b(new_n185), .c(new_n186), .o1(new_n188));
  aoi112aa1n03x5               g093(.a(new_n188), .b(new_n183), .c(new_n125), .d(new_n182), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[16] ), .c(new_n178), .out0(\s[17] ));
  nor042aa1d18x5               g095(.a(\b[16] ), .b(\a[17] ), .o1(new_n191));
  inv040aa1n02x5               g096(.a(new_n191), .o1(new_n192));
  nanp02aa1n06x5               g097(.a(new_n125), .b(new_n182), .o1(new_n193));
  inv000aa1n02x5               g098(.a(new_n183), .o1(new_n194));
  oai112aa1n06x5               g099(.a(new_n193), .b(new_n194), .c(new_n187), .d(new_n165), .o1(new_n195));
  xorc02aa1n02x5               g100(.a(\a[17] ), .b(\b[16] ), .out0(new_n196));
  nanp02aa1n06x5               g101(.a(new_n195), .b(new_n196), .o1(new_n197));
  xorc02aa1n02x5               g102(.a(\a[18] ), .b(\b[17] ), .out0(new_n198));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\b[17] ), .o1(new_n200));
  aoi012aa1n02x5               g105(.a(new_n191), .b(new_n199), .c(new_n200), .o1(new_n201));
  oai112aa1n02x5               g106(.a(new_n197), .b(new_n201), .c(new_n200), .d(new_n199), .o1(new_n202));
  aoai13aa1n02x5               g107(.a(new_n202), .b(new_n198), .c(new_n192), .d(new_n197), .o1(\s[18] ));
  xroi22aa1d06x4               g108(.a(new_n178), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n204));
  tech160nm_fioaoi03aa1n04x5   g109(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n205));
  nor042aa1n09x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand42aa1d28x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nanb02aa1n02x5               g112(.a(new_n206), .b(new_n207), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n04x5               g114(.a(new_n209), .b(new_n205), .c(new_n195), .d(new_n204), .o1(new_n210));
  aoi112aa1n02x5               g115(.a(new_n209), .b(new_n205), .c(new_n195), .d(new_n204), .o1(new_n211));
  norb02aa1n03x4               g116(.a(new_n210), .b(new_n211), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g118(.a(new_n206), .o1(new_n214));
  nor042aa1n04x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  nand42aa1n16x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  norb03aa1n02x5               g122(.a(new_n216), .b(new_n206), .c(new_n215), .out0(new_n218));
  nanp02aa1n03x5               g123(.a(new_n210), .b(new_n218), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n219), .b(new_n217), .c(new_n214), .d(new_n210), .o1(\s[20] ));
  nano23aa1d15x5               g125(.a(new_n206), .b(new_n215), .c(new_n216), .d(new_n207), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  nano22aa1n02x4               g127(.a(new_n222), .b(new_n196), .c(new_n198), .out0(new_n223));
  tech160nm_fioaoi03aa1n04x5   g128(.a(\a[20] ), .b(\b[19] ), .c(new_n214), .o1(new_n224));
  tech160nm_fiao0012aa1n02p5x5 g129(.a(new_n224), .b(new_n221), .c(new_n205), .o(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  aoai13aa1n04x5               g132(.a(new_n227), .b(new_n225), .c(new_n195), .d(new_n223), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n227), .b(new_n225), .c(new_n195), .d(new_n223), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n228), .b(new_n229), .out0(\s[21] ));
  norp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[22] ), .b(\b[21] ), .out0(new_n233));
  nanp02aa1n02x5               g138(.a(\b[21] ), .b(\a[22] ), .o1(new_n234));
  oai022aa1n02x5               g139(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n235));
  norb02aa1n02x5               g140(.a(new_n234), .b(new_n235), .out0(new_n236));
  nanp02aa1n03x5               g141(.a(new_n228), .b(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n233), .c(new_n232), .d(new_n228), .o1(\s[22] ));
  orn002aa1n02x5               g143(.a(\a[22] ), .b(\b[21] ), .o(new_n239));
  nano22aa1n09x5               g144(.a(new_n226), .b(new_n239), .c(new_n234), .out0(new_n240));
  nanp03aa1d12x5               g145(.a(new_n204), .b(new_n240), .c(new_n221), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  aoai13aa1n06x5               g147(.a(new_n240), .b(new_n224), .c(new_n221), .d(new_n205), .o1(new_n243));
  nanp02aa1n02x5               g148(.a(new_n235), .b(new_n234), .o1(new_n244));
  nanp02aa1n02x5               g149(.a(new_n243), .b(new_n244), .o1(new_n245));
  tech160nm_fixnrc02aa1n05x5   g150(.a(\b[22] ), .b(\a[23] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  aoai13aa1n04x5               g152(.a(new_n247), .b(new_n245), .c(new_n195), .d(new_n242), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n247), .b(new_n245), .c(new_n195), .d(new_n242), .o1(new_n249));
  norb02aa1n03x4               g154(.a(new_n248), .b(new_n249), .out0(\s[23] ));
  norp02aa1n02x5               g155(.a(\b[22] ), .b(\a[23] ), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .out0(new_n253));
  nanp02aa1n02x5               g158(.a(\b[23] ), .b(\a[24] ), .o1(new_n254));
  oai022aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n254), .b(new_n255), .out0(new_n256));
  nanp02aa1n03x5               g161(.a(new_n248), .b(new_n256), .o1(new_n257));
  aoai13aa1n03x5               g162(.a(new_n257), .b(new_n253), .c(new_n252), .d(new_n248), .o1(\s[24] ));
  nanb02aa1n02x5               g163(.a(new_n246), .b(new_n253), .out0(new_n259));
  nano32aa1n02x4               g164(.a(new_n259), .b(new_n204), .c(new_n240), .d(new_n221), .out0(new_n260));
  nanp02aa1n02x5               g165(.a(new_n255), .b(new_n254), .o1(new_n261));
  aoai13aa1n12x5               g166(.a(new_n261), .b(new_n259), .c(new_n243), .d(new_n244), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  aoai13aa1n04x5               g168(.a(new_n263), .b(new_n262), .c(new_n195), .d(new_n260), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n262), .c(new_n195), .d(new_n260), .o1(new_n265));
  norb02aa1n03x4               g170(.a(new_n264), .b(new_n265), .out0(\s[25] ));
  orn002aa1n02x5               g171(.a(\a[25] ), .b(\b[24] ), .o(new_n267));
  xorc02aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  nanp02aa1n02x5               g173(.a(\b[25] ), .b(\a[26] ), .o1(new_n269));
  oai022aa1n02x5               g174(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n270));
  norb02aa1n02x5               g175(.a(new_n269), .b(new_n270), .out0(new_n271));
  nanp02aa1n03x5               g176(.a(new_n264), .b(new_n271), .o1(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n268), .c(new_n267), .d(new_n264), .o1(\s[26] ));
  and002aa1n02x5               g178(.a(new_n268), .b(new_n263), .o(new_n274));
  nano32aa1n06x5               g179(.a(new_n241), .b(new_n274), .c(new_n247), .d(new_n253), .out0(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  aoi022aa1n12x5               g181(.a(new_n262), .b(new_n274), .c(new_n269), .d(new_n270), .o1(new_n277));
  oai012aa1n12x5               g182(.a(new_n277), .b(new_n189), .c(new_n276), .o1(new_n278));
  xorb03aa1n02x5               g183(.a(new_n278), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  xorc02aa1n06x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  nanp02aa1n03x5               g187(.a(new_n278), .b(new_n282), .o1(new_n283));
  xorc02aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .out0(new_n284));
  nand02aa1n04x5               g189(.a(new_n195), .b(new_n275), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n282), .o1(new_n286));
  oai022aa1n02x5               g191(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n287));
  aoi012aa1n02x5               g192(.a(new_n287), .b(\a[28] ), .c(\b[27] ), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n286), .c(new_n285), .d(new_n277), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n284), .c(new_n283), .d(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g195(.a(new_n284), .b(new_n282), .o(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  inv000aa1d42x5               g197(.a(\b[27] ), .o1(new_n293));
  oaib12aa1n09x5               g198(.a(new_n287), .b(new_n293), .c(\a[28] ), .out0(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[28] ), .b(\a[29] ), .out0(new_n295));
  norb02aa1n02x5               g200(.a(new_n294), .b(new_n295), .out0(new_n296));
  aoai13aa1n02x5               g201(.a(new_n296), .b(new_n292), .c(new_n285), .d(new_n277), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n294), .o1(new_n298));
  aoai13aa1n03x5               g203(.a(new_n295), .b(new_n298), .c(new_n278), .d(new_n291), .o1(new_n299));
  nanp02aa1n03x5               g204(.a(new_n299), .b(new_n297), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g206(.a(new_n295), .b(new_n282), .c(new_n284), .out0(new_n302));
  oaoi03aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .c(new_n294), .o1(new_n303));
  tech160nm_fixorc02aa1n05x5   g208(.a(\a[30] ), .b(\b[29] ), .out0(new_n304));
  inv000aa1d42x5               g209(.a(new_n304), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n303), .c(new_n278), .d(new_n302), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n302), .o1(new_n307));
  norp02aa1n02x5               g212(.a(new_n303), .b(new_n305), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n307), .c(new_n285), .d(new_n277), .o1(new_n309));
  nanp02aa1n03x5               g214(.a(new_n306), .b(new_n309), .o1(\s[30] ));
  nano32aa1n02x5               g215(.a(new_n295), .b(new_n304), .c(new_n282), .d(new_n284), .out0(new_n311));
  nanp02aa1n03x5               g216(.a(new_n278), .b(new_n311), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[31] ), .b(\b[30] ), .out0(new_n313));
  inv000aa1n02x5               g218(.a(new_n311), .o1(new_n314));
  oai012aa1n02x5               g219(.a(new_n313), .b(\b[29] ), .c(\a[30] ), .o1(new_n315));
  aoi012aa1n02x5               g220(.a(new_n315), .b(new_n303), .c(new_n304), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n314), .c(new_n285), .d(new_n277), .o1(new_n317));
  oao003aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .c(new_n308), .carry(new_n318));
  aoai13aa1n03x5               g223(.a(new_n317), .b(new_n313), .c(new_n312), .d(new_n318), .o1(\s[31] ));
  norb02aa1n02x5               g224(.a(new_n104), .b(new_n103), .out0(new_n320));
  xobna2aa1n03x5               g225(.a(new_n320), .b(new_n108), .c(new_n102), .out0(\s[3] ));
  inv000aa1d42x5               g226(.a(new_n103), .o1(new_n322));
  oai112aa1n02x5               g227(.a(new_n320), .b(new_n102), .c(new_n106), .d(new_n107), .o1(new_n323));
  xnbna2aa1n03x5               g228(.a(new_n101), .b(new_n323), .c(new_n322), .out0(\s[4] ));
  nanp02aa1n02x5               g229(.a(new_n109), .b(new_n110), .o1(new_n325));
  xorb03aa1n02x5               g230(.a(new_n325), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoi012aa1n02x5               g231(.a(new_n113), .b(new_n325), .c(new_n114), .o1(new_n327));
  xnrb03aa1n02x5               g232(.a(new_n327), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g233(.a(new_n123), .b(new_n325), .c(new_n115), .o(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g235(.a(new_n116), .b(new_n117), .out0(new_n331));
  aoai13aa1n02x5               g236(.a(new_n331), .b(new_n118), .c(new_n329), .d(new_n119), .o1(new_n332));
  aoi112aa1n02x5               g237(.a(new_n331), .b(new_n118), .c(new_n329), .d(new_n119), .o1(new_n333));
  nanb02aa1n02x5               g238(.a(new_n333), .b(new_n332), .out0(\s[8] ));
  xorb03aa1n02x5               g239(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


