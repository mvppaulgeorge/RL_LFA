// Benchmark "adder" written by ABC on Wed Jul 17 18:59:04 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n336, new_n338,
    new_n340, new_n342, new_n344, new_n345, new_n346, new_n348, new_n349,
    new_n350;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  nor022aa1n06x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand42aa1n06x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aob012aa1n12x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  nor042aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nanp02aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n03x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor002aa1n06x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanp02aa1n06x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n06x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nanp03aa1n09x5               g014(.a(new_n103), .b(new_n106), .c(new_n109), .o1(new_n110));
  tech160nm_fioai012aa1n04x5   g015(.a(new_n105), .b(new_n107), .c(new_n104), .o1(new_n111));
  tech160nm_finor002aa1n05x5   g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand02aa1d16x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n16x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nanp02aa1n12x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n03x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  norp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand42aa1n06x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nor042aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nand42aa1n03x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  nano23aa1n03x5               g025(.a(new_n117), .b(new_n119), .c(new_n120), .d(new_n118), .out0(new_n121));
  nanp02aa1n03x5               g026(.a(new_n121), .b(new_n116), .o1(new_n122));
  norb02aa1n06x5               g027(.a(new_n115), .b(new_n114), .out0(new_n123));
  oaih22aa1n06x5               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  aoi022aa1d24x5               g029(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  ao0012aa1n03x7               g030(.a(new_n112), .b(new_n114), .c(new_n113), .o(new_n126));
  aoi013aa1n09x5               g031(.a(new_n126), .b(new_n123), .c(new_n124), .d(new_n125), .o1(new_n127));
  aoai13aa1n12x5               g032(.a(new_n127), .b(new_n122), .c(new_n110), .d(new_n111), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[9] ), .b(\b[8] ), .out0(new_n129));
  nanp02aa1n06x5               g034(.a(new_n128), .b(new_n129), .o1(new_n130));
  xorc02aa1n12x5               g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n130), .c(new_n98), .out0(\s[10] ));
  oai022aa1d24x5               g037(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n133), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(new_n130), .b(new_n134), .o1(new_n135));
  nand42aa1n10x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nor042aa1d18x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  aoi012aa1d24x5               g042(.a(new_n137), .b(\a[10] ), .c(\b[9] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(new_n138), .b(new_n136), .o1(new_n139));
  nanb02aa1n02x5               g044(.a(new_n139), .b(new_n135), .out0(new_n140));
  norb02aa1n02x5               g045(.a(new_n136), .b(new_n137), .out0(new_n141));
  aoi022aa1n02x5               g046(.a(new_n130), .b(new_n134), .c(\b[9] ), .d(\a[10] ), .o1(new_n142));
  oa0012aa1n03x5               g047(.a(new_n140), .b(new_n142), .c(new_n141), .o(\s[11] ));
  inv000aa1d42x5               g048(.a(new_n137), .o1(new_n144));
  aoai13aa1n02x5               g049(.a(new_n144), .b(new_n139), .c(new_n130), .d(new_n134), .o1(new_n145));
  nor042aa1n06x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n20x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  aoib12aa1n02x5               g053(.a(new_n137), .b(new_n147), .c(new_n146), .out0(new_n149));
  aoi022aa1n02x5               g054(.a(new_n140), .b(new_n149), .c(new_n145), .d(new_n148), .o1(\s[12] ));
  aoi012aa1n02x5               g055(.a(new_n99), .b(new_n101), .c(new_n102), .o1(new_n151));
  nona23aa1n09x5               g056(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n152));
  oai012aa1n06x5               g057(.a(new_n111), .b(new_n152), .c(new_n151), .o1(new_n153));
  nanb02aa1n06x5               g058(.a(new_n122), .b(new_n153), .out0(new_n154));
  nano23aa1d15x5               g059(.a(new_n146), .b(new_n137), .c(new_n147), .d(new_n136), .out0(new_n155));
  nand23aa1d12x5               g060(.a(new_n155), .b(new_n129), .c(new_n131), .o1(new_n156));
  aoi022aa1d24x5               g061(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n157));
  nand23aa1d12x5               g062(.a(new_n138), .b(new_n133), .c(new_n157), .o1(new_n158));
  aoi012aa1d18x5               g063(.a(new_n146), .b(new_n137), .c(new_n147), .o1(new_n159));
  nand22aa1n12x5               g064(.a(new_n158), .b(new_n159), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n03x5               g066(.a(new_n161), .b(new_n156), .c(new_n154), .d(new_n127), .o1(new_n162));
  nor042aa1n04x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanp02aa1n04x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(new_n165));
  inv000aa1d42x5               g070(.a(new_n156), .o1(new_n166));
  aoi112aa1n02x5               g071(.a(new_n165), .b(new_n160), .c(new_n128), .d(new_n166), .o1(new_n167));
  aoi012aa1n02x5               g072(.a(new_n167), .b(new_n162), .c(new_n165), .o1(\s[13] ));
  nor002aa1n06x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand02aa1n08x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  aoai13aa1n03x5               g076(.a(new_n171), .b(new_n163), .c(new_n162), .d(new_n164), .o1(new_n172));
  aoi112aa1n02x5               g077(.a(new_n163), .b(new_n171), .c(new_n162), .d(new_n165), .o1(new_n173));
  norb02aa1n02x7               g078(.a(new_n172), .b(new_n173), .out0(\s[14] ));
  nano23aa1n06x5               g079(.a(new_n163), .b(new_n169), .c(new_n170), .d(new_n164), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n160), .c(new_n128), .d(new_n166), .o1(new_n176));
  aoi012aa1n09x5               g081(.a(new_n169), .b(new_n163), .c(new_n170), .o1(new_n177));
  nor042aa1d18x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nand42aa1n06x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  norb02aa1n12x5               g084(.a(new_n179), .b(new_n178), .out0(new_n180));
  xnbna2aa1n03x5               g085(.a(new_n180), .b(new_n176), .c(new_n177), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(new_n177), .o1(new_n182));
  aoai13aa1n03x5               g087(.a(new_n180), .b(new_n182), .c(new_n162), .d(new_n175), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n178), .o1(new_n184));
  inv000aa1d42x5               g089(.a(new_n180), .o1(new_n185));
  aoai13aa1n03x5               g090(.a(new_n184), .b(new_n185), .c(new_n176), .d(new_n177), .o1(new_n186));
  nor002aa1n06x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nand42aa1n03x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  norb02aa1n06x4               g093(.a(new_n188), .b(new_n187), .out0(new_n189));
  aoib12aa1n02x5               g094(.a(new_n178), .b(new_n188), .c(new_n187), .out0(new_n190));
  aoi022aa1n03x5               g095(.a(new_n186), .b(new_n189), .c(new_n183), .d(new_n190), .o1(\s[16] ));
  nona23aa1n09x5               g096(.a(new_n170), .b(new_n164), .c(new_n163), .d(new_n169), .out0(new_n192));
  nano22aa1n12x5               g097(.a(new_n192), .b(new_n180), .c(new_n189), .out0(new_n193));
  nanb02aa1n06x5               g098(.a(new_n156), .b(new_n193), .out0(new_n194));
  aoai13aa1n06x5               g099(.a(new_n179), .b(new_n169), .c(new_n163), .d(new_n170), .o1(new_n195));
  aoi022aa1n02x5               g100(.a(new_n195), .b(new_n184), .c(\a[16] ), .d(\b[15] ), .o1(new_n196));
  aoi112aa1n03x5               g101(.a(new_n196), .b(new_n187), .c(new_n193), .d(new_n160), .o1(new_n197));
  aoai13aa1n12x5               g102(.a(new_n197), .b(new_n194), .c(new_n154), .d(new_n127), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g104(.a(\a[17] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(\b[16] ), .b(new_n200), .out0(new_n201));
  nano32aa1n09x5               g106(.a(new_n156), .b(new_n189), .c(new_n175), .d(new_n180), .out0(new_n202));
  nanp02aa1n03x5               g107(.a(new_n193), .b(new_n160), .o1(new_n203));
  nona22aa1n06x5               g108(.a(new_n203), .b(new_n196), .c(new_n187), .out0(new_n204));
  xorc02aa1n02x5               g109(.a(\a[17] ), .b(\b[16] ), .out0(new_n205));
  aoai13aa1n03x5               g110(.a(new_n205), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[18] ), .b(\b[17] ), .out0(new_n207));
  xnbna2aa1n03x5               g112(.a(new_n207), .b(new_n206), .c(new_n201), .out0(\s[18] ));
  inv000aa1d42x5               g113(.a(\a[18] ), .o1(new_n209));
  xroi22aa1d04x5               g114(.a(new_n200), .b(\b[16] ), .c(new_n209), .d(\b[17] ), .out0(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n211));
  nor042aa1n03x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  aoi112aa1n09x5               g117(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n213));
  nor042aa1n04x5               g118(.a(new_n213), .b(new_n212), .o1(new_n214));
  xorc02aa1n12x5               g119(.a(\a[19] ), .b(\b[18] ), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n211), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g122(.a(new_n214), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n215), .b(new_n218), .c(new_n198), .d(new_n210), .o1(new_n219));
  nor042aa1d18x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  inv040aa1n02x5               g125(.a(new_n220), .o1(new_n221));
  tech160nm_fixnrc02aa1n05x5   g126(.a(\b[18] ), .b(\a[19] ), .out0(new_n222));
  aoai13aa1n02x5               g127(.a(new_n221), .b(new_n222), .c(new_n211), .d(new_n214), .o1(new_n223));
  tech160nm_fixorc02aa1n04x5   g128(.a(\a[20] ), .b(\b[19] ), .out0(new_n224));
  norp02aa1n02x5               g129(.a(new_n224), .b(new_n220), .o1(new_n225));
  aoi022aa1n02x5               g130(.a(new_n223), .b(new_n224), .c(new_n219), .d(new_n225), .o1(\s[20] ));
  nano32aa1n02x4               g131(.a(new_n222), .b(new_n224), .c(new_n205), .d(new_n207), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n228));
  and002aa1n12x5               g133(.a(\b[19] ), .b(\a[20] ), .o(new_n229));
  oao003aa1n12x5               g134(.a(\a[20] ), .b(\b[19] ), .c(new_n221), .carry(new_n230));
  oai013aa1d12x5               g135(.a(new_n230), .b(new_n214), .c(new_n222), .d(new_n229), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  nor002aa1d32x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  nand02aa1d24x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n02x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  xnbna2aa1n03x5               g140(.a(new_n235), .b(new_n228), .c(new_n232), .out0(\s[21] ));
  aoai13aa1n03x5               g141(.a(new_n235), .b(new_n231), .c(new_n198), .d(new_n227), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n233), .o1(new_n238));
  inv000aa1d42x5               g143(.a(new_n235), .o1(new_n239));
  aoai13aa1n02x5               g144(.a(new_n238), .b(new_n239), .c(new_n228), .d(new_n232), .o1(new_n240));
  nor022aa1n08x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  nand02aa1d28x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n242), .b(new_n241), .out0(new_n243));
  aoib12aa1n02x5               g148(.a(new_n233), .b(new_n242), .c(new_n241), .out0(new_n244));
  aoi022aa1n03x5               g149(.a(new_n240), .b(new_n243), .c(new_n237), .d(new_n244), .o1(\s[22] ));
  norb02aa1n02x5               g150(.a(new_n224), .b(new_n222), .out0(new_n246));
  nano23aa1n06x5               g151(.a(new_n233), .b(new_n241), .c(new_n242), .d(new_n234), .out0(new_n247));
  and003aa1n02x5               g152(.a(new_n246), .b(new_n210), .c(new_n247), .o(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n249));
  aoi012aa1n06x5               g154(.a(new_n241), .b(new_n233), .c(new_n242), .o1(new_n250));
  inv020aa1n03x5               g155(.a(new_n250), .o1(new_n251));
  aoi012aa1n03x5               g156(.a(new_n251), .b(new_n231), .c(new_n247), .o1(new_n252));
  nanp02aa1n02x5               g157(.a(new_n249), .b(new_n252), .o1(new_n253));
  nor042aa1d18x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  nanp02aa1n09x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  norb02aa1n02x5               g160(.a(new_n255), .b(new_n254), .out0(new_n256));
  aoi112aa1n02x5               g161(.a(new_n256), .b(new_n251), .c(new_n231), .d(new_n247), .o1(new_n257));
  aoi022aa1n02x5               g162(.a(new_n253), .b(new_n256), .c(new_n249), .d(new_n257), .o1(\s[23] ));
  inv000aa1n02x5               g163(.a(new_n252), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n256), .b(new_n259), .c(new_n198), .d(new_n248), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n254), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n256), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n261), .b(new_n262), .c(new_n249), .d(new_n252), .o1(new_n263));
  nor042aa1n03x5               g168(.a(\b[23] ), .b(\a[24] ), .o1(new_n264));
  nand02aa1n16x5               g169(.a(\b[23] ), .b(\a[24] ), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n265), .b(new_n264), .out0(new_n266));
  aoib12aa1n02x5               g171(.a(new_n254), .b(new_n265), .c(new_n264), .out0(new_n267));
  aoi022aa1n03x5               g172(.a(new_n263), .b(new_n266), .c(new_n260), .d(new_n267), .o1(\s[24] ));
  nano23aa1n03x7               g173(.a(new_n254), .b(new_n264), .c(new_n265), .d(new_n255), .out0(new_n269));
  nand22aa1n06x5               g174(.a(new_n269), .b(new_n247), .o1(new_n270));
  nano32aa1n02x4               g175(.a(new_n270), .b(new_n210), .c(new_n215), .d(new_n224), .out0(new_n271));
  aoai13aa1n04x5               g176(.a(new_n271), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n272));
  inv030aa1n04x5               g177(.a(new_n229), .o1(new_n273));
  oai112aa1n06x5               g178(.a(new_n215), .b(new_n273), .c(new_n213), .d(new_n212), .o1(new_n274));
  nano22aa1n03x5               g179(.a(new_n254), .b(new_n255), .c(new_n265), .out0(new_n275));
  tech160nm_fiaoi012aa1n03p5x5 g180(.a(new_n264), .b(new_n254), .c(new_n265), .o1(new_n276));
  aobi12aa1n06x5               g181(.a(new_n276), .b(new_n251), .c(new_n275), .out0(new_n277));
  aoai13aa1n12x5               g182(.a(new_n277), .b(new_n270), .c(new_n274), .d(new_n230), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(new_n272), .b(new_n279), .o1(new_n280));
  xorc02aa1n12x5               g185(.a(\a[25] ), .b(\b[24] ), .out0(new_n281));
  inv000aa1d42x5               g186(.a(new_n281), .o1(new_n282));
  oai112aa1n02x5               g187(.a(new_n277), .b(new_n282), .c(new_n232), .d(new_n270), .o1(new_n283));
  aboi22aa1n03x5               g188(.a(new_n283), .b(new_n272), .c(new_n280), .d(new_n281), .out0(\s[25] ));
  aoai13aa1n03x5               g189(.a(new_n281), .b(new_n278), .c(new_n198), .d(new_n271), .o1(new_n285));
  nor042aa1n03x5               g190(.a(\b[24] ), .b(\a[25] ), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n286), .o1(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n282), .c(new_n272), .d(new_n279), .o1(new_n288));
  tech160nm_fixorc02aa1n02p5x5 g193(.a(\a[26] ), .b(\b[25] ), .out0(new_n289));
  norp02aa1n02x5               g194(.a(new_n289), .b(new_n286), .o1(new_n290));
  aoi022aa1n03x5               g195(.a(new_n288), .b(new_n289), .c(new_n285), .d(new_n290), .o1(\s[26] ));
  and002aa1n12x5               g196(.a(new_n289), .b(new_n281), .o(new_n292));
  nano32aa1n03x7               g197(.a(new_n270), .b(new_n292), .c(new_n246), .d(new_n210), .out0(new_n293));
  aoai13aa1n06x5               g198(.a(new_n293), .b(new_n204), .c(new_n128), .d(new_n202), .o1(new_n294));
  oao003aa1n02x5               g199(.a(\a[26] ), .b(\b[25] ), .c(new_n287), .carry(new_n295));
  aobi12aa1n12x5               g200(.a(new_n295), .b(new_n278), .c(new_n292), .out0(new_n296));
  xorc02aa1n12x5               g201(.a(\a[27] ), .b(\b[26] ), .out0(new_n297));
  xnbna2aa1n03x5               g202(.a(new_n297), .b(new_n294), .c(new_n296), .out0(\s[27] ));
  aob012aa1n06x5               g203(.a(new_n295), .b(new_n278), .c(new_n292), .out0(new_n299));
  aoai13aa1n02x7               g204(.a(new_n297), .b(new_n299), .c(new_n198), .d(new_n293), .o1(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  inv000aa1n03x5               g206(.a(new_n301), .o1(new_n302));
  inv000aa1n02x5               g207(.a(new_n297), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n302), .b(new_n303), .c(new_n294), .d(new_n296), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[28] ), .b(\b[27] ), .out0(new_n305));
  norp02aa1n02x5               g210(.a(new_n305), .b(new_n301), .o1(new_n306));
  aoi022aa1n03x5               g211(.a(new_n304), .b(new_n305), .c(new_n300), .d(new_n306), .o1(\s[28] ));
  and002aa1n02x5               g212(.a(new_n305), .b(new_n297), .o(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n299), .c(new_n198), .d(new_n293), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n308), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[28] ), .b(\b[27] ), .c(new_n302), .carry(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n310), .c(new_n294), .d(new_n296), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n311), .b(new_n313), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[29] ));
  xorb03aa1n02x5               g220(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n09x5               g221(.a(new_n303), .b(new_n305), .c(new_n313), .out0(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n299), .c(new_n198), .d(new_n293), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n317), .o1(new_n319));
  oaoi03aa1n02x5               g224(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .o1(new_n320));
  inv000aa1n03x5               g225(.a(new_n320), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n319), .c(new_n294), .d(new_n296), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(\b[28] ), .b(\a[29] ), .o(new_n324));
  oabi12aa1n02x5               g229(.a(new_n323), .b(\a[29] ), .c(\b[28] ), .out0(new_n325));
  oab012aa1n02x4               g230(.a(new_n325), .b(new_n311), .c(new_n324), .out0(new_n326));
  aoi022aa1n03x5               g231(.a(new_n322), .b(new_n323), .c(new_n318), .d(new_n326), .o1(\s[30] ));
  nano32aa1n06x5               g232(.a(new_n303), .b(new_n323), .c(new_n305), .d(new_n313), .out0(new_n328));
  aoai13aa1n02x7               g233(.a(new_n328), .b(new_n299), .c(new_n198), .d(new_n293), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[31] ), .b(\b[30] ), .out0(new_n330));
  oao003aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .c(new_n321), .carry(new_n331));
  norb02aa1n02x5               g236(.a(new_n331), .b(new_n330), .out0(new_n332));
  inv000aa1d42x5               g237(.a(new_n328), .o1(new_n333));
  aoai13aa1n03x5               g238(.a(new_n331), .b(new_n333), .c(new_n294), .d(new_n296), .o1(new_n334));
  aoi022aa1n03x5               g239(.a(new_n334), .b(new_n330), .c(new_n329), .d(new_n332), .o1(\s[31] ));
  aoi112aa1n02x5               g240(.a(new_n109), .b(new_n99), .c(new_n101), .d(new_n102), .o1(new_n336));
  aoi012aa1n02x5               g241(.a(new_n336), .b(new_n103), .c(new_n109), .o1(\s[3] ));
  aoi112aa1n02x5               g242(.a(new_n107), .b(new_n106), .c(new_n103), .d(new_n108), .o1(new_n338));
  aoib12aa1n02x5               g243(.a(new_n338), .b(new_n153), .c(new_n104), .out0(\s[4] ));
  norb02aa1n02x5               g244(.a(new_n120), .b(new_n119), .out0(new_n340));
  xnbna2aa1n03x5               g245(.a(new_n340), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  aoi012aa1n02x5               g246(.a(new_n119), .b(new_n153), .c(new_n120), .o1(new_n342));
  xnrb03aa1n02x5               g247(.a(new_n342), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g248(.a(new_n124), .b(new_n153), .c(new_n340), .o(new_n344));
  aoai13aa1n02x5               g249(.a(new_n118), .b(new_n124), .c(new_n153), .d(new_n340), .o1(new_n345));
  nano22aa1n02x4               g250(.a(new_n114), .b(new_n115), .c(new_n118), .out0(new_n346));
  aboi22aa1n03x5               g251(.a(new_n123), .b(new_n345), .c(new_n344), .d(new_n346), .out0(\s[7] ));
  norb02aa1n02x5               g252(.a(new_n113), .b(new_n112), .out0(new_n348));
  orn002aa1n02x5               g253(.a(\a[7] ), .b(\b[6] ), .o(new_n349));
  aoai13aa1n02x5               g254(.a(new_n346), .b(new_n124), .c(new_n153), .d(new_n340), .o1(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n348), .b(new_n350), .c(new_n349), .out0(\s[8] ));
  xnbna2aa1n03x5               g256(.a(new_n129), .b(new_n154), .c(new_n127), .out0(\s[9] ));
endmodule


