// Benchmark "adder" written by ABC on Wed Jul 17 23:01:08 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n153, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n342, new_n344, new_n345, new_n347,
    new_n348, new_n350, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nand02aa1n08x5               g006(.a(\b[8] ), .b(\a[9] ), .o1(new_n102));
  nor002aa1d32x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand02aa1d28x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n03x5               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  nand22aa1n12x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nand42aa1d28x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nor042aa1n12x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nona22aa1n03x5               g013(.a(new_n107), .b(new_n108), .c(new_n106), .out0(new_n109));
  nor002aa1d32x5               g014(.a(\b[2] ), .b(\a[3] ), .o1(new_n110));
  nand42aa1n10x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nano22aa1n03x7               g016(.a(new_n110), .b(new_n107), .c(new_n111), .out0(new_n112));
  aoi012aa1d18x5               g017(.a(new_n103), .b(new_n110), .c(new_n104), .o1(new_n113));
  inv000aa1d42x5               g018(.a(new_n113), .o1(new_n114));
  aoi013aa1n06x4               g019(.a(new_n114), .b(new_n112), .c(new_n109), .d(new_n105), .o1(new_n115));
  nor042aa1d18x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand42aa1n16x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nor002aa1d32x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nand42aa1n08x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nano23aa1n09x5               g024(.a(new_n116), .b(new_n118), .c(new_n119), .d(new_n117), .out0(new_n120));
  nor042aa1n09x5               g025(.a(\b[5] ), .b(\a[6] ), .o1(new_n121));
  nand42aa1d28x5               g026(.a(\b[5] ), .b(\a[6] ), .o1(new_n122));
  norb02aa1n03x5               g027(.a(new_n122), .b(new_n121), .out0(new_n123));
  xorc02aa1n12x5               g028(.a(\a[5] ), .b(\b[4] ), .out0(new_n124));
  nand23aa1n03x5               g029(.a(new_n120), .b(new_n123), .c(new_n124), .o1(new_n125));
  orn002aa1n03x5               g030(.a(\a[6] ), .b(\b[5] ), .o(new_n126));
  oai112aa1n03x5               g031(.a(new_n126), .b(new_n122), .c(\b[4] ), .d(\a[5] ), .o1(new_n127));
  oa0012aa1n03x5               g032(.a(new_n117), .b(new_n118), .c(new_n116), .o(new_n128));
  aoi013aa1n06x4               g033(.a(new_n128), .b(new_n120), .c(new_n122), .d(new_n127), .o1(new_n129));
  tech160nm_fioai012aa1n05x5   g034(.a(new_n129), .b(new_n115), .c(new_n125), .o1(new_n130));
  aoai13aa1n02x5               g035(.a(new_n100), .b(new_n101), .c(new_n130), .d(new_n102), .o1(new_n131));
  nanb02aa1n09x5               g036(.a(new_n103), .b(new_n104), .out0(new_n132));
  norb03aa1d15x5               g037(.a(new_n107), .b(new_n106), .c(new_n108), .out0(new_n133));
  nanb03aa1d24x5               g038(.a(new_n110), .b(new_n111), .c(new_n107), .out0(new_n134));
  oai013aa1d12x5               g039(.a(new_n113), .b(new_n133), .c(new_n134), .d(new_n132), .o1(new_n135));
  nona23aa1n09x5               g040(.a(new_n119), .b(new_n117), .c(new_n116), .d(new_n118), .out0(new_n136));
  nano22aa1n03x7               g041(.a(new_n136), .b(new_n124), .c(new_n123), .out0(new_n137));
  inv020aa1n04x5               g042(.a(new_n122), .o1(new_n138));
  inv000aa1d42x5               g043(.a(\a[5] ), .o1(new_n139));
  inv000aa1d42x5               g044(.a(\b[4] ), .o1(new_n140));
  aoi112aa1n06x5               g045(.a(new_n138), .b(new_n121), .c(new_n139), .d(new_n140), .o1(new_n141));
  inv040aa1n03x5               g046(.a(new_n128), .o1(new_n142));
  oai013aa1n03x5               g047(.a(new_n142), .b(new_n136), .c(new_n141), .d(new_n138), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n102), .b(new_n143), .c(new_n135), .d(new_n137), .o1(new_n144));
  nona22aa1n02x4               g049(.a(new_n144), .b(new_n101), .c(new_n100), .out0(new_n145));
  nanp02aa1n02x5               g050(.a(new_n131), .b(new_n145), .o1(\s[10] ));
  aoi022aa1n02x5               g051(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n147));
  oai112aa1n02x5               g052(.a(new_n145), .b(new_n147), .c(\b[10] ), .d(\a[11] ), .o1(new_n148));
  nor002aa1d24x5               g053(.a(\b[10] ), .b(\a[11] ), .o1(new_n149));
  nand42aa1n08x5               g054(.a(\b[10] ), .b(\a[11] ), .o1(new_n150));
  aboi22aa1n03x5               g055(.a(new_n149), .b(new_n150), .c(new_n145), .d(new_n98), .out0(new_n151));
  norb02aa1n02x5               g056(.a(new_n148), .b(new_n151), .out0(\s[11] ));
  aoi012aa1n02x5               g057(.a(new_n149), .b(new_n145), .c(new_n147), .o1(new_n153));
  xnrb03aa1n02x5               g058(.a(new_n153), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor022aa1n16x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand02aa1d28x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  nona23aa1d18x5               g061(.a(new_n156), .b(new_n150), .c(new_n149), .d(new_n155), .out0(new_n157));
  nona23aa1n03x5               g062(.a(new_n102), .b(new_n98), .c(new_n97), .d(new_n101), .out0(new_n158));
  nor042aa1n03x5               g063(.a(new_n158), .b(new_n157), .o1(new_n159));
  oai012aa1d24x5               g064(.a(new_n98), .b(new_n101), .c(new_n97), .o1(new_n160));
  aoi012aa1n06x5               g065(.a(new_n155), .b(new_n149), .c(new_n156), .o1(new_n161));
  oai012aa1n12x5               g066(.a(new_n161), .b(new_n157), .c(new_n160), .o1(new_n162));
  nor042aa1n06x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nand42aa1d28x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanb02aa1n02x5               g069(.a(new_n163), .b(new_n164), .out0(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n162), .c(new_n130), .d(new_n159), .o1(new_n167));
  oai112aa1n02x5               g072(.a(new_n161), .b(new_n165), .c(new_n157), .d(new_n160), .o1(new_n168));
  aoi012aa1n02x5               g073(.a(new_n168), .b(new_n130), .c(new_n159), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n167), .b(new_n169), .out0(\s[13] ));
  nor042aa1n06x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nand42aa1d28x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  obai22aa1n02x7               g077(.a(new_n172), .b(new_n171), .c(\a[13] ), .d(\b[12] ), .out0(new_n173));
  nona23aa1n02x4               g078(.a(new_n172), .b(new_n164), .c(new_n163), .d(new_n171), .out0(new_n174));
  nona32aa1n02x4               g079(.a(new_n130), .b(new_n174), .c(new_n158), .d(new_n157), .out0(new_n175));
  nano23aa1n06x5               g080(.a(new_n163), .b(new_n171), .c(new_n172), .d(new_n164), .out0(new_n176));
  aoi012aa1n02x5               g081(.a(new_n171), .b(new_n163), .c(new_n172), .o1(new_n177));
  inv020aa1n02x5               g082(.a(new_n177), .o1(new_n178));
  aoi012aa1n02x5               g083(.a(new_n178), .b(new_n162), .c(new_n176), .o1(new_n179));
  aoi012aa1n02x5               g084(.a(new_n171), .b(new_n175), .c(new_n179), .o1(new_n180));
  aoib12aa1n02x5               g085(.a(new_n180), .b(new_n167), .c(new_n173), .out0(\s[14] ));
  norp02aa1n12x5               g086(.a(\b[14] ), .b(\a[15] ), .o1(new_n182));
  nand22aa1n04x5               g087(.a(\b[14] ), .b(\a[15] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n175), .c(new_n179), .out0(\s[15] ));
  aob012aa1n02x5               g090(.a(new_n184), .b(new_n175), .c(new_n179), .out0(new_n186));
  nor002aa1d32x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(new_n187), .o1(new_n188));
  nand22aa1n06x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  aoi012aa1n02x5               g094(.a(new_n182), .b(new_n188), .c(new_n189), .o1(new_n190));
  nano23aa1n02x5               g095(.a(new_n97), .b(new_n101), .c(new_n102), .d(new_n98), .out0(new_n191));
  nano23aa1n06x5               g096(.a(new_n182), .b(new_n187), .c(new_n189), .d(new_n183), .out0(new_n192));
  nano32aa1n03x7               g097(.a(new_n157), .b(new_n192), .c(new_n191), .d(new_n176), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n143), .c(new_n135), .d(new_n137), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n192), .b(new_n178), .c(new_n162), .d(new_n176), .o1(new_n195));
  aoi012aa1n09x5               g100(.a(new_n187), .b(new_n182), .c(new_n189), .o1(new_n196));
  nanp03aa1d12x5               g101(.a(new_n194), .b(new_n195), .c(new_n196), .o1(new_n197));
  aoi022aa1n02x5               g102(.a(new_n186), .b(new_n190), .c(new_n188), .d(new_n197), .o1(\s[16] ));
  xorc02aa1n12x5               g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  nano22aa1n02x4               g104(.a(new_n199), .b(new_n195), .c(new_n196), .out0(new_n200));
  aoi022aa1n02x5               g105(.a(new_n200), .b(new_n194), .c(new_n197), .d(new_n199), .o1(\s[17] ));
  nona23aa1n03x5               g106(.a(new_n189), .b(new_n183), .c(new_n182), .d(new_n187), .out0(new_n202));
  nona22aa1n09x5               g107(.a(new_n159), .b(new_n174), .c(new_n202), .out0(new_n203));
  oaoi13aa1n09x5               g108(.a(new_n203), .b(new_n129), .c(new_n115), .d(new_n125), .o1(new_n204));
  nano23aa1n02x4               g109(.a(new_n149), .b(new_n155), .c(new_n156), .d(new_n150), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n160), .o1(new_n206));
  inv030aa1n02x5               g111(.a(new_n161), .o1(new_n207));
  aoai13aa1n03x5               g112(.a(new_n176), .b(new_n207), .c(new_n205), .d(new_n206), .o1(new_n208));
  aoai13aa1n04x5               g113(.a(new_n196), .b(new_n202), .c(new_n208), .d(new_n177), .o1(new_n209));
  nor042aa1n06x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nand02aa1d28x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  obai22aa1n02x7               g116(.a(new_n211), .b(new_n210), .c(\a[17] ), .d(\b[16] ), .out0(new_n212));
  oaoi13aa1n02x5               g117(.a(new_n212), .b(new_n199), .c(new_n209), .d(new_n204), .o1(new_n213));
  nano22aa1n03x7               g118(.a(new_n210), .b(new_n199), .c(new_n211), .out0(new_n214));
  oaih12aa1n02x5               g119(.a(new_n214), .b(new_n209), .c(new_n204), .o1(new_n215));
  nor042aa1n06x5               g120(.a(\b[16] ), .b(\a[17] ), .o1(new_n216));
  tech160nm_fiaoi012aa1n04x5   g121(.a(new_n210), .b(new_n216), .c(new_n211), .o1(new_n217));
  aoi012aa1n02x5               g122(.a(new_n210), .b(new_n215), .c(new_n217), .o1(new_n218));
  norp02aa1n02x5               g123(.a(new_n218), .b(new_n213), .o1(\s[18] ));
  nor002aa1d32x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nand42aa1n06x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n215), .c(new_n217), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g129(.a(new_n220), .o1(new_n225));
  inv000aa1n03x5               g130(.a(new_n217), .o1(new_n226));
  aoai13aa1n06x5               g131(.a(new_n222), .b(new_n226), .c(new_n197), .d(new_n214), .o1(new_n227));
  nor002aa1n16x5               g132(.a(\b[19] ), .b(\a[20] ), .o1(new_n228));
  nand42aa1n06x5               g133(.a(\b[19] ), .b(\a[20] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  norb03aa1n02x5               g135(.a(new_n229), .b(new_n220), .c(new_n228), .out0(new_n231));
  nanp02aa1n03x5               g136(.a(new_n227), .b(new_n231), .o1(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n230), .c(new_n225), .d(new_n227), .o1(\s[20] ));
  nona23aa1n09x5               g138(.a(new_n229), .b(new_n221), .c(new_n220), .d(new_n228), .out0(new_n234));
  nano23aa1n02x4               g139(.a(new_n234), .b(new_n210), .c(new_n199), .d(new_n211), .out0(new_n235));
  oaoi03aa1n09x5               g140(.a(\a[20] ), .b(\b[19] ), .c(new_n225), .o1(new_n236));
  oabi12aa1n06x5               g141(.a(new_n236), .b(new_n234), .c(new_n217), .out0(new_n237));
  nor042aa1n06x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  nanp02aa1n02x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n238), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n237), .c(new_n197), .d(new_n235), .o1(new_n241));
  nano23aa1d15x5               g146(.a(new_n220), .b(new_n228), .c(new_n229), .d(new_n221), .out0(new_n242));
  aoi112aa1n02x5               g147(.a(new_n236), .b(new_n240), .c(new_n242), .d(new_n226), .o1(new_n243));
  aobi12aa1n02x5               g148(.a(new_n243), .b(new_n197), .c(new_n235), .out0(new_n244));
  norb02aa1n03x4               g149(.a(new_n241), .b(new_n244), .out0(\s[21] ));
  inv040aa1n08x5               g150(.a(new_n238), .o1(new_n246));
  xnrc02aa1n12x5               g151(.a(\b[21] ), .b(\a[22] ), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  and002aa1n02x5               g153(.a(\b[21] ), .b(\a[22] ), .o(new_n249));
  oai022aa1n02x5               g154(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n250));
  nona22aa1n03x5               g155(.a(new_n241), .b(new_n249), .c(new_n250), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n248), .c(new_n246), .d(new_n241), .o1(\s[22] ));
  nano22aa1d15x5               g157(.a(new_n247), .b(new_n246), .c(new_n239), .out0(new_n253));
  nand23aa1d12x5               g158(.a(new_n214), .b(new_n253), .c(new_n242), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n253), .b(new_n236), .c(new_n242), .d(new_n226), .o1(new_n256));
  oaoi03aa1n12x5               g161(.a(\a[22] ), .b(\b[21] ), .c(new_n246), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(new_n256), .b(new_n258), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[22] ), .b(\a[23] ), .out0(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n259), .c(new_n197), .d(new_n255), .o1(new_n262));
  aoi112aa1n02x7               g167(.a(new_n261), .b(new_n259), .c(new_n197), .d(new_n255), .o1(new_n263));
  norb02aa1n03x4               g168(.a(new_n262), .b(new_n263), .out0(\s[23] ));
  norp02aa1n02x5               g169(.a(\b[22] ), .b(\a[23] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  xorc02aa1n03x5               g171(.a(\a[24] ), .b(\b[23] ), .out0(new_n267));
  and002aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .o(new_n268));
  oai022aa1n02x5               g173(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n269));
  nona22aa1n03x5               g174(.a(new_n262), .b(new_n268), .c(new_n269), .out0(new_n270));
  aoai13aa1n03x5               g175(.a(new_n270), .b(new_n267), .c(new_n266), .d(new_n262), .o1(\s[24] ));
  norb02aa1n06x4               g176(.a(new_n267), .b(new_n260), .out0(new_n272));
  inv000aa1n02x5               g177(.a(new_n272), .o1(new_n273));
  nano32aa1n02x5               g178(.a(new_n273), .b(new_n214), .c(new_n253), .d(new_n242), .out0(new_n274));
  aob012aa1n02x5               g179(.a(new_n269), .b(\b[23] ), .c(\a[24] ), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n273), .c(new_n256), .d(new_n258), .o1(new_n276));
  xorc02aa1n06x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n276), .c(new_n197), .d(new_n274), .o1(new_n278));
  aoi112aa1n02x7               g183(.a(new_n277), .b(new_n276), .c(new_n197), .d(new_n274), .o1(new_n279));
  norb02aa1n03x4               g184(.a(new_n278), .b(new_n279), .out0(\s[25] ));
  norp02aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n281), .o1(new_n282));
  xorc02aa1n02x5               g187(.a(\a[26] ), .b(\b[25] ), .out0(new_n283));
  and002aa1n02x5               g188(.a(\b[25] ), .b(\a[26] ), .o(new_n284));
  oai022aa1n02x5               g189(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n285));
  nona22aa1n03x5               g190(.a(new_n278), .b(new_n284), .c(new_n285), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n283), .c(new_n282), .d(new_n278), .o1(\s[26] ));
  and002aa1n06x5               g192(.a(new_n283), .b(new_n277), .o(new_n288));
  nano22aa1n12x5               g193(.a(new_n254), .b(new_n288), .c(new_n272), .out0(new_n289));
  tech160nm_fioai012aa1n04x5   g194(.a(new_n289), .b(new_n209), .c(new_n204), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n284), .o1(new_n291));
  aoi022aa1n06x5               g196(.a(new_n276), .b(new_n288), .c(new_n291), .d(new_n285), .o1(new_n292));
  xorc02aa1n12x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  xnbna2aa1n03x5               g198(.a(new_n293), .b(new_n290), .c(new_n292), .out0(\s[27] ));
  inv000aa1d42x5               g199(.a(\a[27] ), .o1(new_n295));
  nanb02aa1n12x5               g200(.a(\b[26] ), .b(new_n295), .out0(new_n296));
  aoai13aa1n06x5               g201(.a(new_n272), .b(new_n257), .c(new_n237), .d(new_n253), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n288), .o1(new_n298));
  aob012aa1n02x5               g203(.a(new_n285), .b(\b[25] ), .c(\a[26] ), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n298), .c(new_n297), .d(new_n275), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n293), .b(new_n300), .c(new_n197), .d(new_n289), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[28] ), .b(\b[27] ), .out0(new_n302));
  oai022aa1n02x5               g207(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n303));
  aoi012aa1n02x5               g208(.a(new_n303), .b(\a[28] ), .c(\b[27] ), .o1(new_n304));
  nand02aa1n02x5               g209(.a(new_n301), .b(new_n304), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n305), .b(new_n302), .c(new_n296), .d(new_n301), .o1(\s[28] ));
  xorc02aa1n12x5               g211(.a(\a[29] ), .b(\b[28] ), .out0(new_n307));
  inv000aa1d42x5               g212(.a(\b[27] ), .o1(new_n308));
  xroi22aa1d04x5               g213(.a(new_n308), .b(\a[28] ), .c(new_n295), .d(\b[26] ), .out0(new_n309));
  aoai13aa1n04x5               g214(.a(new_n309), .b(new_n300), .c(new_n197), .d(new_n289), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n307), .o1(new_n311));
  oaoi03aa1n02x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n296), .o1(new_n312));
  nona22aa1n03x5               g217(.a(new_n310), .b(new_n311), .c(new_n312), .out0(new_n313));
  inv000aa1n06x5               g218(.a(new_n289), .o1(new_n314));
  aoi013aa1n03x5               g219(.a(new_n314), .b(new_n194), .c(new_n195), .d(new_n196), .o1(new_n315));
  oaoi13aa1n03x5               g220(.a(new_n312), .b(new_n309), .c(new_n315), .d(new_n300), .o1(new_n316));
  oai012aa1n03x5               g221(.a(new_n313), .b(new_n316), .c(new_n307), .o1(\s[29] ));
  xorb03aa1n02x5               g222(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g223(.a(new_n311), .b(new_n293), .c(new_n302), .out0(new_n319));
  aob012aa1n02x5               g224(.a(new_n312), .b(\b[28] ), .c(\a[29] ), .out0(new_n320));
  oai012aa1n06x5               g225(.a(new_n320), .b(\b[28] ), .c(\a[29] ), .o1(new_n321));
  oaoi13aa1n03x5               g226(.a(new_n321), .b(new_n319), .c(new_n315), .d(new_n300), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .out0(new_n323));
  inv000aa1n02x5               g228(.a(new_n319), .o1(new_n324));
  norb02aa1n02x5               g229(.a(new_n323), .b(new_n321), .out0(new_n325));
  aoai13aa1n03x5               g230(.a(new_n325), .b(new_n324), .c(new_n290), .d(new_n292), .o1(new_n326));
  oai012aa1n03x5               g231(.a(new_n326), .b(new_n322), .c(new_n323), .o1(\s[30] ));
  xnrc02aa1n02x5               g232(.a(\b[30] ), .b(\a[31] ), .out0(new_n328));
  nano32aa1n02x4               g233(.a(new_n311), .b(new_n323), .c(new_n293), .d(new_n302), .out0(new_n329));
  inv000aa1n02x5               g234(.a(new_n329), .o1(new_n330));
  inv000aa1d42x5               g235(.a(\a[30] ), .o1(new_n331));
  inv000aa1d42x5               g236(.a(\b[29] ), .o1(new_n332));
  oao003aa1n02x5               g237(.a(new_n331), .b(new_n332), .c(new_n321), .carry(new_n333));
  inv000aa1n02x5               g238(.a(new_n333), .o1(new_n334));
  aoai13aa1n06x5               g239(.a(new_n334), .b(new_n330), .c(new_n290), .d(new_n292), .o1(new_n335));
  nanp02aa1n03x5               g240(.a(new_n335), .b(new_n328), .o1(new_n336));
  aoai13aa1n02x7               g241(.a(new_n329), .b(new_n300), .c(new_n197), .d(new_n289), .o1(new_n337));
  nona22aa1n03x5               g242(.a(new_n337), .b(new_n333), .c(new_n328), .out0(new_n338));
  nanp02aa1n03x5               g243(.a(new_n336), .b(new_n338), .o1(\s[31] ));
  norb02aa1n02x5               g244(.a(new_n111), .b(new_n110), .out0(new_n340));
  xobna2aa1n03x5               g245(.a(new_n340), .b(new_n109), .c(new_n107), .out0(\s[3] ));
  oabi12aa1n02x5               g246(.a(new_n110), .b(new_n133), .c(new_n134), .out0(new_n342));
  xorb03aa1n02x5               g247(.a(new_n342), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  nanp03aa1n02x5               g248(.a(new_n112), .b(new_n109), .c(new_n105), .o1(new_n344));
  aoi112aa1n02x5               g249(.a(new_n124), .b(new_n103), .c(new_n104), .d(new_n110), .o1(new_n345));
  aoi022aa1n02x5               g250(.a(new_n135), .b(new_n124), .c(new_n344), .d(new_n345), .o1(\s[5] ));
  oaoi03aa1n02x5               g251(.a(new_n139), .b(new_n140), .c(new_n135), .o1(new_n347));
  oaib12aa1n02x5               g252(.a(new_n141), .b(new_n115), .c(new_n124), .out0(new_n348));
  oai012aa1n02x5               g253(.a(new_n348), .b(new_n347), .c(new_n123), .o1(\s[6] ));
  aoai13aa1n02x5               g254(.a(new_n122), .b(new_n127), .c(new_n135), .d(new_n124), .o1(new_n350));
  xnrb03aa1n02x5               g255(.a(new_n350), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g256(.a(\a[7] ), .b(\b[6] ), .c(new_n350), .o1(new_n352));
  xorb03aa1n02x5               g257(.a(new_n352), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g258(.a(new_n130), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


