// Benchmark "adder" written by ABC on Wed Jul 17 18:19:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n293, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n311, new_n313, new_n314, new_n317, new_n319, new_n321;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n16x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nand02aa1d08x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nor022aa1n16x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nanp02aa1n06x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nano23aa1d15x5               g005(.a(new_n97), .b(new_n99), .c(new_n100), .d(new_n98), .out0(new_n101));
  oai022aa1n04x5               g006(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n102));
  inv030aa1n02x5               g007(.a(new_n102), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand02aa1d08x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  norb02aa1n06x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor002aa1n03x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  aoi022aa1d24x5               g012(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n108));
  oai012aa1n06x5               g013(.a(new_n106), .b(new_n108), .c(new_n107), .o1(new_n109));
  nanp02aa1n09x5               g014(.a(new_n109), .b(new_n103), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  inv040aa1d32x5               g016(.a(\a[6] ), .o1(new_n112));
  inv040aa1d28x5               g017(.a(\b[5] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(new_n113), .b(new_n112), .o1(new_n114));
  nand02aa1n03x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand22aa1n03x5               g020(.a(new_n114), .b(new_n115), .o1(new_n116));
  nor002aa1d32x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  tech160nm_finand02aa1n05x5   g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nano23aa1n06x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .d(new_n111), .out0(new_n119));
  nona23aa1d18x5               g024(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n120));
  oaoi03aa1n02x5               g025(.a(new_n112), .b(new_n113), .c(new_n117), .o1(new_n121));
  tech160nm_fiaoi012aa1n04x5   g026(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n122));
  oai012aa1n04x7               g027(.a(new_n122), .b(new_n120), .c(new_n121), .o1(new_n123));
  aoi013aa1n09x5               g028(.a(new_n123), .b(new_n110), .c(new_n119), .d(new_n101), .o1(new_n124));
  oaoi03aa1n09x5               g029(.a(\a[9] ), .b(\b[8] ), .c(new_n124), .o1(new_n125));
  xorb03aa1n02x5               g030(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  xorc02aa1n12x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  inv000aa1d42x5               g032(.a(\a[10] ), .o1(new_n128));
  inv000aa1d42x5               g033(.a(\b[9] ), .o1(new_n129));
  oai022aa1d18x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  oa0012aa1n02x5               g035(.a(new_n130), .b(new_n129), .c(new_n128), .o(new_n131));
  xnrc02aa1n12x5               g036(.a(\b[10] ), .b(\a[11] ), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n132), .b(new_n131), .c(new_n125), .d(new_n127), .o1(new_n133));
  aoi112aa1n06x5               g038(.a(new_n132), .b(new_n131), .c(new_n125), .d(new_n127), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(\s[11] ));
  and002aa1n02x5               g040(.a(\b[10] ), .b(\a[11] ), .o(new_n136));
  xorc02aa1n12x5               g041(.a(\a[12] ), .b(\b[11] ), .out0(new_n137));
  orn003aa1n03x7               g042(.a(new_n134), .b(new_n136), .c(new_n137), .o(new_n138));
  tech160nm_fioai012aa1n04x5   g043(.a(new_n137), .b(new_n134), .c(new_n136), .o1(new_n139));
  nanp02aa1n03x5               g044(.a(new_n138), .b(new_n139), .o1(\s[12] ));
  xnrc02aa1n02x5               g045(.a(\b[8] ), .b(\a[9] ), .out0(new_n141));
  nona23aa1n09x5               g046(.a(new_n137), .b(new_n127), .c(new_n141), .d(new_n132), .out0(new_n142));
  nanp02aa1n02x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n02x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  oai112aa1n06x5               g049(.a(new_n130), .b(new_n144), .c(new_n129), .d(new_n128), .o1(new_n145));
  oai122aa1n12x5               g050(.a(new_n145), .b(\a[12] ), .c(\b[11] ), .d(\a[11] ), .e(\b[10] ), .o1(new_n146));
  nanp02aa1n09x5               g051(.a(new_n146), .b(new_n143), .o1(new_n147));
  oai012aa1n12x5               g052(.a(new_n147), .b(new_n124), .c(new_n142), .o1(new_n148));
  xorb03aa1n02x5               g053(.a(new_n148), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nand02aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  tech160nm_fiaoi012aa1n05x5   g056(.a(new_n150), .b(new_n148), .c(new_n151), .o1(new_n152));
  xnrb03aa1n03x5               g057(.a(new_n152), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nand02aa1n06x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nano23aa1n09x5               g060(.a(new_n150), .b(new_n154), .c(new_n155), .d(new_n151), .out0(new_n156));
  oa0012aa1n02x5               g061(.a(new_n155), .b(new_n154), .c(new_n150), .o(new_n157));
  xorc02aa1n12x5               g062(.a(\a[15] ), .b(\b[14] ), .out0(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n157), .c(new_n148), .d(new_n156), .o1(new_n159));
  aoi112aa1n02x5               g064(.a(new_n158), .b(new_n157), .c(new_n148), .d(new_n156), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n159), .b(new_n160), .out0(\s[15] ));
  inv000aa1d42x5               g066(.a(\a[15] ), .o1(new_n162));
  inv000aa1d42x5               g067(.a(\b[14] ), .o1(new_n163));
  nanp02aa1n02x5               g068(.a(new_n163), .b(new_n162), .o1(new_n164));
  xnrc02aa1n12x5               g069(.a(\b[15] ), .b(\a[16] ), .out0(new_n165));
  nand23aa1n03x5               g070(.a(new_n159), .b(new_n164), .c(new_n165), .o1(new_n166));
  aoi012aa1n03x5               g071(.a(new_n165), .b(new_n159), .c(new_n164), .o1(new_n167));
  norb02aa1n03x4               g072(.a(new_n166), .b(new_n167), .out0(\s[16] ));
  norb02aa1n02x5               g073(.a(new_n137), .b(new_n141), .out0(new_n169));
  inv000aa1d42x5               g074(.a(\b[10] ), .o1(new_n170));
  xroi22aa1d04x5               g075(.a(new_n128), .b(\b[9] ), .c(new_n170), .d(\a[11] ), .out0(new_n171));
  nona23aa1n09x5               g076(.a(new_n155), .b(new_n151), .c(new_n150), .d(new_n154), .out0(new_n172));
  norb03aa1n12x5               g077(.a(new_n158), .b(new_n172), .c(new_n165), .out0(new_n173));
  nand23aa1n03x5               g078(.a(new_n173), .b(new_n169), .c(new_n171), .o1(new_n174));
  orn002aa1n02x5               g079(.a(\a[16] ), .b(\b[15] ), .o(new_n175));
  and002aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o(new_n176));
  oai122aa1n06x5               g081(.a(new_n155), .b(new_n154), .c(new_n150), .d(new_n163), .e(new_n162), .o1(new_n177));
  aoai13aa1n03x5               g082(.a(new_n175), .b(new_n176), .c(new_n177), .d(new_n164), .o1(new_n178));
  aoi013aa1n09x5               g083(.a(new_n178), .b(new_n173), .c(new_n146), .d(new_n143), .o1(new_n179));
  tech160nm_fioai012aa1n05x5   g084(.a(new_n179), .b(new_n124), .c(new_n174), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(\b[16] ), .o1(new_n183));
  oaoi03aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n180), .o1(new_n184));
  xnrb03aa1n03x5               g089(.a(new_n184), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  oaoi13aa1n09x5               g090(.a(new_n102), .b(new_n106), .c(new_n108), .d(new_n107), .o1(new_n186));
  norb02aa1n03x5               g091(.a(new_n118), .b(new_n117), .out0(new_n187));
  nanb03aa1n09x5               g092(.a(new_n116), .b(new_n187), .c(new_n111), .out0(new_n188));
  inv000aa1d42x5               g093(.a(new_n117), .o1(new_n189));
  oaoi03aa1n02x5               g094(.a(\a[6] ), .b(\b[5] ), .c(new_n189), .o1(new_n190));
  aobi12aa1n06x5               g095(.a(new_n122), .b(new_n101), .c(new_n190), .out0(new_n191));
  oai013aa1n09x5               g096(.a(new_n191), .b(new_n188), .c(new_n186), .d(new_n120), .o1(new_n192));
  nanb03aa1n06x5               g097(.a(new_n165), .b(new_n156), .c(new_n158), .out0(new_n193));
  nor042aa1n03x5               g098(.a(new_n142), .b(new_n193), .o1(new_n194));
  nand02aa1d06x5               g099(.a(new_n192), .b(new_n194), .o1(new_n195));
  nand42aa1n03x5               g100(.a(new_n183), .b(new_n182), .o1(new_n196));
  nand42aa1n03x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  nor002aa1d32x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nand42aa1n08x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nano32aa1d12x5               g104(.a(new_n198), .b(new_n196), .c(new_n199), .d(new_n197), .out0(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n199), .b(new_n198), .c(new_n182), .d(new_n183), .o1(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n201), .c(new_n195), .d(new_n179), .o1(new_n203));
  xorb03aa1n02x5               g108(.a(new_n203), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g109(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  nand02aa1d10x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nor042aa1n06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1n10x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi112aa1n03x5               g115(.a(new_n206), .b(new_n210), .c(new_n203), .d(new_n207), .o1(new_n211));
  aoai13aa1n03x5               g116(.a(new_n210), .b(new_n206), .c(new_n203), .d(new_n207), .o1(new_n212));
  norb02aa1n02x7               g117(.a(new_n212), .b(new_n211), .out0(\s[20] ));
  nano23aa1n09x5               g118(.a(new_n206), .b(new_n208), .c(new_n209), .d(new_n207), .out0(new_n214));
  nand02aa1d04x5               g119(.a(new_n200), .b(new_n214), .o1(new_n215));
  nona23aa1d18x5               g120(.a(new_n209), .b(new_n207), .c(new_n206), .d(new_n208), .out0(new_n216));
  aoi012aa1n12x5               g121(.a(new_n208), .b(new_n206), .c(new_n209), .o1(new_n217));
  oai012aa1n18x5               g122(.a(new_n217), .b(new_n216), .c(new_n202), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoai13aa1n04x5               g124(.a(new_n219), .b(new_n215), .c(new_n195), .d(new_n179), .o1(new_n220));
  xorb03aa1n02x5               g125(.a(new_n220), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  xorc02aa1n02x5               g127(.a(\a[21] ), .b(\b[20] ), .out0(new_n223));
  xorc02aa1n02x5               g128(.a(\a[22] ), .b(\b[21] ), .out0(new_n224));
  aoi112aa1n02x7               g129(.a(new_n222), .b(new_n224), .c(new_n220), .d(new_n223), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n224), .b(new_n222), .c(new_n220), .d(new_n223), .o1(new_n226));
  norb02aa1n03x4               g131(.a(new_n226), .b(new_n225), .out0(\s[22] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  inv040aa1d32x5               g133(.a(\a[22] ), .o1(new_n229));
  xroi22aa1d06x4               g134(.a(new_n228), .b(\b[20] ), .c(new_n229), .d(\b[21] ), .out0(new_n230));
  nand23aa1n03x5               g135(.a(new_n230), .b(new_n200), .c(new_n214), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\b[21] ), .o1(new_n232));
  oaoi03aa1n09x5               g137(.a(new_n229), .b(new_n232), .c(new_n222), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  aoi012aa1n02x5               g139(.a(new_n234), .b(new_n218), .c(new_n230), .o1(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n231), .c(new_n195), .d(new_n179), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g142(.a(\b[22] ), .b(\a[23] ), .o1(new_n238));
  tech160nm_fixorc02aa1n02p5x5 g143(.a(\a[23] ), .b(\b[22] ), .out0(new_n239));
  tech160nm_fixorc02aa1n02p5x5 g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  aoi112aa1n02x7               g145(.a(new_n238), .b(new_n240), .c(new_n236), .d(new_n239), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n240), .b(new_n238), .c(new_n236), .d(new_n239), .o1(new_n242));
  norb02aa1n03x4               g147(.a(new_n242), .b(new_n241), .out0(\s[24] ));
  and002aa1n06x5               g148(.a(new_n240), .b(new_n239), .o(new_n244));
  inv000aa1n02x5               g149(.a(new_n244), .o1(new_n245));
  nor042aa1n02x5               g150(.a(new_n231), .b(new_n245), .o1(new_n246));
  inv030aa1n03x5               g151(.a(new_n202), .o1(new_n247));
  inv000aa1n04x5               g152(.a(new_n217), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n230), .b(new_n248), .c(new_n214), .d(new_n247), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n250));
  oab012aa1n02x4               g155(.a(new_n250), .b(\a[24] ), .c(\b[23] ), .out0(new_n251));
  aoai13aa1n04x5               g156(.a(new_n251), .b(new_n245), .c(new_n249), .d(new_n233), .o1(new_n252));
  aoi012aa1n03x5               g157(.a(new_n252), .b(new_n180), .c(new_n246), .o1(new_n253));
  xnrc02aa1n12x5               g158(.a(\b[24] ), .b(\a[25] ), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  xnrc02aa1n03x5               g160(.a(new_n253), .b(new_n255), .out0(\s[25] ));
  nor042aa1n03x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n03x5               g163(.a(new_n255), .b(new_n252), .c(new_n180), .d(new_n246), .o1(new_n259));
  tech160nm_fixnrc02aa1n05x5   g164(.a(\b[25] ), .b(\a[26] ), .out0(new_n260));
  nand23aa1n03x5               g165(.a(new_n259), .b(new_n258), .c(new_n260), .o1(new_n261));
  aoi012aa1n02x7               g166(.a(new_n260), .b(new_n259), .c(new_n258), .o1(new_n262));
  norb02aa1n03x4               g167(.a(new_n261), .b(new_n262), .out0(\s[26] ));
  oabi12aa1n03x5               g168(.a(new_n178), .b(new_n147), .c(new_n193), .out0(new_n264));
  nor042aa1n03x5               g169(.a(new_n260), .b(new_n254), .o1(new_n265));
  nano22aa1n06x5               g170(.a(new_n231), .b(new_n244), .c(new_n265), .out0(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n264), .c(new_n192), .d(new_n194), .o1(new_n267));
  oao003aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .c(new_n258), .carry(new_n268));
  aobi12aa1n06x5               g173(.a(new_n268), .b(new_n252), .c(new_n265), .out0(new_n269));
  xorc02aa1n12x5               g174(.a(\a[27] ), .b(\b[26] ), .out0(new_n270));
  xnbna2aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n267), .out0(\s[27] ));
  norp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  inv040aa1n03x5               g177(.a(new_n272), .o1(new_n273));
  aobi12aa1n06x5               g178(.a(new_n270), .b(new_n269), .c(new_n267), .out0(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[27] ), .b(\a[28] ), .out0(new_n275));
  nano22aa1n02x4               g180(.a(new_n274), .b(new_n273), .c(new_n275), .out0(new_n276));
  inv040aa1n03x5               g181(.a(new_n265), .o1(new_n277));
  nona23aa1n09x5               g182(.a(new_n230), .b(new_n244), .c(new_n215), .d(new_n277), .out0(new_n278));
  oaoi13aa1n09x5               g183(.a(new_n278), .b(new_n179), .c(new_n124), .d(new_n174), .o1(new_n279));
  aoai13aa1n06x5               g184(.a(new_n244), .b(new_n234), .c(new_n218), .d(new_n230), .o1(new_n280));
  aoai13aa1n04x5               g185(.a(new_n268), .b(new_n277), .c(new_n280), .d(new_n251), .o1(new_n281));
  oaih12aa1n02x5               g186(.a(new_n270), .b(new_n281), .c(new_n279), .o1(new_n282));
  tech160nm_fiaoi012aa1n02p5x5 g187(.a(new_n275), .b(new_n282), .c(new_n273), .o1(new_n283));
  norp02aa1n03x5               g188(.a(new_n283), .b(new_n276), .o1(\s[28] ));
  xnrc02aa1n02x5               g189(.a(\b[28] ), .b(\a[29] ), .out0(new_n285));
  norb02aa1n02x5               g190(.a(new_n270), .b(new_n275), .out0(new_n286));
  oaih12aa1n02x5               g191(.a(new_n286), .b(new_n281), .c(new_n279), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[28] ), .b(\b[27] ), .c(new_n273), .carry(new_n288));
  tech160nm_fiaoi012aa1n02p5x5 g193(.a(new_n285), .b(new_n287), .c(new_n288), .o1(new_n289));
  aobi12aa1n02x7               g194(.a(new_n286), .b(new_n269), .c(new_n267), .out0(new_n290));
  nano22aa1n03x5               g195(.a(new_n290), .b(new_n285), .c(new_n288), .out0(new_n291));
  norp02aa1n03x5               g196(.a(new_n289), .b(new_n291), .o1(\s[29] ));
  nanp02aa1n02x5               g197(.a(\b[0] ), .b(\a[1] ), .o1(new_n293));
  xorb03aa1n02x5               g198(.a(new_n293), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  xnrc02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .out0(new_n295));
  norb03aa1n02x5               g200(.a(new_n270), .b(new_n285), .c(new_n275), .out0(new_n296));
  oaih12aa1n02x5               g201(.a(new_n296), .b(new_n281), .c(new_n279), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n288), .carry(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n295), .b(new_n297), .c(new_n298), .o1(new_n299));
  aobi12aa1n02x7               g204(.a(new_n296), .b(new_n269), .c(new_n267), .out0(new_n300));
  nano22aa1n03x5               g205(.a(new_n300), .b(new_n295), .c(new_n298), .out0(new_n301));
  norp02aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[30] ));
  xnrc02aa1n02x5               g207(.a(\b[30] ), .b(\a[31] ), .out0(new_n303));
  norb02aa1n03x4               g208(.a(new_n296), .b(new_n295), .out0(new_n304));
  aobi12aa1n06x5               g209(.a(new_n304), .b(new_n269), .c(new_n267), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n306));
  nano22aa1n03x5               g211(.a(new_n305), .b(new_n303), .c(new_n306), .out0(new_n307));
  oaih12aa1n02x5               g212(.a(new_n304), .b(new_n281), .c(new_n279), .o1(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n303), .b(new_n308), .c(new_n306), .o1(new_n309));
  nor002aa1n02x5               g214(.a(new_n309), .b(new_n307), .o1(\s[31] ));
  norp03aa1n02x5               g215(.a(new_n106), .b(new_n107), .c(new_n108), .o1(new_n311));
  norb02aa1n02x5               g216(.a(new_n109), .b(new_n311), .out0(\s[3] ));
  xorc02aa1n02x5               g217(.a(\a[4] ), .b(\b[3] ), .out0(new_n313));
  norp02aa1n02x5               g218(.a(new_n313), .b(new_n104), .o1(new_n314));
  aoi022aa1n02x5               g219(.a(new_n110), .b(new_n313), .c(new_n109), .d(new_n314), .o1(\s[4] ));
  xobna2aa1n03x5               g220(.a(new_n187), .b(new_n110), .c(new_n111), .out0(\s[5] ));
  nanp03aa1n02x5               g221(.a(new_n110), .b(new_n111), .c(new_n187), .o1(new_n317));
  xobna2aa1n03x5               g222(.a(new_n116), .b(new_n317), .c(new_n189), .out0(\s[6] ));
  oai012aa1n02x5               g223(.a(new_n121), .b(new_n188), .c(new_n186), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g225(.a(new_n99), .b(new_n319), .c(new_n100), .o1(new_n321));
  xnrb03aa1n02x5               g226(.a(new_n321), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g227(.a(new_n192), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


