// Benchmark "adder" written by ABC on Wed Jul 17 19:44:51 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n335, new_n336, new_n338, new_n339,
    new_n340, new_n342, new_n343, new_n345, new_n346, new_n347;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  xnrc02aa1n02x5               g002(.a(\b[2] ), .b(\a[3] ), .out0(new_n98));
  orn002aa1n02x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nanp02aa1n04x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n06x5               g005(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(new_n101));
  nor002aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n04x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor022aa1n06x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb03aa1n12x5               g009(.a(new_n103), .b(new_n102), .c(new_n104), .out0(new_n105));
  aoai13aa1n09x5               g010(.a(new_n105), .b(new_n98), .c(new_n101), .d(new_n99), .o1(new_n106));
  nand42aa1n04x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nor042aa1n04x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand42aa1n02x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nanb03aa1n02x5               g014(.a(new_n108), .b(new_n109), .c(new_n107), .out0(new_n110));
  xnrc02aa1n02x5               g015(.a(\b[7] ), .b(\a[8] ), .out0(new_n111));
  inv000aa1d42x5               g016(.a(\b[4] ), .o1(new_n112));
  nanb02aa1d36x5               g017(.a(\a[5] ), .b(new_n112), .out0(new_n113));
  aoi022aa1n06x5               g018(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n114));
  oai112aa1n03x5               g019(.a(new_n114), .b(new_n113), .c(\b[5] ), .d(\a[6] ), .o1(new_n115));
  nor043aa1n03x5               g020(.a(new_n115), .b(new_n110), .c(new_n111), .o1(new_n116));
  nano22aa1n03x7               g021(.a(new_n108), .b(new_n107), .c(new_n109), .out0(new_n117));
  xorc02aa1n06x5               g022(.a(\a[8] ), .b(\b[7] ), .out0(new_n118));
  nor002aa1n02x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  nanb03aa1n06x5               g024(.a(new_n119), .b(new_n113), .c(new_n107), .out0(new_n120));
  nanp03aa1n02x5               g025(.a(new_n120), .b(new_n117), .c(new_n118), .o1(new_n121));
  inv030aa1n02x5               g026(.a(new_n108), .o1(new_n122));
  tech160nm_fioaoi03aa1n03p5x5 g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  nanb02aa1n06x5               g028(.a(new_n123), .b(new_n121), .out0(new_n124));
  xorc02aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n106), .d(new_n116), .o1(new_n126));
  xorc02aa1n02x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  and002aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  oai022aa1d18x5               g033(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n129));
  nor042aa1n06x5               g034(.a(new_n129), .b(new_n128), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(new_n126), .b(new_n130), .o1(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n127), .c(new_n97), .d(new_n126), .o1(\s[10] ));
  inv000aa1d42x5               g037(.a(new_n129), .o1(new_n133));
  aoi022aa1n09x5               g038(.a(new_n126), .b(new_n133), .c(\b[9] ), .d(\a[10] ), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n06x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  and002aa1n02x5               g041(.a(\b[10] ), .b(\a[11] ), .o(new_n137));
  norp02aa1n02x5               g042(.a(new_n137), .b(new_n136), .o1(new_n138));
  nor042aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n12x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n09x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  aoai13aa1n02x5               g047(.a(new_n142), .b(new_n136), .c(new_n134), .d(new_n138), .o1(new_n143));
  aoi112aa1n03x5               g048(.a(new_n142), .b(new_n136), .c(new_n134), .d(new_n138), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(\s[12] ));
  nanp02aa1n03x5               g050(.a(new_n116), .b(new_n106), .o1(new_n146));
  aoi013aa1n06x4               g051(.a(new_n123), .b(new_n117), .c(new_n120), .d(new_n118), .o1(new_n147));
  and002aa1n02x5               g052(.a(\b[8] ), .b(\a[9] ), .o(new_n148));
  aoi112aa1n03x5               g053(.a(new_n137), .b(new_n136), .c(\a[10] ), .d(\b[9] ), .o1(new_n149));
  nona23aa1n02x4               g054(.a(new_n149), .b(new_n141), .c(new_n148), .d(new_n129), .out0(new_n150));
  aoi022aa1n06x5               g055(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n151));
  nona23aa1n09x5               g056(.a(new_n151), .b(new_n140), .c(new_n136), .d(new_n139), .out0(new_n152));
  tech160nm_fioai012aa1n03p5x5 g057(.a(new_n140), .b(new_n139), .c(new_n136), .o1(new_n153));
  oai012aa1n18x5               g058(.a(new_n153), .b(new_n152), .c(new_n130), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  aoai13aa1n03x5               g060(.a(new_n155), .b(new_n150), .c(new_n146), .d(new_n147), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n02x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand42aa1n03x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  aoi012aa1n03x5               g064(.a(new_n158), .b(new_n156), .c(new_n159), .o1(new_n160));
  xnrb03aa1n03x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  tech160nm_fixorc02aa1n02p5x5 g066(.a(\a[3] ), .b(\b[2] ), .out0(new_n162));
  nand42aa1n02x5               g067(.a(new_n101), .b(new_n99), .o1(new_n163));
  inv040aa1n03x5               g068(.a(new_n105), .o1(new_n164));
  tech160nm_fiaoi012aa1n04x5   g069(.a(new_n164), .b(new_n163), .c(new_n162), .o1(new_n165));
  nanb03aa1n03x5               g070(.a(new_n115), .b(new_n117), .c(new_n118), .out0(new_n166));
  oai012aa1n06x5               g071(.a(new_n147), .b(new_n166), .c(new_n165), .o1(new_n167));
  nor043aa1n02x5               g072(.a(new_n152), .b(new_n129), .c(new_n148), .o1(new_n168));
  nor002aa1n02x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand42aa1n03x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nano23aa1n03x5               g075(.a(new_n158), .b(new_n169), .c(new_n170), .d(new_n159), .out0(new_n171));
  aoai13aa1n06x5               g076(.a(new_n171), .b(new_n154), .c(new_n167), .d(new_n168), .o1(new_n172));
  oai012aa1n06x5               g077(.a(new_n170), .b(new_n169), .c(new_n158), .o1(new_n173));
  norp02aa1n04x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  nand42aa1n02x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n172), .c(new_n173), .out0(\s[15] ));
  nand42aa1n02x5               g082(.a(new_n172), .b(new_n173), .o1(new_n178));
  norp02aa1n04x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand02aa1n03x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  nanb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n174), .c(new_n178), .d(new_n176), .o1(new_n182));
  inv030aa1n02x5               g087(.a(new_n173), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n176), .b(new_n183), .c(new_n156), .d(new_n171), .o1(new_n184));
  nona22aa1n02x4               g089(.a(new_n184), .b(new_n181), .c(new_n174), .out0(new_n185));
  nanp02aa1n02x5               g090(.a(new_n182), .b(new_n185), .o1(\s[16] ));
  norb02aa1n02x5               g091(.a(new_n159), .b(new_n158), .out0(new_n187));
  orn002aa1n02x5               g092(.a(\a[14] ), .b(\b[13] ), .o(new_n188));
  nona23aa1n03x5               g093(.a(new_n180), .b(new_n175), .c(new_n174), .d(new_n179), .out0(new_n189));
  nano32aa1n02x4               g094(.a(new_n189), .b(new_n187), .c(new_n188), .d(new_n170), .out0(new_n190));
  nanp02aa1n02x5               g095(.a(new_n168), .b(new_n190), .o1(new_n191));
  tech160nm_fiao0012aa1n02p5x5 g096(.a(new_n179), .b(new_n174), .c(new_n180), .o(new_n192));
  oabi12aa1n03x5               g097(.a(new_n192), .b(new_n189), .c(new_n173), .out0(new_n193));
  aoi012aa1n06x5               g098(.a(new_n193), .b(new_n154), .c(new_n190), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n191), .c(new_n146), .d(new_n147), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d28x5               g101(.a(\a[17] ), .o1(new_n197));
  inv040aa1d32x5               g102(.a(\b[16] ), .o1(new_n198));
  oaoi03aa1n03x5               g103(.a(new_n197), .b(new_n198), .c(new_n195), .o1(new_n199));
  xnrb03aa1n03x5               g104(.a(new_n199), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nano23aa1n02x4               g105(.a(new_n174), .b(new_n179), .c(new_n180), .d(new_n175), .out0(new_n201));
  nanp02aa1n03x5               g106(.a(new_n201), .b(new_n171), .o1(new_n202));
  nor042aa1n03x5               g107(.a(new_n150), .b(new_n202), .o1(new_n203));
  oai112aa1n02x5               g108(.a(new_n149), .b(new_n141), .c(new_n129), .d(new_n128), .o1(new_n204));
  tech160nm_fiaoi012aa1n02p5x5 g109(.a(new_n192), .b(new_n201), .c(new_n183), .o1(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n202), .c(new_n204), .d(new_n153), .o1(new_n206));
  norp02aa1n02x5               g111(.a(\b[16] ), .b(\a[17] ), .o1(new_n207));
  nand42aa1n03x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  nor002aa1d32x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  nano23aa1n06x5               g115(.a(new_n207), .b(new_n209), .c(new_n210), .d(new_n208), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n206), .c(new_n167), .d(new_n203), .o1(new_n212));
  aoai13aa1n12x5               g117(.a(new_n210), .b(new_n209), .c(new_n197), .d(new_n198), .o1(new_n213));
  xnrc02aa1n12x5               g118(.a(\b[18] ), .b(\a[19] ), .out0(new_n214));
  inv000aa1n04x5               g119(.a(new_n214), .o1(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n212), .c(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand42aa1n02x5               g122(.a(new_n212), .b(new_n213), .o1(new_n218));
  norp02aa1n02x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  xnrc02aa1n12x5               g124(.a(\b[19] ), .b(\a[20] ), .out0(new_n220));
  aoai13aa1n03x5               g125(.a(new_n220), .b(new_n219), .c(new_n218), .d(new_n215), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n213), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n215), .b(new_n222), .c(new_n195), .d(new_n211), .o1(new_n223));
  nona22aa1n02x5               g128(.a(new_n223), .b(new_n220), .c(new_n219), .out0(new_n224));
  nanp02aa1n03x5               g129(.a(new_n221), .b(new_n224), .o1(\s[20] ));
  aoai13aa1n06x5               g130(.a(new_n203), .b(new_n124), .c(new_n106), .d(new_n116), .o1(new_n226));
  norb03aa1d15x5               g131(.a(new_n211), .b(new_n220), .c(new_n214), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  orn002aa1n02x5               g133(.a(\a[19] ), .b(\b[18] ), .o(new_n229));
  oao003aa1n02x5               g134(.a(\a[20] ), .b(\b[19] ), .c(new_n229), .carry(new_n230));
  oai013aa1d12x5               g135(.a(new_n230), .b(new_n214), .c(new_n220), .d(new_n213), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n04x5               g137(.a(new_n232), .b(new_n228), .c(new_n226), .d(new_n194), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nand42aa1n03x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  nanb02aa1n03x5               g141(.a(new_n235), .b(new_n236), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  nor022aa1n08x5               g143(.a(\b[21] ), .b(\a[22] ), .o1(new_n239));
  nand02aa1n04x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nanb02aa1n02x5               g145(.a(new_n239), .b(new_n240), .out0(new_n241));
  aoai13aa1n02x5               g146(.a(new_n241), .b(new_n235), .c(new_n233), .d(new_n238), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n238), .b(new_n231), .c(new_n195), .d(new_n227), .o1(new_n243));
  nona22aa1n02x4               g148(.a(new_n243), .b(new_n241), .c(new_n235), .out0(new_n244));
  nanp02aa1n02x5               g149(.a(new_n242), .b(new_n244), .o1(\s[22] ));
  nano23aa1n09x5               g150(.a(new_n235), .b(new_n239), .c(new_n240), .d(new_n236), .out0(new_n246));
  nona23aa1d18x5               g151(.a(new_n211), .b(new_n246), .c(new_n220), .d(new_n214), .out0(new_n247));
  inv000aa1d42x5               g152(.a(new_n247), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n206), .c(new_n167), .d(new_n203), .o1(new_n249));
  tech160nm_fioai012aa1n04x5   g154(.a(new_n240), .b(new_n239), .c(new_n235), .o1(new_n250));
  inv000aa1n02x5               g155(.a(new_n250), .o1(new_n251));
  aoi012aa1n03x5               g156(.a(new_n251), .b(new_n231), .c(new_n246), .o1(new_n252));
  nor022aa1n08x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  nand42aa1n08x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  xnbna2aa1n03x5               g160(.a(new_n255), .b(new_n249), .c(new_n252), .out0(\s[23] ));
  aoai13aa1n04x5               g161(.a(new_n252), .b(new_n247), .c(new_n226), .d(new_n194), .o1(new_n257));
  nor022aa1n08x5               g162(.a(\b[23] ), .b(\a[24] ), .o1(new_n258));
  nand42aa1n06x5               g163(.a(\b[23] ), .b(\a[24] ), .o1(new_n259));
  nanb02aa1n02x5               g164(.a(new_n258), .b(new_n259), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n253), .c(new_n257), .d(new_n255), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(new_n257), .b(new_n255), .o1(new_n262));
  nona22aa1n02x4               g167(.a(new_n262), .b(new_n260), .c(new_n253), .out0(new_n263));
  nanp02aa1n02x5               g168(.a(new_n263), .b(new_n261), .o1(\s[24] ));
  nona23aa1n02x4               g169(.a(new_n259), .b(new_n254), .c(new_n253), .d(new_n258), .out0(new_n265));
  nor042aa1n03x5               g170(.a(new_n247), .b(new_n265), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n206), .c(new_n167), .d(new_n203), .o1(new_n267));
  nona22aa1n09x5               g172(.a(new_n215), .b(new_n220), .c(new_n213), .out0(new_n268));
  nano23aa1n03x5               g173(.a(new_n253), .b(new_n258), .c(new_n259), .d(new_n254), .out0(new_n269));
  nanp02aa1n02x5               g174(.a(new_n269), .b(new_n246), .o1(new_n270));
  oai012aa1n02x5               g175(.a(new_n259), .b(new_n258), .c(new_n253), .o1(new_n271));
  aobi12aa1n02x5               g176(.a(new_n271), .b(new_n269), .c(new_n251), .out0(new_n272));
  aoai13aa1n12x5               g177(.a(new_n272), .b(new_n270), .c(new_n268), .d(new_n230), .o1(new_n273));
  inv000aa1n02x5               g178(.a(new_n273), .o1(new_n274));
  nanp02aa1n04x5               g179(.a(new_n267), .b(new_n274), .o1(new_n275));
  tech160nm_fixorc02aa1n04x5   g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  nor003aa1n03x5               g181(.a(new_n265), .b(new_n241), .c(new_n237), .o1(new_n277));
  oai012aa1n02x5               g182(.a(new_n271), .b(new_n265), .c(new_n250), .o1(new_n278));
  aoi112aa1n02x5               g183(.a(new_n276), .b(new_n278), .c(new_n231), .d(new_n277), .o1(new_n279));
  aoi022aa1n02x5               g184(.a(new_n275), .b(new_n276), .c(new_n267), .d(new_n279), .o1(\s[25] ));
  norp02aa1n02x5               g185(.a(\b[24] ), .b(\a[25] ), .o1(new_n281));
  xnrc02aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .out0(new_n282));
  aoai13aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n275), .d(new_n276), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n276), .b(new_n273), .c(new_n195), .d(new_n266), .o1(new_n284));
  nona22aa1n03x5               g189(.a(new_n284), .b(new_n282), .c(new_n281), .out0(new_n285));
  nanp02aa1n02x5               g190(.a(new_n283), .b(new_n285), .o1(\s[26] ));
  norb02aa1n02x7               g191(.a(new_n276), .b(new_n282), .out0(new_n287));
  nano22aa1n06x5               g192(.a(new_n247), .b(new_n287), .c(new_n269), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n206), .c(new_n167), .d(new_n203), .o1(new_n289));
  aoi112aa1n02x5               g194(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n290));
  oab012aa1n02x4               g195(.a(new_n290), .b(\a[26] ), .c(\b[25] ), .out0(new_n291));
  aobi12aa1n06x5               g196(.a(new_n291), .b(new_n273), .c(new_n287), .out0(new_n292));
  xorc02aa1n02x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  xnbna2aa1n03x5               g198(.a(new_n293), .b(new_n289), .c(new_n292), .out0(\s[27] ));
  nand42aa1n03x5               g199(.a(new_n289), .b(new_n292), .o1(new_n295));
  norp02aa1n02x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  norp02aa1n02x5               g201(.a(\b[27] ), .b(\a[28] ), .o1(new_n297));
  nanp02aa1n02x5               g202(.a(\b[27] ), .b(\a[28] ), .o1(new_n298));
  norb02aa1n06x4               g203(.a(new_n298), .b(new_n297), .out0(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n296), .c(new_n295), .d(new_n293), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n287), .b(new_n278), .c(new_n231), .d(new_n277), .o1(new_n302));
  nand42aa1n04x5               g207(.a(new_n302), .b(new_n291), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n293), .b(new_n303), .c(new_n195), .d(new_n288), .o1(new_n304));
  nona22aa1n02x5               g209(.a(new_n304), .b(new_n300), .c(new_n296), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n301), .b(new_n305), .o1(\s[28] ));
  norb02aa1n02x5               g211(.a(new_n293), .b(new_n300), .out0(new_n307));
  aoai13aa1n06x5               g212(.a(new_n307), .b(new_n303), .c(new_n195), .d(new_n288), .o1(new_n308));
  oai012aa1n02x5               g213(.a(new_n298), .b(new_n297), .c(new_n296), .o1(new_n309));
  nand42aa1n04x5               g214(.a(new_n308), .b(new_n309), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  norb02aa1n02x5               g216(.a(new_n309), .b(new_n311), .out0(new_n312));
  aoi022aa1n02x7               g217(.a(new_n310), .b(new_n311), .c(new_n308), .d(new_n312), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanp03aa1n02x5               g219(.a(new_n311), .b(new_n293), .c(new_n299), .o1(new_n315));
  nanb02aa1n03x5               g220(.a(new_n315), .b(new_n295), .out0(new_n316));
  oao003aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n309), .carry(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n315), .c(new_n289), .d(new_n292), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  norp02aa1n02x5               g224(.a(\b[28] ), .b(\a[29] ), .o1(new_n320));
  aoi012aa1n02x5               g225(.a(new_n309), .b(\a[29] ), .c(\b[28] ), .o1(new_n321));
  norp03aa1n02x5               g226(.a(new_n321), .b(new_n319), .c(new_n320), .o1(new_n322));
  aoi022aa1n03x5               g227(.a(new_n322), .b(new_n316), .c(new_n318), .d(new_n319), .o1(\s[30] ));
  norb02aa1n02x5               g228(.a(new_n319), .b(new_n315), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n303), .c(new_n195), .d(new_n288), .o1(new_n325));
  oao003aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n326));
  nanb02aa1n02x5               g231(.a(\b[30] ), .b(\a[31] ), .out0(new_n327));
  nanb02aa1n02x5               g232(.a(\a[31] ), .b(\b[30] ), .out0(new_n328));
  aoi022aa1n03x5               g233(.a(new_n325), .b(new_n326), .c(new_n328), .d(new_n327), .o1(new_n329));
  aobi12aa1n06x5               g234(.a(new_n324), .b(new_n289), .c(new_n292), .out0(new_n330));
  xnrc02aa1n02x5               g235(.a(\b[30] ), .b(\a[31] ), .out0(new_n331));
  nano22aa1n03x5               g236(.a(new_n330), .b(new_n326), .c(new_n331), .out0(new_n332));
  norp02aa1n03x5               g237(.a(new_n329), .b(new_n332), .o1(\s[31] ));
  xnbna2aa1n03x5               g238(.a(new_n162), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  norb02aa1n02x5               g239(.a(new_n103), .b(new_n104), .out0(new_n335));
  aoi012aa1n02x5               g240(.a(new_n102), .b(new_n163), .c(new_n162), .o1(new_n336));
  oai012aa1n02x5               g241(.a(new_n106), .b(new_n336), .c(new_n335), .o1(\s[4] ));
  and002aa1n02x5               g242(.a(new_n114), .b(new_n113), .o(new_n338));
  aoai13aa1n02x5               g243(.a(new_n103), .b(new_n164), .c(new_n163), .d(new_n162), .o1(new_n339));
  xnrc02aa1n02x5               g244(.a(\b[4] ), .b(\a[5] ), .out0(new_n340));
  aoi022aa1n02x5               g245(.a(new_n339), .b(new_n340), .c(new_n338), .d(new_n106), .o1(\s[5] ));
  norb02aa1n02x5               g246(.a(new_n107), .b(new_n119), .out0(new_n342));
  aoai13aa1n02x5               g247(.a(new_n338), .b(new_n164), .c(new_n163), .d(new_n162), .o1(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n342), .b(new_n343), .c(new_n113), .out0(\s[6] ));
  aoai13aa1n02x5               g249(.a(new_n117), .b(new_n120), .c(new_n106), .d(new_n338), .o1(new_n345));
  nanb02aa1n02x5               g250(.a(new_n120), .b(new_n343), .out0(new_n346));
  aoi022aa1n02x5               g251(.a(new_n346), .b(new_n107), .c(new_n122), .d(new_n109), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n345), .b(new_n347), .out0(\s[7] ));
  xnbna2aa1n03x5               g253(.a(new_n118), .b(new_n345), .c(new_n122), .out0(\s[8] ));
  xnbna2aa1n03x5               g254(.a(new_n125), .b(new_n146), .c(new_n147), .out0(\s[9] ));
endmodule


