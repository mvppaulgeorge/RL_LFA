// Benchmark "adder" written by ABC on Thu Jul 18 05:16:41 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n311, new_n313, new_n314, new_n315, new_n317, new_n318,
    new_n320, new_n321, new_n323, new_n324, new_n326;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[9] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[8] ), .o1(new_n99));
  orn002aa1n06x5               g004(.a(\a[2] ), .b(\b[1] ), .o(new_n100));
  nand22aa1n03x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n12x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  aob012aa1n06x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  xorc02aa1n12x5               g008(.a(\a[3] ), .b(\b[2] ), .out0(new_n104));
  oai022aa1n02x5               g009(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n105));
  aoi012aa1n06x5               g010(.a(new_n105), .b(new_n103), .c(new_n104), .o1(new_n106));
  nor042aa1n09x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand02aa1n16x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nand42aa1n16x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nano22aa1n03x7               g014(.a(new_n107), .b(new_n108), .c(new_n109), .out0(new_n110));
  nand22aa1n04x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  nor002aa1d24x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nand02aa1n04x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nano22aa1n03x7               g018(.a(new_n112), .b(new_n111), .c(new_n113), .out0(new_n114));
  nor042aa1n09x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand22aa1n09x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nor002aa1d32x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  norb03aa1n03x5               g022(.a(new_n116), .b(new_n115), .c(new_n117), .out0(new_n118));
  nand23aa1n03x5               g023(.a(new_n114), .b(new_n110), .c(new_n118), .o1(new_n119));
  nano23aa1n09x5               g024(.a(new_n115), .b(new_n107), .c(new_n108), .d(new_n109), .out0(new_n120));
  inv030aa1n02x5               g025(.a(new_n116), .o1(new_n121));
  oab012aa1n03x5               g026(.a(new_n121), .b(new_n112), .c(new_n117), .out0(new_n122));
  norb03aa1n12x5               g027(.a(new_n108), .b(new_n107), .c(new_n115), .out0(new_n123));
  aboi22aa1n09x5               g028(.a(new_n123), .b(new_n108), .c(new_n120), .d(new_n122), .out0(new_n124));
  oai012aa1n18x5               g029(.a(new_n124), .b(new_n106), .c(new_n119), .o1(new_n125));
  oaoi03aa1n02x5               g030(.a(new_n98), .b(new_n99), .c(new_n125), .o1(new_n126));
  xorb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  nand42aa1n08x5               g032(.a(\b[10] ), .b(\a[11] ), .o1(new_n128));
  nor002aa1n12x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  norb02aa1n02x5               g034(.a(new_n128), .b(new_n129), .out0(new_n130));
  oaib12aa1n06x5               g035(.a(new_n125), .b(new_n99), .c(\a[9] ), .out0(new_n131));
  oai022aa1d18x5               g036(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n132));
  aboi22aa1n03x5               g037(.a(new_n132), .b(new_n131), .c(\b[9] ), .d(\a[10] ), .out0(new_n133));
  inv000aa1d42x5               g038(.a(new_n129), .o1(new_n134));
  nanb02aa1n02x5               g039(.a(new_n132), .b(new_n131), .out0(new_n135));
  aoi022aa1d24x5               g040(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n136));
  nanp03aa1n03x5               g041(.a(new_n135), .b(new_n134), .c(new_n136), .o1(new_n137));
  oa0012aa1n02x5               g042(.a(new_n137), .b(new_n133), .c(new_n130), .o(\s[11] ));
  norp02aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand02aa1d20x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  oai022aa1n04x5               g046(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n142));
  nanb03aa1n02x5               g047(.a(new_n142), .b(new_n137), .c(new_n140), .out0(new_n143));
  aoai13aa1n02x5               g048(.a(new_n143), .b(new_n141), .c(new_n134), .d(new_n137), .o1(\s[12] ));
  nor002aa1n02x5               g049(.a(\b[1] ), .b(\a[2] ), .o1(new_n145));
  aoi012aa1n02x5               g050(.a(new_n145), .b(new_n101), .c(new_n102), .o1(new_n146));
  xnrc02aa1n02x5               g051(.a(\b[2] ), .b(\a[3] ), .out0(new_n147));
  oabi12aa1n02x7               g052(.a(new_n105), .b(new_n147), .c(new_n146), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n112), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n117), .o1(new_n150));
  oai112aa1n02x5               g055(.a(new_n150), .b(new_n116), .c(\b[7] ), .d(\a[8] ), .o1(new_n151));
  nano32aa1n03x7               g056(.a(new_n151), .b(new_n113), .c(new_n149), .d(new_n111), .out0(new_n152));
  nanp03aa1n03x5               g057(.a(new_n148), .b(new_n152), .c(new_n110), .o1(new_n153));
  xorc02aa1n02x5               g058(.a(\a[10] ), .b(\b[9] ), .out0(new_n154));
  nano23aa1n03x5               g059(.a(new_n139), .b(new_n129), .c(new_n140), .d(new_n128), .out0(new_n155));
  xorc02aa1n02x5               g060(.a(\a[9] ), .b(\b[8] ), .out0(new_n156));
  nand23aa1n03x5               g061(.a(new_n155), .b(new_n154), .c(new_n156), .o1(new_n157));
  aoai13aa1n04x5               g062(.a(new_n140), .b(new_n142), .c(new_n132), .d(new_n136), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n158), .b(new_n157), .c(new_n153), .d(new_n124), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nand42aa1n08x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nanp03aa1n02x5               g068(.a(new_n159), .b(new_n162), .c(new_n163), .o1(new_n164));
  nor022aa1n08x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand42aa1n16x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  oai022aa1n02x5               g072(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n168));
  nanb03aa1n02x5               g073(.a(new_n168), .b(new_n164), .c(new_n166), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n167), .c(new_n164), .d(new_n162), .o1(\s[14] ));
  nano23aa1n06x5               g075(.a(new_n161), .b(new_n165), .c(new_n166), .d(new_n163), .out0(new_n171));
  aoi022aa1n06x5               g076(.a(new_n159), .b(new_n171), .c(new_n166), .d(new_n168), .o1(new_n172));
  inv040aa1d28x5               g077(.a(\a[15] ), .o1(new_n173));
  inv040aa1d30x5               g078(.a(\b[14] ), .o1(new_n174));
  nand02aa1d06x5               g079(.a(new_n174), .b(new_n173), .o1(new_n175));
  nand02aa1n03x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n172), .b(new_n176), .c(new_n175), .out0(\s[15] ));
  nanp02aa1n02x5               g082(.a(new_n175), .b(new_n176), .o1(new_n178));
  tech160nm_fixnrc02aa1n02p5x5 g083(.a(\b[15] ), .b(\a[16] ), .out0(new_n179));
  oaoi13aa1n02x7               g084(.a(new_n179), .b(new_n175), .c(new_n172), .d(new_n178), .o1(new_n180));
  nor042aa1n03x5               g085(.a(new_n172), .b(new_n178), .o1(new_n181));
  nano22aa1n02x4               g086(.a(new_n181), .b(new_n175), .c(new_n179), .out0(new_n182));
  norp02aa1n03x5               g087(.a(new_n180), .b(new_n182), .o1(\s[16] ));
  inv040aa1d32x5               g088(.a(\a[17] ), .o1(new_n184));
  nona22aa1n09x5               g089(.a(new_n171), .b(new_n179), .c(new_n178), .out0(new_n185));
  nor042aa1n06x5               g090(.a(new_n185), .b(new_n157), .o1(new_n186));
  tech160nm_fioai012aa1n03p5x5 g091(.a(new_n166), .b(new_n165), .c(new_n161), .o1(new_n187));
  orn002aa1n02x5               g092(.a(\a[16] ), .b(\b[15] ), .o(new_n188));
  aob012aa1n02x5               g093(.a(new_n176), .b(\b[15] ), .c(\a[16] ), .out0(new_n189));
  aoai13aa1n03x5               g094(.a(new_n188), .b(new_n189), .c(new_n187), .d(new_n175), .o1(new_n190));
  oabi12aa1n12x5               g095(.a(new_n190), .b(new_n185), .c(new_n158), .out0(new_n191));
  aoi012aa1n02x5               g096(.a(new_n191), .b(new_n125), .c(new_n186), .o1(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[16] ), .c(new_n184), .out0(\s[17] ));
  oaoi03aa1n03x5               g098(.a(\a[17] ), .b(\b[16] ), .c(new_n192), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  inv040aa1d32x5               g100(.a(\a[18] ), .o1(new_n196));
  xroi22aa1d06x4               g101(.a(new_n184), .b(\b[16] ), .c(new_n196), .d(\b[17] ), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n191), .c(new_n125), .d(new_n186), .o1(new_n198));
  nanb02aa1n06x5               g103(.a(\b[16] ), .b(new_n184), .out0(new_n199));
  oaoi03aa1n12x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n199), .o1(new_n200));
  inv000aa1n03x5               g105(.a(new_n200), .o1(new_n201));
  nor042aa1d18x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nand42aa1d28x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n198), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n02x5               g111(.a(new_n202), .o1(new_n207));
  aob012aa1n03x5               g112(.a(new_n204), .b(new_n198), .c(new_n201), .out0(new_n208));
  nor042aa1n09x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  norb03aa1n02x5               g116(.a(new_n210), .b(new_n202), .c(new_n209), .out0(new_n212));
  nand42aa1n02x5               g117(.a(new_n208), .b(new_n212), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n211), .c(new_n207), .d(new_n208), .o1(\s[20] ));
  nano23aa1n09x5               g119(.a(new_n202), .b(new_n209), .c(new_n210), .d(new_n203), .out0(new_n215));
  nand02aa1d04x5               g120(.a(new_n197), .b(new_n215), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n06x5               g122(.a(new_n217), .b(new_n191), .c(new_n125), .d(new_n186), .o1(new_n218));
  nona23aa1n09x5               g123(.a(new_n210), .b(new_n203), .c(new_n202), .d(new_n209), .out0(new_n219));
  oaoi03aa1n09x5               g124(.a(\a[20] ), .b(\b[19] ), .c(new_n207), .o1(new_n220));
  oabi12aa1n12x5               g125(.a(new_n220), .b(new_n201), .c(new_n219), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  xnrc02aa1n12x5               g127(.a(\b[20] ), .b(\a[21] ), .out0(new_n223));
  xobna2aa1n03x5               g128(.a(new_n223), .b(new_n218), .c(new_n222), .out0(\s[21] ));
  tech160nm_fiaoi012aa1n05x5   g129(.a(new_n223), .b(new_n218), .c(new_n222), .o1(new_n225));
  xnrc02aa1n06x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  norp02aa1n02x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  norp02aa1n03x5               g132(.a(new_n225), .b(new_n227), .o1(new_n228));
  nanp02aa1n02x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  oai022aa1n02x5               g134(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n230));
  nanb02aa1n02x5               g135(.a(new_n230), .b(new_n229), .out0(new_n231));
  obai22aa1n03x5               g136(.a(new_n226), .b(new_n228), .c(new_n225), .d(new_n231), .out0(\s[22] ));
  nor042aa1n06x5               g137(.a(new_n226), .b(new_n223), .o1(new_n233));
  and003aa1n02x5               g138(.a(new_n197), .b(new_n233), .c(new_n215), .o(new_n234));
  aoai13aa1n06x5               g139(.a(new_n234), .b(new_n191), .c(new_n125), .d(new_n186), .o1(new_n235));
  aoi022aa1n06x5               g140(.a(new_n221), .b(new_n233), .c(new_n229), .d(new_n230), .o1(new_n236));
  xorc02aa1n02x5               g141(.a(\a[23] ), .b(\b[22] ), .out0(new_n237));
  xnbna2aa1n03x5               g142(.a(new_n237), .b(new_n235), .c(new_n236), .out0(\s[23] ));
  nor042aa1n12x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  aob012aa1n03x5               g145(.a(new_n237), .b(new_n235), .c(new_n236), .out0(new_n241));
  xorc02aa1n02x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  nanp02aa1n04x5               g147(.a(\b[23] ), .b(\a[24] ), .o1(new_n243));
  oai022aa1n02x5               g148(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n243), .b(new_n244), .out0(new_n245));
  nanp02aa1n06x5               g150(.a(new_n241), .b(new_n245), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n246), .b(new_n242), .c(new_n240), .d(new_n241), .o1(\s[24] ));
  nanp02aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  nor042aa1n02x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  nano23aa1n03x7               g154(.a(new_n239), .b(new_n249), .c(new_n243), .d(new_n248), .out0(new_n250));
  nano22aa1n02x4               g155(.a(new_n216), .b(new_n233), .c(new_n250), .out0(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n191), .c(new_n125), .d(new_n186), .o1(new_n252));
  aoai13aa1n06x5               g157(.a(new_n233), .b(new_n220), .c(new_n215), .d(new_n200), .o1(new_n253));
  nand02aa1d04x5               g158(.a(new_n230), .b(new_n229), .o1(new_n254));
  inv000aa1n02x5               g159(.a(new_n250), .o1(new_n255));
  tech160nm_fioai012aa1n04x5   g160(.a(new_n243), .b(new_n249), .c(new_n239), .o1(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n255), .c(new_n253), .d(new_n254), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[25] ), .b(\b[24] ), .out0(new_n259));
  xnbna2aa1n03x5               g164(.a(new_n259), .b(new_n252), .c(new_n258), .out0(\s[25] ));
  norp02aa1n02x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  aob012aa1n03x5               g167(.a(new_n259), .b(new_n252), .c(new_n258), .out0(new_n263));
  tech160nm_fixorc02aa1n03p5x5 g168(.a(\a[26] ), .b(\b[25] ), .out0(new_n264));
  nanp02aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .o1(new_n265));
  oai022aa1n02x5               g170(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n266));
  norb02aa1n02x5               g171(.a(new_n265), .b(new_n266), .out0(new_n267));
  nand42aa1n02x5               g172(.a(new_n263), .b(new_n267), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n264), .c(new_n263), .d(new_n262), .o1(\s[26] ));
  and002aa1n02x5               g174(.a(new_n264), .b(new_n259), .o(new_n270));
  nano32aa1n03x7               g175(.a(new_n216), .b(new_n270), .c(new_n233), .d(new_n250), .out0(new_n271));
  aoai13aa1n12x5               g176(.a(new_n271), .b(new_n191), .c(new_n125), .d(new_n186), .o1(new_n272));
  aoi022aa1n12x5               g177(.a(new_n257), .b(new_n270), .c(new_n265), .d(new_n266), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n272), .out0(\s[27] ));
  nand42aa1n04x5               g180(.a(new_n257), .b(new_n270), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(new_n266), .b(new_n265), .o1(new_n277));
  nanp03aa1n06x5               g182(.a(new_n276), .b(new_n272), .c(new_n277), .o1(new_n278));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  xnrc02aa1n12x5               g184(.a(\b[27] ), .b(\a[28] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n279), .c(new_n278), .d(new_n274), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n274), .o1(new_n282));
  norp02aa1n02x5               g187(.a(new_n280), .b(new_n279), .o1(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n282), .c(new_n273), .d(new_n272), .o1(new_n284));
  nanp02aa1n03x5               g189(.a(new_n281), .b(new_n284), .o1(\s[28] ));
  norb02aa1n15x5               g190(.a(new_n274), .b(new_n280), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n278), .b(new_n286), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n286), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[27] ), .b(\a[28] ), .o1(new_n289));
  oai012aa1n02x5               g194(.a(new_n289), .b(new_n280), .c(new_n279), .o1(new_n290));
  aoai13aa1n03x5               g195(.a(new_n290), .b(new_n288), .c(new_n273), .d(new_n272), .o1(new_n291));
  xorc02aa1n02x5               g196(.a(\a[29] ), .b(\b[28] ), .out0(new_n292));
  oaoi13aa1n02x5               g197(.a(new_n292), .b(new_n289), .c(new_n280), .d(new_n279), .o1(new_n293));
  aoi022aa1n03x5               g198(.a(new_n291), .b(new_n292), .c(new_n287), .d(new_n293), .o1(\s[29] ));
  xorb03aa1n02x5               g199(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g200(.a(new_n280), .b(new_n274), .c(new_n292), .out0(new_n296));
  nanp02aa1n02x5               g201(.a(new_n278), .b(new_n296), .o1(new_n297));
  inv000aa1n02x5               g202(.a(new_n296), .o1(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n298), .c(new_n273), .d(new_n272), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  norb02aa1n02x5               g206(.a(new_n299), .b(new_n301), .out0(new_n302));
  aoi022aa1n03x5               g207(.a(new_n300), .b(new_n301), .c(new_n297), .d(new_n302), .o1(\s[30] ));
  nanp03aa1n02x5               g208(.a(new_n286), .b(new_n292), .c(new_n301), .o1(new_n304));
  nanb02aa1n03x5               g209(.a(new_n304), .b(new_n278), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n304), .c(new_n273), .d(new_n272), .o1(new_n307));
  xorc02aa1n02x5               g212(.a(\a[31] ), .b(\b[30] ), .out0(new_n308));
  norb02aa1n02x5               g213(.a(new_n306), .b(new_n308), .out0(new_n309));
  aoi022aa1n03x5               g214(.a(new_n307), .b(new_n308), .c(new_n305), .d(new_n309), .o1(\s[31] ));
  inv000aa1d42x5               g215(.a(\a[3] ), .o1(new_n311));
  xorb03aa1n02x5               g216(.a(new_n146), .b(\b[2] ), .c(new_n311), .out0(\s[3] ));
  nanp02aa1n02x5               g217(.a(new_n103), .b(new_n104), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[4] ), .b(\b[3] ), .out0(new_n314));
  aoib12aa1n02x5               g219(.a(new_n314), .b(new_n311), .c(\b[2] ), .out0(new_n315));
  aoi022aa1n02x5               g220(.a(new_n148), .b(new_n314), .c(new_n315), .d(new_n313), .o1(\s[4] ));
  aoai13aa1n02x5               g221(.a(new_n114), .b(new_n105), .c(new_n103), .d(new_n104), .o1(new_n317));
  aoi022aa1n02x5               g222(.a(new_n148), .b(new_n111), .c(new_n113), .d(new_n149), .o1(new_n318));
  norb02aa1n02x5               g223(.a(new_n317), .b(new_n318), .out0(\s[5] ));
  aoi012aa1n02x5               g224(.a(new_n112), .b(new_n148), .c(new_n114), .o1(new_n320));
  nona32aa1n02x4               g225(.a(new_n317), .b(new_n117), .c(new_n121), .d(new_n112), .out0(new_n321));
  aoai13aa1n02x5               g226(.a(new_n321), .b(new_n320), .c(new_n116), .d(new_n150), .o1(\s[6] ));
  aboi22aa1n03x5               g227(.a(new_n107), .b(new_n109), .c(new_n321), .d(new_n116), .out0(new_n323));
  nano32aa1n02x4               g228(.a(new_n107), .b(new_n321), .c(new_n109), .d(new_n116), .out0(new_n324));
  norp02aa1n02x5               g229(.a(new_n324), .b(new_n323), .o1(\s[7] ));
  obai22aa1n02x7               g230(.a(new_n108), .b(new_n115), .c(new_n324), .d(new_n107), .out0(new_n326));
  oaib12aa1n02x5               g231(.a(new_n326), .b(new_n324), .c(new_n123), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


