// Benchmark "adder" written by ABC on Wed Jul 17 16:43:44 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n341, new_n343, new_n346, new_n347,
    new_n350, new_n351, new_n352, new_n354, new_n355;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[2] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[1] ), .o1(new_n98));
  nanp02aa1n04x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand42aa1d28x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand42aa1d28x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  aob012aa1n03x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  xorc02aa1n12x5               g007(.a(\a[4] ), .b(\b[3] ), .out0(new_n103));
  xorc02aa1n12x5               g008(.a(\a[3] ), .b(\b[2] ), .out0(new_n104));
  nand03aa1n04x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor042aa1n04x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  inv040aa1n03x5               g011(.a(new_n106), .o1(new_n107));
  oao003aa1n02x5               g012(.a(\a[4] ), .b(\b[3] ), .c(new_n107), .carry(new_n108));
  nand22aa1n04x5               g013(.a(new_n105), .b(new_n108), .o1(new_n109));
  nand02aa1n03x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  norp02aa1n09x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  norb02aa1n09x5               g016(.a(new_n110), .b(new_n111), .out0(new_n112));
  xnrc02aa1n12x5               g017(.a(\b[4] ), .b(\a[5] ), .out0(new_n113));
  inv000aa1n02x5               g018(.a(new_n113), .o1(new_n114));
  xorc02aa1n12x5               g019(.a(\a[8] ), .b(\b[7] ), .out0(new_n115));
  xorc02aa1n12x5               g020(.a(\a[7] ), .b(\b[6] ), .out0(new_n116));
  nanp02aa1n02x5               g021(.a(new_n116), .b(new_n115), .o1(new_n117));
  nano22aa1n03x7               g022(.a(new_n117), .b(new_n114), .c(new_n112), .out0(new_n118));
  inv040aa1n02x5               g023(.a(new_n111), .o1(new_n119));
  nor042aa1n02x5               g024(.a(\b[4] ), .b(\a[5] ), .o1(new_n120));
  aob012aa1n06x5               g025(.a(new_n119), .b(new_n120), .c(new_n110), .out0(new_n121));
  inv000aa1d42x5               g026(.a(\a[8] ), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\b[7] ), .o1(new_n123));
  nor042aa1n06x5               g028(.a(\b[6] ), .b(\a[7] ), .o1(new_n124));
  oaoi03aa1n09x5               g029(.a(new_n122), .b(new_n123), .c(new_n124), .o1(new_n125));
  inv000aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  aoi013aa1n06x4               g031(.a(new_n126), .b(new_n121), .c(new_n116), .d(new_n115), .o1(new_n127));
  inv020aa1n03x5               g032(.a(new_n127), .o1(new_n128));
  xnrc02aa1n12x5               g033(.a(\b[8] ), .b(\a[9] ), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n129), .o1(new_n130));
  aoai13aa1n06x5               g035(.a(new_n130), .b(new_n128), .c(new_n109), .d(new_n118), .o1(new_n131));
  xorc02aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .out0(new_n132));
  oaoi13aa1n02x5               g037(.a(new_n132), .b(new_n131), .c(\a[9] ), .d(\b[8] ), .o1(new_n133));
  nand22aa1n03x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  oa0022aa1n06x5               g039(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n135));
  nanp03aa1n02x5               g040(.a(new_n131), .b(new_n134), .c(new_n135), .o1(new_n136));
  nanb02aa1n03x5               g041(.a(new_n133), .b(new_n136), .out0(\s[10] ));
  nanp02aa1n02x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nor042aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nanb03aa1n02x5               g044(.a(new_n139), .b(new_n134), .c(new_n138), .out0(new_n140));
  ao0012aa1n03x7               g045(.a(new_n140), .b(new_n131), .c(new_n135), .o(new_n141));
  nanb02aa1n06x5               g046(.a(new_n139), .b(new_n138), .out0(new_n142));
  aob012aa1n02x5               g047(.a(new_n134), .b(new_n131), .c(new_n135), .out0(new_n143));
  aobi12aa1n02x5               g048(.a(new_n141), .b(new_n143), .c(new_n142), .out0(\s[11] ));
  nor042aa1n04x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  and002aa1n12x5               g050(.a(\b[11] ), .b(\a[12] ), .o(new_n146));
  nor042aa1n02x5               g051(.a(new_n146), .b(new_n145), .o1(new_n147));
  oab012aa1n02x4               g052(.a(new_n139), .b(new_n146), .c(new_n145), .out0(new_n148));
  inv000aa1n02x5               g053(.a(new_n139), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n140), .c(new_n131), .d(new_n135), .o1(new_n150));
  aoi022aa1n02x5               g055(.a(new_n141), .b(new_n148), .c(new_n150), .d(new_n147), .o1(\s[12] ));
  nona23aa1d18x5               g056(.a(new_n147), .b(new_n132), .c(new_n129), .d(new_n142), .out0(new_n152));
  inv040aa1n02x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n03x5               g058(.a(new_n153), .b(new_n128), .c(new_n109), .d(new_n118), .o1(new_n154));
  aoi112aa1n06x5               g059(.a(new_n146), .b(new_n145), .c(\a[11] ), .d(\b[10] ), .o1(new_n155));
  nona23aa1n12x5               g060(.a(new_n155), .b(new_n134), .c(new_n135), .d(new_n139), .out0(new_n156));
  oab012aa1n06x5               g061(.a(new_n145), .b(new_n149), .c(new_n146), .out0(new_n157));
  nanp02aa1n04x5               g062(.a(new_n156), .b(new_n157), .o1(new_n158));
  nanb02aa1n02x5               g063(.a(new_n158), .b(new_n154), .out0(new_n159));
  xorc02aa1n02x5               g064(.a(\a[13] ), .b(\b[12] ), .out0(new_n160));
  nano22aa1n02x4               g065(.a(new_n160), .b(new_n156), .c(new_n157), .out0(new_n161));
  aoi022aa1n02x5               g066(.a(new_n159), .b(new_n160), .c(new_n154), .d(new_n161), .o1(\s[13] ));
  inv040aa1d32x5               g067(.a(\a[13] ), .o1(new_n163));
  nanb02aa1d24x5               g068(.a(\b[12] ), .b(new_n163), .out0(new_n164));
  xnrc02aa1n02x5               g069(.a(\b[6] ), .b(\a[7] ), .out0(new_n165));
  nona23aa1n09x5               g070(.a(new_n115), .b(new_n112), .c(new_n165), .d(new_n113), .out0(new_n166));
  aoai13aa1n09x5               g071(.a(new_n127), .b(new_n166), .c(new_n105), .d(new_n108), .o1(new_n167));
  aoai13aa1n03x5               g072(.a(new_n160), .b(new_n158), .c(new_n167), .d(new_n153), .o1(new_n168));
  xorc02aa1n02x5               g073(.a(\a[14] ), .b(\b[13] ), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n168), .c(new_n164), .out0(\s[14] ));
  inv040aa1d32x5               g075(.a(\a[14] ), .o1(new_n171));
  xroi22aa1d06x4               g076(.a(new_n163), .b(\b[12] ), .c(new_n171), .d(\b[13] ), .out0(new_n172));
  aoai13aa1n03x5               g077(.a(new_n172), .b(new_n158), .c(new_n167), .d(new_n153), .o1(new_n173));
  oaoi03aa1n12x5               g078(.a(\a[14] ), .b(\b[13] ), .c(new_n164), .o1(new_n174));
  inv000aa1d42x5               g079(.a(new_n174), .o1(new_n175));
  xorc02aa1n12x5               g080(.a(\a[15] ), .b(\b[14] ), .out0(new_n176));
  xnbna2aa1n03x5               g081(.a(new_n176), .b(new_n173), .c(new_n175), .out0(\s[15] ));
  aoai13aa1n02x5               g082(.a(new_n176), .b(new_n174), .c(new_n159), .d(new_n172), .o1(new_n178));
  xorc02aa1n02x5               g083(.a(\a[16] ), .b(\b[15] ), .out0(new_n179));
  nor042aa1n06x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  norp02aa1n02x5               g085(.a(new_n179), .b(new_n180), .o1(new_n181));
  inv040aa1n03x5               g086(.a(new_n180), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n176), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n173), .d(new_n175), .o1(new_n184));
  aoi022aa1n02x7               g089(.a(new_n184), .b(new_n179), .c(new_n178), .d(new_n181), .o1(\s[16] ));
  nanp02aa1n02x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  tech160nm_fixnrc02aa1n02p5x5 g091(.a(\b[15] ), .b(\a[16] ), .out0(new_n187));
  nano22aa1n03x7               g092(.a(new_n187), .b(new_n182), .c(new_n186), .out0(new_n188));
  nano22aa1d15x5               g093(.a(new_n152), .b(new_n172), .c(new_n188), .out0(new_n189));
  aoai13aa1n06x5               g094(.a(new_n189), .b(new_n128), .c(new_n118), .d(new_n109), .o1(new_n190));
  nand22aa1n06x5               g095(.a(new_n172), .b(new_n188), .o1(new_n191));
  inv000aa1n02x5               g096(.a(new_n191), .o1(new_n192));
  nand23aa1n04x5               g097(.a(new_n174), .b(new_n176), .c(new_n179), .o1(new_n193));
  oao003aa1n02x5               g098(.a(\a[16] ), .b(\b[15] ), .c(new_n182), .carry(new_n194));
  nanp02aa1n02x5               g099(.a(new_n193), .b(new_n194), .o1(new_n195));
  aoi012aa1n12x5               g100(.a(new_n195), .b(new_n192), .c(new_n158), .o1(new_n196));
  nanp02aa1n09x5               g101(.a(new_n190), .b(new_n196), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  nanb03aa1n02x5               g103(.a(new_n198), .b(new_n193), .c(new_n194), .out0(new_n199));
  aoi012aa1n02x5               g104(.a(new_n199), .b(new_n192), .c(new_n158), .o1(new_n200));
  aoi022aa1n02x5               g105(.a(new_n197), .b(new_n198), .c(new_n190), .d(new_n200), .o1(\s[17] ));
  inv040aa1d32x5               g106(.a(\a[17] ), .o1(new_n202));
  inv040aa1d28x5               g107(.a(\b[16] ), .o1(new_n203));
  nanp02aa1n02x5               g108(.a(new_n203), .b(new_n202), .o1(new_n204));
  aobi12aa1n06x5               g109(.a(new_n194), .b(new_n188), .c(new_n174), .out0(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n191), .c(new_n156), .d(new_n157), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n198), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n207));
  norp02aa1n06x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nand02aa1d28x5               g113(.a(\b[17] ), .b(\a[18] ), .o1(new_n209));
  norb02aa1n06x4               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  xnbna2aa1n03x5               g115(.a(new_n210), .b(new_n207), .c(new_n204), .out0(\s[18] ));
  and002aa1n02x5               g116(.a(new_n198), .b(new_n210), .o(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n213));
  aoi013aa1n09x5               g118(.a(new_n208), .b(new_n209), .c(new_n202), .d(new_n203), .o1(new_n214));
  nor002aa1d32x5               g119(.a(\b[18] ), .b(\a[19] ), .o1(new_n215));
  nand02aa1d24x5               g120(.a(\b[18] ), .b(\a[19] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n213), .c(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n02x5               g124(.a(\a[18] ), .b(\b[17] ), .c(new_n204), .o1(new_n220));
  aoai13aa1n03x5               g125(.a(new_n217), .b(new_n220), .c(new_n197), .d(new_n212), .o1(new_n221));
  nor002aa1d32x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand02aa1d24x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n02x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  inv000aa1d42x5               g129(.a(\a[19] ), .o1(new_n225));
  inv000aa1d42x5               g130(.a(\b[18] ), .o1(new_n226));
  aboi22aa1n03x5               g131(.a(new_n222), .b(new_n223), .c(new_n225), .d(new_n226), .out0(new_n227));
  inv040aa1n08x5               g132(.a(new_n215), .o1(new_n228));
  inv000aa1n02x5               g133(.a(new_n217), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n228), .b(new_n229), .c(new_n213), .d(new_n214), .o1(new_n230));
  aoi022aa1n03x5               g135(.a(new_n230), .b(new_n224), .c(new_n221), .d(new_n227), .o1(\s[20] ));
  nano23aa1n06x5               g136(.a(new_n215), .b(new_n222), .c(new_n223), .d(new_n216), .out0(new_n232));
  nand23aa1n06x5               g137(.a(new_n232), .b(new_n198), .c(new_n210), .o1(new_n233));
  tech160nm_fiaoi012aa1n03p5x5 g138(.a(new_n233), .b(new_n190), .c(new_n196), .o1(new_n234));
  nona23aa1d18x5               g139(.a(new_n223), .b(new_n216), .c(new_n215), .d(new_n222), .out0(new_n235));
  oaoi03aa1n09x5               g140(.a(\a[20] ), .b(\b[19] ), .c(new_n228), .o1(new_n236));
  inv040aa1n02x5               g141(.a(new_n236), .o1(new_n237));
  oai012aa1d24x5               g142(.a(new_n237), .b(new_n235), .c(new_n214), .o1(new_n238));
  xnrc02aa1n06x5               g143(.a(\b[20] ), .b(\a[21] ), .out0(new_n239));
  oabi12aa1n03x5               g144(.a(new_n239), .b(new_n234), .c(new_n238), .out0(new_n240));
  oai112aa1n02x5               g145(.a(new_n237), .b(new_n239), .c(new_n235), .d(new_n214), .o1(new_n241));
  oa0012aa1n03x5               g146(.a(new_n240), .b(new_n234), .c(new_n241), .o(\s[21] ));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  nor042aa1n06x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n243), .b(new_n245), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n233), .o1(new_n247));
  aoai13aa1n02x5               g152(.a(new_n247), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n238), .o1(new_n249));
  inv000aa1n09x5               g154(.a(new_n245), .o1(new_n250));
  aoai13aa1n02x7               g155(.a(new_n250), .b(new_n239), .c(new_n248), .d(new_n249), .o1(new_n251));
  aoi022aa1n03x5               g156(.a(new_n251), .b(new_n244), .c(new_n240), .d(new_n246), .o1(\s[22] ));
  nor042aa1n06x5               g157(.a(new_n243), .b(new_n239), .o1(new_n253));
  norb02aa1n09x5               g158(.a(new_n253), .b(new_n233), .out0(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n255));
  oaoi03aa1n12x5               g160(.a(\a[22] ), .b(\b[21] ), .c(new_n250), .o1(new_n256));
  aoi012aa1d18x5               g161(.a(new_n256), .b(new_n238), .c(new_n253), .o1(new_n257));
  inv040aa1d30x5               g162(.a(new_n257), .o1(new_n258));
  xorc02aa1n12x5               g163(.a(\a[23] ), .b(\b[22] ), .out0(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n258), .c(new_n197), .d(new_n254), .o1(new_n260));
  aoi112aa1n02x5               g165(.a(new_n259), .b(new_n256), .c(new_n238), .d(new_n253), .o1(new_n261));
  aobi12aa1n02x7               g166(.a(new_n260), .b(new_n261), .c(new_n255), .out0(\s[23] ));
  tech160nm_fixorc02aa1n05x5   g167(.a(\a[24] ), .b(\b[23] ), .out0(new_n263));
  nor042aa1n09x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  norp02aa1n02x5               g169(.a(new_n263), .b(new_n264), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n264), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n259), .o1(new_n267));
  aoai13aa1n02x7               g172(.a(new_n266), .b(new_n267), .c(new_n255), .d(new_n257), .o1(new_n268));
  aoi022aa1n02x7               g173(.a(new_n268), .b(new_n263), .c(new_n260), .d(new_n265), .o1(\s[24] ));
  nano32aa1n03x7               g174(.a(new_n233), .b(new_n263), .c(new_n253), .d(new_n259), .out0(new_n270));
  aoai13aa1n02x5               g175(.a(new_n270), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n253), .b(new_n236), .c(new_n232), .d(new_n220), .o1(new_n272));
  inv000aa1n02x5               g177(.a(new_n256), .o1(new_n273));
  and002aa1n06x5               g178(.a(new_n263), .b(new_n259), .o(new_n274));
  inv030aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[24] ), .b(\b[23] ), .c(new_n266), .carry(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n275), .c(new_n272), .d(new_n273), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n197), .d(new_n270), .o1(new_n279));
  aoai13aa1n04x5               g184(.a(new_n274), .b(new_n256), .c(new_n238), .d(new_n253), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n278), .o1(new_n281));
  and003aa1n02x5               g186(.a(new_n280), .b(new_n281), .c(new_n276), .o(new_n282));
  aobi12aa1n03x7               g187(.a(new_n279), .b(new_n282), .c(new_n271), .out0(\s[25] ));
  xorc02aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .out0(new_n284));
  norp02aa1n02x5               g189(.a(\b[24] ), .b(\a[25] ), .o1(new_n285));
  norp02aa1n02x5               g190(.a(new_n284), .b(new_n285), .o1(new_n286));
  inv000aa1n02x5               g191(.a(new_n277), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  aoai13aa1n02x7               g193(.a(new_n288), .b(new_n281), .c(new_n271), .d(new_n287), .o1(new_n289));
  aoi022aa1n02x7               g194(.a(new_n289), .b(new_n284), .c(new_n279), .d(new_n286), .o1(\s[26] ));
  and002aa1n06x5               g195(.a(new_n284), .b(new_n278), .o(new_n291));
  inv000aa1n03x5               g196(.a(new_n291), .o1(new_n292));
  nano23aa1n06x5               g197(.a(new_n292), .b(new_n233), .c(new_n274), .d(new_n253), .out0(new_n293));
  aoai13aa1n06x5               g198(.a(new_n293), .b(new_n206), .c(new_n167), .d(new_n189), .o1(new_n294));
  nanp02aa1n02x5               g199(.a(\b[25] ), .b(\a[26] ), .o1(new_n295));
  oai022aa1n02x5               g200(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n296));
  nanp02aa1n02x5               g201(.a(new_n296), .b(new_n295), .o1(new_n297));
  aoai13aa1n04x5               g202(.a(new_n297), .b(new_n292), .c(new_n280), .d(new_n276), .o1(new_n298));
  xorc02aa1n12x5               g203(.a(\a[27] ), .b(\b[26] ), .out0(new_n299));
  aoai13aa1n06x5               g204(.a(new_n299), .b(new_n298), .c(new_n197), .d(new_n293), .o1(new_n300));
  aoi122aa1n03x5               g205(.a(new_n299), .b(new_n295), .c(new_n296), .d(new_n277), .e(new_n291), .o1(new_n301));
  aobi12aa1n03x7               g206(.a(new_n300), .b(new_n301), .c(new_n294), .out0(\s[27] ));
  xorc02aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .out0(new_n303));
  nor042aa1n03x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  norp02aa1n02x5               g209(.a(new_n303), .b(new_n304), .o1(new_n305));
  aoi022aa1n02x7               g210(.a(new_n277), .b(new_n291), .c(new_n295), .d(new_n296), .o1(new_n306));
  inv000aa1n06x5               g211(.a(new_n304), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n299), .o1(new_n308));
  aoai13aa1n02x7               g213(.a(new_n307), .b(new_n308), .c(new_n306), .d(new_n294), .o1(new_n309));
  aoi022aa1n02x7               g214(.a(new_n309), .b(new_n303), .c(new_n300), .d(new_n305), .o1(\s[28] ));
  and002aa1n02x5               g215(.a(new_n303), .b(new_n299), .o(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n298), .c(new_n197), .d(new_n293), .o1(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  oaoi03aa1n12x5               g218(.a(\a[28] ), .b(\b[27] ), .c(new_n307), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n306), .d(new_n294), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .out0(new_n317));
  norp02aa1n02x5               g222(.a(new_n314), .b(new_n317), .o1(new_n318));
  aoi022aa1n03x5               g223(.a(new_n316), .b(new_n317), .c(new_n312), .d(new_n318), .o1(\s[29] ));
  xorb03aa1n02x5               g224(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g225(.a(new_n308), .b(new_n303), .c(new_n317), .out0(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n298), .c(new_n197), .d(new_n293), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n321), .o1(new_n323));
  inv000aa1d42x5               g228(.a(\b[28] ), .o1(new_n324));
  oaib12aa1n09x5               g229(.a(new_n314), .b(new_n324), .c(\a[29] ), .out0(new_n325));
  oa0012aa1n02x5               g230(.a(new_n325), .b(\b[28] ), .c(\a[29] ), .o(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n323), .c(new_n306), .d(new_n294), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[30] ), .b(\b[29] ), .out0(new_n328));
  oabi12aa1n02x5               g233(.a(new_n328), .b(\a[29] ), .c(\b[28] ), .out0(new_n329));
  norb02aa1n02x5               g234(.a(new_n325), .b(new_n329), .out0(new_n330));
  aoi022aa1n03x5               g235(.a(new_n327), .b(new_n328), .c(new_n322), .d(new_n330), .o1(\s[30] ));
  nano32aa1n06x5               g236(.a(new_n308), .b(new_n328), .c(new_n303), .d(new_n317), .out0(new_n332));
  aoai13aa1n03x5               g237(.a(new_n332), .b(new_n298), .c(new_n197), .d(new_n293), .o1(new_n333));
  xorc02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  oai122aa1n06x5               g239(.a(new_n325), .b(\a[30] ), .c(\b[29] ), .d(\a[29] ), .e(\b[28] ), .o1(new_n335));
  aob012aa1n02x5               g240(.a(new_n335), .b(\b[29] ), .c(\a[30] ), .out0(new_n336));
  norb02aa1n02x5               g241(.a(new_n336), .b(new_n334), .out0(new_n337));
  inv000aa1d42x5               g242(.a(new_n332), .o1(new_n338));
  aoai13aa1n03x5               g243(.a(new_n336), .b(new_n338), .c(new_n306), .d(new_n294), .o1(new_n339));
  aoi022aa1n03x5               g244(.a(new_n339), .b(new_n334), .c(new_n333), .d(new_n337), .o1(\s[31] ));
  nanp03aa1n02x5               g245(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n341));
  xnbna2aa1n03x5               g246(.a(new_n104), .b(new_n341), .c(new_n99), .out0(\s[3] ));
  nanp02aa1n02x5               g247(.a(new_n102), .b(new_n104), .o1(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n103), .b(new_n343), .c(new_n107), .out0(\s[4] ));
  xnbna2aa1n03x5               g249(.a(new_n114), .b(new_n105), .c(new_n108), .out0(\s[5] ));
  aoai13aa1n03x5               g250(.a(new_n112), .b(new_n120), .c(new_n109), .d(new_n114), .o1(new_n346));
  aoi112aa1n02x5               g251(.a(new_n120), .b(new_n112), .c(new_n109), .d(new_n114), .o1(new_n347));
  norb02aa1n02x5               g252(.a(new_n346), .b(new_n347), .out0(\s[6] ));
  xnbna2aa1n03x5               g253(.a(new_n116), .b(new_n346), .c(new_n119), .out0(\s[7] ));
  aob012aa1n03x5               g254(.a(new_n116), .b(new_n346), .c(new_n119), .out0(new_n350));
  oai012aa1n02x7               g255(.a(new_n350), .b(\b[6] ), .c(\a[7] ), .o1(new_n351));
  norp02aa1n02x5               g256(.a(new_n115), .b(new_n124), .o1(new_n352));
  aoi022aa1n02x5               g257(.a(new_n351), .b(new_n115), .c(new_n350), .d(new_n352), .o1(\s[8] ));
  nanp02aa1n02x5               g258(.a(new_n109), .b(new_n118), .o1(new_n354));
  aoi113aa1n02x5               g259(.a(new_n126), .b(new_n130), .c(new_n121), .d(new_n116), .e(new_n115), .o1(new_n355));
  aoi022aa1n02x5               g260(.a(new_n167), .b(new_n130), .c(new_n354), .d(new_n355), .o1(\s[9] ));
endmodule


