// Benchmark "adder" written by ABC on Wed Jul 17 19:08:30 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n324,
    new_n325, new_n328, new_n330, new_n331, new_n332, new_n333, new_n335;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor022aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  norp02aa1n04x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand22aa1n06x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor022aa1n16x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nand02aa1d04x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nona23aa1d18x5               g007(.a(new_n102), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n103));
  xorc02aa1n02x5               g008(.a(\a[5] ), .b(\b[4] ), .out0(new_n104));
  tech160nm_fixorc02aa1n02p5x5 g009(.a(\a[6] ), .b(\b[5] ), .out0(new_n105));
  nano22aa1n03x7               g010(.a(new_n103), .b(new_n104), .c(new_n105), .out0(new_n106));
  and002aa1n18x5               g011(.a(\b[3] ), .b(\a[4] ), .o(new_n107));
  nor042aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nor043aa1n06x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nanb02aa1n12x5               g016(.a(new_n109), .b(new_n111), .out0(new_n112));
  nor002aa1n03x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand22aa1n09x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  tech160nm_fioai012aa1n05x5   g020(.a(new_n115), .b(new_n113), .c(new_n114), .o1(new_n116));
  oaoi13aa1n12x5               g021(.a(new_n107), .b(new_n110), .c(new_n116), .d(new_n112), .o1(new_n117));
  norp02aa1n24x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nor042aa1n03x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  and002aa1n12x5               g024(.a(\b[5] ), .b(\a[6] ), .o(new_n120));
  oab012aa1n03x5               g025(.a(new_n120), .b(new_n118), .c(new_n119), .out0(new_n121));
  oai012aa1n02x5               g026(.a(new_n100), .b(new_n101), .c(new_n99), .o1(new_n122));
  oaib12aa1n06x5               g027(.a(new_n122), .b(new_n103), .c(new_n121), .out0(new_n123));
  xorc02aa1n03x5               g028(.a(\a[9] ), .b(\b[8] ), .out0(new_n124));
  aoai13aa1n02x5               g029(.a(new_n124), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n125));
  nor002aa1n03x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand42aa1n08x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  norb02aa1n06x4               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n125), .c(new_n98), .out0(\s[10] ));
  inv030aa1n02x5               g034(.a(new_n118), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[4] ), .b(\a[5] ), .o1(new_n131));
  nano23aa1n02x4               g036(.a(new_n120), .b(new_n119), .c(new_n130), .d(new_n131), .out0(new_n132));
  tech160nm_fioai012aa1n05x5   g037(.a(new_n110), .b(new_n116), .c(new_n112), .o1(new_n133));
  nona23aa1n06x5               g038(.a(new_n133), .b(new_n132), .c(new_n103), .d(new_n107), .out0(new_n134));
  nona22aa1n02x4               g039(.a(new_n100), .b(new_n101), .c(new_n99), .out0(new_n135));
  aboi22aa1n06x5               g040(.a(new_n103), .b(new_n121), .c(new_n135), .d(new_n100), .out0(new_n136));
  nanp02aa1n02x5               g041(.a(new_n124), .b(new_n128), .o1(new_n137));
  oai012aa1n18x5               g042(.a(new_n127), .b(new_n126), .c(new_n97), .o1(new_n138));
  aoai13aa1n02x5               g043(.a(new_n138), .b(new_n137), .c(new_n134), .d(new_n136), .o1(new_n139));
  xorb03aa1n02x5               g044(.a(new_n139), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  orn002aa1n02x5               g045(.a(\a[11] ), .b(\b[10] ), .o(new_n141));
  nor002aa1n16x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand42aa1n03x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  norb02aa1n02x5               g048(.a(new_n143), .b(new_n142), .out0(new_n144));
  nanp02aa1n03x5               g049(.a(new_n139), .b(new_n144), .o1(new_n145));
  nor022aa1n16x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nanp02aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1n02x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n145), .c(new_n141), .out0(\s[12] ));
  nona23aa1n03x5               g054(.a(new_n147), .b(new_n143), .c(new_n142), .d(new_n146), .out0(new_n150));
  nano22aa1n03x5               g055(.a(new_n150), .b(new_n124), .c(new_n128), .out0(new_n151));
  aoai13aa1n06x5               g056(.a(new_n151), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n152));
  tech160nm_fioai012aa1n03p5x5 g057(.a(new_n147), .b(new_n146), .c(new_n142), .o1(new_n153));
  tech160nm_fioai012aa1n05x5   g058(.a(new_n153), .b(new_n150), .c(new_n138), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n154), .b(new_n152), .out0(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nanp02aa1n09x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nano22aa1n02x4               g063(.a(new_n157), .b(new_n155), .c(new_n158), .out0(new_n159));
  norp02aa1n12x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nanp02aa1n09x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n163));
  nona22aa1n02x4               g068(.a(new_n161), .b(new_n160), .c(new_n157), .out0(new_n164));
  oai012aa1n03x5               g069(.a(new_n163), .b(new_n159), .c(new_n164), .o1(\s[14] ));
  nona23aa1n09x5               g070(.a(new_n161), .b(new_n158), .c(new_n157), .d(new_n160), .out0(new_n166));
  nano23aa1n03x7               g071(.a(new_n157), .b(new_n160), .c(new_n161), .d(new_n158), .out0(new_n167));
  aoi022aa1n02x5               g072(.a(new_n154), .b(new_n167), .c(new_n161), .d(new_n164), .o1(new_n168));
  tech160nm_fioai012aa1n03p5x5 g073(.a(new_n168), .b(new_n152), .c(new_n166), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanp02aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nanb02aa1n03x5               g077(.a(new_n171), .b(new_n172), .out0(new_n173));
  oaoi13aa1n02x5               g078(.a(new_n173), .b(new_n168), .c(new_n152), .d(new_n166), .o1(new_n174));
  nor042aa1n06x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand42aa1n04x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n03x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n171), .c(new_n169), .d(new_n172), .o1(new_n178));
  norb03aa1n02x5               g083(.a(new_n176), .b(new_n171), .c(new_n175), .out0(new_n179));
  oaib12aa1n03x5               g084(.a(new_n178), .b(new_n174), .c(new_n179), .out0(\s[16] ));
  nor003aa1n03x5               g085(.a(new_n166), .b(new_n173), .c(new_n177), .o1(new_n181));
  nand02aa1n02x5               g086(.a(new_n151), .b(new_n181), .o1(new_n182));
  oaih12aa1n02x5               g087(.a(new_n161), .b(new_n160), .c(new_n157), .o1(new_n183));
  oai012aa1n02x5               g088(.a(new_n176), .b(new_n175), .c(new_n171), .o1(new_n184));
  oai013aa1n03x4               g089(.a(new_n184), .b(new_n183), .c(new_n173), .d(new_n177), .o1(new_n185));
  aoi012aa1n12x5               g090(.a(new_n185), .b(new_n154), .c(new_n181), .o1(new_n186));
  aoai13aa1n09x5               g091(.a(new_n186), .b(new_n182), .c(new_n134), .d(new_n136), .o1(new_n187));
  xorb03aa1n02x5               g092(.a(new_n187), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor002aa1d32x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n189), .o1(new_n190));
  xorc02aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  nanp02aa1n03x5               g096(.a(new_n187), .b(new_n191), .o1(new_n192));
  xnrc02aa1n02x5               g097(.a(\b[17] ), .b(\a[18] ), .out0(new_n193));
  xobna2aa1n03x5               g098(.a(new_n193), .b(new_n192), .c(new_n190), .out0(\s[18] ));
  nano23aa1n02x5               g099(.a(new_n142), .b(new_n146), .c(new_n147), .d(new_n143), .out0(new_n195));
  nano23aa1n02x4               g100(.a(new_n171), .b(new_n175), .c(new_n176), .d(new_n172), .out0(new_n196));
  nano32aa1n03x7               g101(.a(new_n137), .b(new_n196), .c(new_n195), .d(new_n167), .out0(new_n197));
  aoai13aa1n09x5               g102(.a(new_n197), .b(new_n123), .c(new_n117), .d(new_n106), .o1(new_n198));
  inv000aa1d42x5               g103(.a(\a[17] ), .o1(new_n199));
  inv000aa1d42x5               g104(.a(\a[18] ), .o1(new_n200));
  xroi22aa1d06x4               g105(.a(new_n199), .b(\b[16] ), .c(new_n200), .d(\b[17] ), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  oaoi03aa1n12x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n190), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n202), .c(new_n198), .d(new_n186), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nand42aa1n06x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nor042aa1n04x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nand42aa1n08x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nanb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  aoai13aa1n03x5               g117(.a(new_n212), .b(new_n208), .c(new_n205), .d(new_n209), .o1(new_n213));
  nanp02aa1n03x5               g118(.a(new_n187), .b(new_n201), .o1(new_n214));
  nanb02aa1n02x5               g119(.a(new_n208), .b(new_n209), .out0(new_n215));
  norb03aa1n02x5               g120(.a(new_n211), .b(new_n208), .c(new_n210), .out0(new_n216));
  aoai13aa1n03x5               g121(.a(new_n216), .b(new_n215), .c(new_n214), .d(new_n204), .o1(new_n217));
  nanp02aa1n03x5               g122(.a(new_n213), .b(new_n217), .o1(\s[20] ));
  nano23aa1d15x5               g123(.a(new_n208), .b(new_n210), .c(new_n211), .d(new_n209), .out0(new_n219));
  nanb03aa1n06x5               g124(.a(new_n193), .b(new_n219), .c(new_n191), .out0(new_n220));
  nand02aa1d04x5               g125(.a(new_n219), .b(new_n203), .o1(new_n221));
  oaih12aa1n06x5               g126(.a(new_n211), .b(new_n210), .c(new_n208), .o1(new_n222));
  nanp02aa1n06x5               g127(.a(new_n221), .b(new_n222), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n220), .c(new_n198), .d(new_n186), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  nanp02aa1n24x5               g132(.a(\b[20] ), .b(\a[21] ), .o1(new_n228));
  norb02aa1n02x5               g133(.a(new_n228), .b(new_n227), .out0(new_n229));
  nor042aa1n12x5               g134(.a(\b[21] ), .b(\a[22] ), .o1(new_n230));
  nanp02aa1n12x5               g135(.a(\b[21] ), .b(\a[22] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  aoai13aa1n02x5               g138(.a(new_n233), .b(new_n227), .c(new_n225), .d(new_n229), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(new_n225), .b(new_n229), .o1(new_n235));
  norb03aa1n02x5               g140(.a(new_n231), .b(new_n227), .c(new_n230), .out0(new_n236));
  nand42aa1n02x5               g141(.a(new_n235), .b(new_n236), .o1(new_n237));
  nanp02aa1n03x5               g142(.a(new_n234), .b(new_n237), .o1(\s[22] ));
  nano23aa1d15x5               g143(.a(new_n227), .b(new_n230), .c(new_n231), .d(new_n228), .out0(new_n239));
  nanp03aa1n02x5               g144(.a(new_n201), .b(new_n219), .c(new_n239), .o1(new_n240));
  and002aa1n02x5               g145(.a(\b[21] ), .b(\a[22] ), .o(new_n241));
  oab012aa1n02x4               g146(.a(new_n241), .b(new_n227), .c(new_n230), .out0(new_n242));
  tech160nm_fiaoi012aa1n05x5   g147(.a(new_n242), .b(new_n223), .c(new_n239), .o1(new_n243));
  aoai13aa1n04x5               g148(.a(new_n243), .b(new_n240), .c(new_n198), .d(new_n186), .o1(new_n244));
  xorb03aa1n02x5               g149(.a(new_n244), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n02x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  nand42aa1n10x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  norb02aa1n02x5               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  nor002aa1d32x5               g153(.a(\b[23] ), .b(\a[24] ), .o1(new_n249));
  nand42aa1d28x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  nanb02aa1n02x5               g155(.a(new_n249), .b(new_n250), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n246), .c(new_n244), .d(new_n248), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n219), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n239), .o1(new_n254));
  nona32aa1n03x5               g159(.a(new_n187), .b(new_n254), .c(new_n253), .d(new_n202), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n248), .o1(new_n256));
  inv040aa1n09x5               g161(.a(new_n249), .o1(new_n257));
  oai112aa1n06x5               g162(.a(new_n257), .b(new_n250), .c(\b[22] ), .d(\a[23] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  aoai13aa1n03x5               g164(.a(new_n259), .b(new_n256), .c(new_n255), .d(new_n243), .o1(new_n260));
  nanp02aa1n03x5               g165(.a(new_n252), .b(new_n260), .o1(\s[24] ));
  nano23aa1n03x7               g166(.a(new_n246), .b(new_n249), .c(new_n250), .d(new_n247), .out0(new_n262));
  nona23aa1n02x4               g167(.a(new_n201), .b(new_n262), .c(new_n254), .d(new_n253), .out0(new_n263));
  nand02aa1n02x5               g168(.a(new_n262), .b(new_n239), .o1(new_n264));
  aoi022aa1n06x5               g169(.a(new_n262), .b(new_n242), .c(new_n250), .d(new_n258), .o1(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n264), .c(new_n221), .d(new_n222), .o1(new_n266));
  inv030aa1n02x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n263), .c(new_n198), .d(new_n186), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  xnrc02aa1n12x5               g175(.a(\b[24] ), .b(\a[25] ), .out0(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  xnrc02aa1n02x5               g177(.a(\b[25] ), .b(\a[26] ), .out0(new_n273));
  aoai13aa1n02x7               g178(.a(new_n273), .b(new_n270), .c(new_n268), .d(new_n272), .o1(new_n274));
  nona32aa1n03x5               g179(.a(new_n187), .b(new_n264), .c(new_n253), .d(new_n202), .out0(new_n275));
  oabi12aa1n12x5               g180(.a(new_n273), .b(\a[25] ), .c(\b[24] ), .out0(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n277), .b(new_n271), .c(new_n275), .d(new_n267), .o1(new_n278));
  nanp02aa1n03x5               g183(.a(new_n274), .b(new_n278), .o1(\s[26] ));
  nor022aa1n04x5               g184(.a(new_n273), .b(new_n271), .o1(new_n280));
  nano32aa1n06x5               g185(.a(new_n220), .b(new_n280), .c(new_n239), .d(new_n262), .out0(new_n281));
  inv020aa1n03x5               g186(.a(new_n281), .o1(new_n282));
  nanp02aa1n02x5               g187(.a(\b[25] ), .b(\a[26] ), .o1(new_n283));
  aoi022aa1n06x5               g188(.a(new_n266), .b(new_n280), .c(new_n283), .d(new_n276), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n282), .c(new_n198), .d(new_n186), .o1(new_n285));
  xorb03aa1n03x5               g190(.a(new_n285), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor002aa1n02x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  xorc02aa1n02x5               g192(.a(\a[27] ), .b(\b[26] ), .out0(new_n288));
  xnrc02aa1n02x5               g193(.a(\b[27] ), .b(\a[28] ), .out0(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n287), .c(new_n285), .d(new_n288), .o1(new_n290));
  tech160nm_finand02aa1n03p5x5 g195(.a(new_n266), .b(new_n280), .o1(new_n291));
  oaib12aa1n06x5               g196(.a(new_n291), .b(new_n277), .c(new_n283), .out0(new_n292));
  aoai13aa1n03x5               g197(.a(new_n288), .b(new_n292), .c(new_n187), .d(new_n281), .o1(new_n293));
  nona22aa1n02x4               g198(.a(new_n293), .b(new_n289), .c(new_n287), .out0(new_n294));
  nanp02aa1n03x5               g199(.a(new_n290), .b(new_n294), .o1(\s[28] ));
  norb02aa1n02x5               g200(.a(new_n288), .b(new_n289), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n296), .b(new_n292), .c(new_n187), .d(new_n281), .o1(new_n297));
  tech160nm_fixorc02aa1n03p5x5 g202(.a(\a[29] ), .b(\b[28] ), .out0(new_n298));
  inv000aa1d42x5               g203(.a(new_n298), .o1(new_n299));
  inv000aa1d42x5               g204(.a(\a[28] ), .o1(new_n300));
  inv000aa1d42x5               g205(.a(\b[27] ), .o1(new_n301));
  oao003aa1n02x5               g206(.a(new_n300), .b(new_n301), .c(new_n287), .carry(new_n302));
  nona22aa1n03x5               g207(.a(new_n297), .b(new_n299), .c(new_n302), .out0(new_n303));
  aoai13aa1n03x5               g208(.a(new_n299), .b(new_n302), .c(new_n285), .d(new_n296), .o1(new_n304));
  nanp02aa1n03x5               g209(.a(new_n304), .b(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g211(.a(new_n289), .b(new_n288), .c(new_n298), .out0(new_n307));
  inv000aa1n03x5               g212(.a(new_n302), .o1(new_n308));
  oaoi03aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .o1(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[29] ), .b(\a[30] ), .out0(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n309), .c(new_n285), .d(new_n307), .o1(new_n311));
  aoai13aa1n02x5               g216(.a(new_n307), .b(new_n292), .c(new_n187), .d(new_n281), .o1(new_n312));
  nona22aa1n02x4               g217(.a(new_n312), .b(new_n309), .c(new_n310), .out0(new_n313));
  nanp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[30] ));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  nano23aa1n02x4               g220(.a(new_n310), .b(new_n289), .c(new_n288), .d(new_n298), .out0(new_n316));
  and002aa1n02x5               g221(.a(\b[29] ), .b(\a[30] ), .o(new_n317));
  oab012aa1n02x4               g222(.a(new_n317), .b(new_n309), .c(new_n310), .out0(new_n318));
  aoai13aa1n03x5               g223(.a(new_n315), .b(new_n318), .c(new_n285), .d(new_n316), .o1(new_n319));
  aoai13aa1n03x5               g224(.a(new_n316), .b(new_n292), .c(new_n187), .d(new_n281), .o1(new_n320));
  nona22aa1n03x5               g225(.a(new_n320), .b(new_n318), .c(new_n315), .out0(new_n321));
  nanp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[31] ));
  xnrb03aa1n02x5               g227(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  norp02aa1n02x5               g228(.a(new_n107), .b(new_n108), .o1(new_n324));
  oab012aa1n02x4               g229(.a(new_n109), .b(new_n116), .c(new_n112), .out0(new_n325));
  oai012aa1n02x5               g230(.a(new_n133), .b(new_n325), .c(new_n324), .o1(\s[4] ));
  xorb03aa1n02x5               g231(.a(new_n117), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb03aa1n03x5               g232(.a(new_n107), .b(new_n133), .c(new_n104), .out0(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n105), .b(new_n328), .c(new_n130), .out0(\s[6] ));
  nona32aa1n02x4               g234(.a(new_n328), .b(new_n120), .c(new_n119), .d(new_n118), .out0(new_n330));
  nona23aa1n03x5               g235(.a(new_n330), .b(new_n102), .c(new_n101), .d(new_n120), .out0(new_n331));
  inv000aa1d42x5               g236(.a(new_n101), .o1(new_n332));
  aboi22aa1n03x5               g237(.a(new_n120), .b(new_n330), .c(new_n332), .d(new_n102), .out0(new_n333));
  norb02aa1n02x5               g238(.a(new_n331), .b(new_n333), .out0(\s[7] ));
  norb02aa1n02x5               g239(.a(new_n100), .b(new_n99), .out0(new_n335));
  xnbna2aa1n03x5               g240(.a(new_n335), .b(new_n331), .c(new_n332), .out0(\s[8] ));
  xnbna2aa1n03x5               g241(.a(new_n124), .b(new_n134), .c(new_n136), .out0(\s[9] ));
endmodule


