// Benchmark "adder" written by ABC on Wed Jul 17 22:30:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n133,
    new_n135, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n180, new_n181,
    new_n182, new_n183, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n330,
    new_n332, new_n335, new_n337, new_n339;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nand22aa1n12x5               g001(.a(\b[0] ), .b(\a[1] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nor042aa1n06x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  oai112aa1n06x5               g005(.a(new_n100), .b(new_n98), .c(new_n99), .d(new_n97), .o1(new_n101));
  oa0022aa1n06x5               g006(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n102));
  aoi022aa1n12x5               g007(.a(new_n101), .b(new_n102), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  inv040aa1d32x5               g008(.a(\a[5] ), .o1(new_n104));
  inv040aa1d32x5               g009(.a(\b[4] ), .o1(new_n105));
  tech160nm_finand02aa1n03p5x5 g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nor042aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  nand02aa1d08x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  norb02aa1n06x5               g014(.a(new_n109), .b(new_n108), .out0(new_n110));
  norp02aa1n04x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nand22aa1n12x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nor022aa1n06x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nona23aa1n03x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  nano32aa1n03x7               g020(.a(new_n115), .b(new_n110), .c(new_n107), .d(new_n106), .out0(new_n116));
  nano22aa1n03x5               g021(.a(new_n113), .b(new_n112), .c(new_n114), .out0(new_n117));
  oaoi03aa1n03x5               g022(.a(\a[6] ), .b(\b[5] ), .c(new_n106), .o1(new_n118));
  ao0012aa1n03x7               g023(.a(new_n111), .b(new_n113), .c(new_n112), .o(new_n119));
  ao0012aa1n12x5               g024(.a(new_n119), .b(new_n118), .c(new_n117), .o(new_n120));
  xorc02aa1n12x5               g025(.a(\a[9] ), .b(\b[8] ), .out0(new_n121));
  aoai13aa1n02x5               g026(.a(new_n121), .b(new_n120), .c(new_n103), .d(new_n116), .o1(new_n122));
  oai012aa1n02x5               g027(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .o1(new_n123));
  xorb03aa1n02x5               g028(.a(new_n123), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand02aa1d16x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  nor002aa1d32x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nand02aa1d08x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n126), .b(new_n127), .out0(new_n128));
  nor002aa1d32x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nor002aa1n16x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nona22aa1n02x4               g035(.a(new_n122), .b(new_n130), .c(new_n129), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n128), .b(new_n131), .c(new_n125), .out0(\s[11] ));
  aoi013aa1n03x5               g037(.a(new_n126), .b(new_n131), .c(new_n127), .d(new_n125), .o1(new_n133));
  xnrb03aa1n02x5               g038(.a(new_n133), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norb03aa1n12x5               g039(.a(new_n125), .b(new_n129), .c(new_n126), .out0(new_n135));
  nor042aa1n12x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nand02aa1n16x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  nano22aa1n12x5               g042(.a(new_n136), .b(new_n127), .c(new_n137), .out0(new_n138));
  nand23aa1d12x5               g043(.a(new_n138), .b(new_n121), .c(new_n135), .o1(new_n139));
  inv040aa1n03x5               g044(.a(new_n139), .o1(new_n140));
  aoai13aa1n06x5               g045(.a(new_n140), .b(new_n120), .c(new_n103), .d(new_n116), .o1(new_n141));
  nanb03aa1d24x5               g046(.a(new_n136), .b(new_n137), .c(new_n127), .out0(new_n142));
  inv020aa1n04x5               g047(.a(new_n126), .o1(new_n143));
  oai112aa1n06x5               g048(.a(new_n143), .b(new_n125), .c(new_n130), .d(new_n129), .o1(new_n144));
  aoi012aa1d18x5               g049(.a(new_n136), .b(new_n126), .c(new_n137), .o1(new_n145));
  oai012aa1d24x5               g050(.a(new_n145), .b(new_n144), .c(new_n142), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  tech160nm_fixorc02aa1n04x5   g052(.a(\a[13] ), .b(\b[12] ), .out0(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n141), .c(new_n147), .out0(\s[13] ));
  inv000aa1d42x5               g054(.a(\a[13] ), .o1(new_n150));
  inv000aa1d42x5               g055(.a(\b[12] ), .o1(new_n151));
  nand02aa1d12x5               g056(.a(new_n151), .b(new_n150), .o1(new_n152));
  aob012aa1n02x5               g057(.a(new_n148), .b(new_n141), .c(new_n147), .out0(new_n153));
  nor042aa1n02x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nand22aa1n02x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  norb02aa1n03x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n153), .c(new_n152), .out0(\s[14] ));
  nand42aa1n02x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand23aa1n03x5               g063(.a(new_n156), .b(new_n152), .c(new_n158), .o1(new_n159));
  oaoi03aa1n12x5               g064(.a(\a[14] ), .b(\b[13] ), .c(new_n152), .o1(new_n160));
  inv030aa1n02x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n04x5               g066(.a(new_n161), .b(new_n159), .c(new_n141), .d(new_n147), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand22aa1n09x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nor002aa1n03x5               g070(.a(\b[15] ), .b(\a[16] ), .o1(new_n166));
  nand22aa1n09x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoi112aa1n02x5               g073(.a(new_n164), .b(new_n168), .c(new_n162), .d(new_n165), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n168), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(\s[16] ));
  nano23aa1n06x5               g076(.a(new_n164), .b(new_n166), .c(new_n167), .d(new_n165), .out0(new_n172));
  nano32aa1n03x7               g077(.a(new_n139), .b(new_n172), .c(new_n148), .d(new_n156), .out0(new_n173));
  aoai13aa1n06x5               g078(.a(new_n173), .b(new_n120), .c(new_n103), .d(new_n116), .o1(new_n174));
  nano32aa1n03x7               g079(.a(new_n154), .b(new_n152), .c(new_n155), .d(new_n158), .out0(new_n175));
  aoai13aa1n12x5               g080(.a(new_n172), .b(new_n160), .c(new_n146), .d(new_n175), .o1(new_n176));
  tech160nm_fiaoi012aa1n03p5x5 g081(.a(new_n166), .b(new_n164), .c(new_n167), .o1(new_n177));
  nanp03aa1d12x5               g082(.a(new_n174), .b(new_n176), .c(new_n177), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g084(.a(\a[18] ), .o1(new_n180));
  inv000aa1d42x5               g085(.a(\a[17] ), .o1(new_n181));
  inv040aa1d32x5               g086(.a(\b[16] ), .o1(new_n182));
  tech160nm_fioaoi03aa1n03p5x5 g087(.a(new_n181), .b(new_n182), .c(new_n178), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[17] ), .c(new_n180), .out0(\s[18] ));
  and002aa1n02x5               g089(.a(\b[17] ), .b(\a[18] ), .o(new_n185));
  nand42aa1n02x5               g090(.a(new_n116), .b(new_n103), .o1(new_n186));
  aoi012aa1n02x5               g091(.a(new_n119), .b(new_n118), .c(new_n117), .o1(new_n187));
  inv020aa1n03x5               g092(.a(new_n172), .o1(new_n188));
  nona22aa1n03x5               g093(.a(new_n140), .b(new_n159), .c(new_n188), .out0(new_n189));
  aoi012aa1n06x5               g094(.a(new_n189), .b(new_n186), .c(new_n187), .o1(new_n190));
  oai012aa1n02x5               g095(.a(new_n125), .b(\b[10] ), .c(\a[11] ), .o1(new_n191));
  oab012aa1n02x4               g096(.a(new_n191), .b(new_n129), .c(new_n130), .out0(new_n192));
  inv020aa1n03x5               g097(.a(new_n145), .o1(new_n193));
  aoai13aa1n04x5               g098(.a(new_n175), .b(new_n193), .c(new_n192), .d(new_n138), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n177), .b(new_n188), .c(new_n194), .d(new_n161), .o1(new_n195));
  xroi22aa1d06x4               g100(.a(new_n181), .b(\b[16] ), .c(new_n180), .d(\b[17] ), .out0(new_n196));
  tech160nm_fioai012aa1n05x5   g101(.a(new_n196), .b(new_n190), .c(new_n195), .o1(new_n197));
  aboi22aa1n02x7               g102(.a(\b[17] ), .b(new_n180), .c(new_n181), .d(new_n182), .out0(new_n198));
  inv000aa1d42x5               g103(.a(\a[19] ), .o1(new_n199));
  nanb02aa1d24x5               g104(.a(\b[18] ), .b(new_n199), .out0(new_n200));
  nand42aa1d28x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  tech160nm_finand02aa1n05x5   g106(.a(new_n200), .b(new_n201), .o1(new_n202));
  oaoi13aa1n06x5               g107(.a(new_n202), .b(new_n197), .c(new_n185), .d(new_n198), .o1(new_n203));
  oaih22aa1n06x5               g108(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n204), .b(new_n185), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n202), .o1(new_n206));
  aoi112aa1n02x5               g111(.a(new_n206), .b(new_n205), .c(new_n178), .d(new_n196), .o1(new_n207));
  norp02aa1n02x5               g112(.a(new_n203), .b(new_n207), .o1(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g114(.a(\a[20] ), .o1(new_n210));
  inv000aa1d42x5               g115(.a(\b[19] ), .o1(new_n211));
  nand22aa1n09x5               g116(.a(new_n211), .b(new_n210), .o1(new_n212));
  nand22aa1n04x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nanp02aa1n02x5               g118(.a(new_n212), .b(new_n213), .o1(new_n214));
  nano22aa1n02x4               g119(.a(new_n203), .b(new_n200), .c(new_n214), .out0(new_n215));
  aoai13aa1n03x5               g120(.a(new_n206), .b(new_n205), .c(new_n178), .d(new_n196), .o1(new_n216));
  aoi012aa1n03x5               g121(.a(new_n214), .b(new_n216), .c(new_n200), .o1(new_n217));
  nor002aa1n02x5               g122(.a(new_n217), .b(new_n215), .o1(\s[20] ));
  nor002aa1n06x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n201), .o1(new_n220));
  nona32aa1d18x5               g125(.a(new_n196), .b(new_n214), .c(new_n220), .d(new_n219), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  tech160nm_fioai012aa1n05x5   g127(.a(new_n222), .b(new_n190), .c(new_n195), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[17] ), .o1(new_n224));
  oai112aa1n06x5               g129(.a(new_n200), .b(new_n201), .c(new_n224), .d(new_n180), .o1(new_n225));
  nand23aa1n04x5               g130(.a(new_n204), .b(new_n212), .c(new_n213), .o1(new_n226));
  oaoi03aa1n12x5               g131(.a(new_n210), .b(new_n211), .c(new_n219), .o1(new_n227));
  oai012aa1d24x5               g132(.a(new_n227), .b(new_n226), .c(new_n225), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  nor042aa1n04x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nanp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n02x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  xnbna2aa1n03x5               g137(.a(new_n232), .b(new_n223), .c(new_n229), .out0(\s[21] ));
  inv000aa1n06x5               g138(.a(new_n230), .o1(new_n234));
  aobi12aa1n06x5               g139(.a(new_n232), .b(new_n223), .c(new_n229), .out0(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[21] ), .b(\a[22] ), .out0(new_n236));
  nano22aa1n03x5               g141(.a(new_n235), .b(new_n234), .c(new_n236), .out0(new_n237));
  aoai13aa1n03x5               g142(.a(new_n232), .b(new_n228), .c(new_n178), .d(new_n222), .o1(new_n238));
  tech160nm_fiaoi012aa1n02p5x5 g143(.a(new_n236), .b(new_n238), .c(new_n234), .o1(new_n239));
  nor002aa1n02x5               g144(.a(new_n239), .b(new_n237), .o1(\s[22] ));
  nano22aa1n03x7               g145(.a(new_n236), .b(new_n234), .c(new_n231), .out0(new_n241));
  nano32aa1n06x5               g146(.a(new_n214), .b(new_n196), .c(new_n241), .d(new_n206), .out0(new_n242));
  oai012aa1n03x5               g147(.a(new_n242), .b(new_n190), .c(new_n195), .o1(new_n243));
  aoi112aa1n02x5               g148(.a(new_n220), .b(new_n219), .c(\a[18] ), .d(\b[17] ), .o1(new_n244));
  nano22aa1n03x5               g149(.a(new_n198), .b(new_n212), .c(new_n213), .out0(new_n245));
  aob012aa1n02x5               g150(.a(new_n212), .b(new_n219), .c(new_n213), .out0(new_n246));
  aoai13aa1n03x5               g151(.a(new_n241), .b(new_n246), .c(new_n245), .d(new_n244), .o1(new_n247));
  oao003aa1n02x5               g152(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .carry(new_n248));
  nanp02aa1n02x5               g153(.a(new_n247), .b(new_n248), .o1(new_n249));
  xnrc02aa1n12x5               g154(.a(\b[22] ), .b(\a[23] ), .out0(new_n250));
  aoib12aa1n06x5               g155(.a(new_n250), .b(new_n243), .c(new_n249), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n250), .o1(new_n252));
  aoi112aa1n02x5               g157(.a(new_n252), .b(new_n249), .c(new_n178), .d(new_n242), .o1(new_n253));
  norp02aa1n02x5               g158(.a(new_n251), .b(new_n253), .o1(\s[23] ));
  nor042aa1n03x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  tech160nm_fixnrc02aa1n04x5   g161(.a(\b[23] ), .b(\a[24] ), .out0(new_n257));
  nano22aa1n03x5               g162(.a(new_n251), .b(new_n256), .c(new_n257), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n252), .b(new_n249), .c(new_n178), .d(new_n242), .o1(new_n259));
  aoi012aa1n03x5               g164(.a(new_n257), .b(new_n259), .c(new_n256), .o1(new_n260));
  norp02aa1n03x5               g165(.a(new_n258), .b(new_n260), .o1(\s[24] ));
  nor042aa1n03x5               g166(.a(new_n257), .b(new_n250), .o1(new_n262));
  nano22aa1n03x7               g167(.a(new_n221), .b(new_n241), .c(new_n262), .out0(new_n263));
  oai012aa1n03x5               g168(.a(new_n263), .b(new_n190), .c(new_n195), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n262), .o1(new_n265));
  oao003aa1n02x5               g170(.a(\a[24] ), .b(\b[23] ), .c(new_n256), .carry(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n265), .c(new_n247), .d(new_n248), .o1(new_n267));
  xnrc02aa1n12x5               g172(.a(\b[24] ), .b(\a[25] ), .out0(new_n268));
  aoib12aa1n06x5               g173(.a(new_n268), .b(new_n264), .c(new_n267), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n268), .o1(new_n270));
  aoi112aa1n02x5               g175(.a(new_n270), .b(new_n267), .c(new_n178), .d(new_n263), .o1(new_n271));
  norp02aa1n02x5               g176(.a(new_n269), .b(new_n271), .o1(\s[25] ));
  nor042aa1n09x5               g177(.a(\b[24] ), .b(\a[25] ), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n273), .o1(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[25] ), .b(\a[26] ), .out0(new_n275));
  nano22aa1n03x5               g180(.a(new_n269), .b(new_n274), .c(new_n275), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n270), .b(new_n267), .c(new_n178), .d(new_n263), .o1(new_n277));
  aoi012aa1n03x5               g182(.a(new_n275), .b(new_n277), .c(new_n274), .o1(new_n278));
  nor002aa1n02x5               g183(.a(new_n276), .b(new_n278), .o1(\s[26] ));
  nor042aa1n06x5               g184(.a(new_n275), .b(new_n268), .o1(new_n280));
  nano32aa1d12x5               g185(.a(new_n221), .b(new_n280), .c(new_n241), .d(new_n262), .out0(new_n281));
  oai012aa1n06x5               g186(.a(new_n281), .b(new_n190), .c(new_n195), .o1(new_n282));
  oao003aa1n06x5               g187(.a(\a[26] ), .b(\b[25] ), .c(new_n274), .carry(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  aoi012aa1n06x5               g189(.a(new_n284), .b(new_n267), .c(new_n280), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n282), .out0(\s[27] ));
  nor042aa1n06x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n286), .o1(new_n290));
  aoi012aa1n02x7               g195(.a(new_n290), .b(new_n285), .c(new_n282), .o1(new_n291));
  xnrc02aa1n02x5               g196(.a(\b[27] ), .b(\a[28] ), .out0(new_n292));
  nano22aa1n03x5               g197(.a(new_n291), .b(new_n289), .c(new_n292), .out0(new_n293));
  inv000aa1n02x5               g198(.a(new_n248), .o1(new_n294));
  aoai13aa1n06x5               g199(.a(new_n262), .b(new_n294), .c(new_n228), .d(new_n241), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n280), .o1(new_n296));
  aoai13aa1n12x5               g201(.a(new_n283), .b(new_n296), .c(new_n295), .d(new_n266), .o1(new_n297));
  aoai13aa1n06x5               g202(.a(new_n286), .b(new_n297), .c(new_n178), .d(new_n281), .o1(new_n298));
  tech160nm_fiaoi012aa1n02p5x5 g203(.a(new_n292), .b(new_n298), .c(new_n289), .o1(new_n299));
  norp02aa1n03x5               g204(.a(new_n299), .b(new_n293), .o1(\s[28] ));
  norb02aa1n02x5               g205(.a(new_n286), .b(new_n292), .out0(new_n301));
  aoai13aa1n02x7               g206(.a(new_n301), .b(new_n297), .c(new_n178), .d(new_n281), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  tech160nm_fiaoi012aa1n02p5x5 g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  inv000aa1n02x5               g210(.a(new_n301), .o1(new_n306));
  aoi012aa1n02x7               g211(.a(new_n306), .b(new_n285), .c(new_n282), .o1(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n304), .out0(new_n308));
  nor002aa1n02x5               g213(.a(new_n305), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n97), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n03x5               g215(.a(new_n286), .b(new_n304), .c(new_n292), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n297), .c(new_n178), .d(new_n281), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[29] ), .b(\a[30] ), .out0(new_n314));
  tech160nm_fiaoi012aa1n02p5x5 g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  aoi012aa1n02x7               g221(.a(new_n316), .b(new_n285), .c(new_n282), .o1(new_n317));
  nano22aa1n02x4               g222(.a(new_n317), .b(new_n313), .c(new_n314), .out0(new_n318));
  norp02aa1n03x5               g223(.a(new_n315), .b(new_n318), .o1(\s[30] ));
  nanb02aa1n02x5               g224(.a(\b[30] ), .b(\a[31] ), .out0(new_n320));
  nanb02aa1n02x5               g225(.a(\a[31] ), .b(\b[30] ), .out0(new_n321));
  norb02aa1n03x4               g226(.a(new_n311), .b(new_n314), .out0(new_n322));
  aoai13aa1n06x5               g227(.a(new_n322), .b(new_n297), .c(new_n178), .d(new_n281), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n324));
  aoi022aa1n02x7               g229(.a(new_n323), .b(new_n324), .c(new_n321), .d(new_n320), .o1(new_n325));
  nanp02aa1n02x5               g230(.a(new_n321), .b(new_n320), .o1(new_n326));
  inv000aa1n02x5               g231(.a(new_n324), .o1(new_n327));
  nona22aa1n02x5               g232(.a(new_n323), .b(new_n327), .c(new_n326), .out0(new_n328));
  norb02aa1n03x4               g233(.a(new_n328), .b(new_n325), .out0(\s[31] ));
  oai012aa1n02x5               g234(.a(new_n98), .b(new_n99), .c(new_n97), .o1(new_n330));
  xnrb03aa1n02x5               g235(.a(new_n330), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g236(.a(\a[3] ), .b(\b[2] ), .c(new_n330), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g238(.a(new_n103), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g239(.a(new_n104), .b(new_n105), .c(new_n103), .o1(new_n335));
  xnrc02aa1n02x5               g240(.a(new_n335), .b(new_n110), .out0(\s[6] ));
  aob012aa1n02x5               g241(.a(new_n109), .b(new_n335), .c(new_n110), .out0(new_n337));
  xnrb03aa1n02x5               g242(.a(new_n337), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g243(.a(\a[7] ), .b(\b[6] ), .c(new_n337), .o1(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g245(.a(new_n121), .b(new_n186), .c(new_n187), .out0(\s[9] ));
endmodule


