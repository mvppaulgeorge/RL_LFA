// Benchmark "adder" written by ABC on Thu Jul 18 06:51:26 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n367, new_n370, new_n371, new_n373, new_n374, new_n375, new_n376,
    new_n378;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  and002aa1n24x5               g002(.a(\b[9] ), .b(\a[10] ), .o(new_n98));
  nor042aa1n03x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  orn002aa1n02x5               g004(.a(\a[9] ), .b(\b[8] ), .o(new_n100));
  inv000aa1d42x5               g005(.a(\a[5] ), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\b[4] ), .o1(new_n102));
  nand02aa1n06x5               g007(.a(\b[5] ), .b(\a[6] ), .o1(new_n103));
  nor002aa1n04x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  aoai13aa1n06x5               g009(.a(new_n103), .b(new_n104), .c(new_n102), .d(new_n101), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand42aa1n02x5               g011(.a(\b[7] ), .b(\a[8] ), .o1(new_n107));
  nanb02aa1n06x5               g012(.a(new_n106), .b(new_n107), .out0(new_n108));
  nand02aa1n06x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nor002aa1d24x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanb02aa1d24x5               g015(.a(new_n110), .b(new_n109), .out0(new_n111));
  oai012aa1n02x5               g016(.a(new_n107), .b(new_n110), .c(new_n106), .o1(new_n112));
  oai013aa1n03x5               g017(.a(new_n112), .b(new_n105), .c(new_n108), .d(new_n111), .o1(new_n113));
  nor042aa1n06x5               g018(.a(\b[1] ), .b(\a[2] ), .o1(new_n114));
  nand22aa1n03x5               g019(.a(\b[0] ), .b(\a[1] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  aoi012aa1n06x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  nanp02aa1n02x5               g022(.a(\b[3] ), .b(\a[4] ), .o1(new_n118));
  nor042aa1n02x5               g023(.a(\b[3] ), .b(\a[4] ), .o1(new_n119));
  nanb02aa1n06x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  inv000aa1d42x5               g025(.a(\a[3] ), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\b[2] ), .o1(new_n122));
  nanp02aa1n12x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(\b[2] ), .b(\a[3] ), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(new_n123), .b(new_n124), .o1(new_n125));
  tech160nm_fioaoi03aa1n03p5x5 g030(.a(\a[4] ), .b(\b[3] ), .c(new_n123), .o1(new_n126));
  inv000aa1n02x5               g031(.a(new_n126), .o1(new_n127));
  oai013aa1n09x5               g032(.a(new_n127), .b(new_n117), .c(new_n120), .d(new_n125), .o1(new_n128));
  nor002aa1n02x5               g033(.a(\b[4] ), .b(\a[5] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[4] ), .b(\a[5] ), .o1(new_n130));
  nona23aa1n02x4               g035(.a(new_n103), .b(new_n130), .c(new_n129), .d(new_n104), .out0(new_n131));
  nor043aa1n03x5               g036(.a(new_n131), .b(new_n111), .c(new_n108), .o1(new_n132));
  norp02aa1n02x5               g037(.a(\b[8] ), .b(\a[9] ), .o1(new_n133));
  nand42aa1n03x5               g038(.a(\b[8] ), .b(\a[9] ), .o1(new_n134));
  norb02aa1n03x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n135), .b(new_n113), .c(new_n128), .d(new_n132), .o1(new_n136));
  xnbna2aa1n03x5               g041(.a(new_n99), .b(new_n136), .c(new_n100), .out0(\s[10] ));
  inv000aa1d42x5               g042(.a(new_n98), .o1(new_n138));
  norp02aa1n04x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1n10x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n15x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  nona22aa1n02x4               g047(.a(new_n136), .b(new_n133), .c(new_n97), .out0(new_n143));
  xnbna2aa1n03x5               g048(.a(new_n142), .b(new_n143), .c(new_n138), .out0(\s[11] ));
  nona22aa1n02x4               g049(.a(new_n143), .b(new_n142), .c(new_n98), .out0(new_n145));
  norp02aa1n04x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nand42aa1n06x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  norb02aa1d21x5               g052(.a(new_n147), .b(new_n146), .out0(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  oaoi13aa1n02x5               g054(.a(new_n149), .b(new_n145), .c(\a[11] ), .d(\b[10] ), .o1(new_n150));
  aoi113aa1n02x5               g055(.a(new_n139), .b(new_n148), .c(new_n143), .d(new_n140), .e(new_n138), .o1(new_n151));
  norp02aa1n02x5               g056(.a(new_n150), .b(new_n151), .o1(\s[12] ));
  inv020aa1n02x5               g057(.a(new_n105), .o1(new_n153));
  nano23aa1n02x5               g058(.a(new_n110), .b(new_n106), .c(new_n107), .d(new_n109), .out0(new_n154));
  aobi12aa1n06x5               g059(.a(new_n112), .b(new_n154), .c(new_n153), .out0(new_n155));
  norp03aa1n02x5               g060(.a(new_n117), .b(new_n120), .c(new_n125), .o1(new_n156));
  oai012aa1n03x5               g061(.a(new_n132), .b(new_n156), .c(new_n126), .o1(new_n157));
  inv040aa1n02x5               g062(.a(new_n99), .o1(new_n158));
  nano32aa1d15x5               g063(.a(new_n158), .b(new_n148), .c(new_n135), .d(new_n141), .out0(new_n159));
  inv000aa1d42x5               g064(.a(new_n159), .o1(new_n160));
  oai022aa1n02x5               g065(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n161));
  oai022aa1n02x5               g066(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n162));
  aoi022aa1n02x5               g067(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n147), .b(new_n161), .c(new_n162), .d(new_n163), .o1(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n160), .c(new_n157), .d(new_n155), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  aoai13aa1n06x5               g071(.a(new_n159), .b(new_n113), .c(new_n128), .d(new_n132), .o1(new_n167));
  nor042aa1n06x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  nand42aa1n06x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  aoai13aa1n02x5               g076(.a(new_n169), .b(new_n171), .c(new_n167), .d(new_n164), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n03x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nand02aa1n06x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nona23aa1d18x5               g080(.a(new_n175), .b(new_n170), .c(new_n168), .d(new_n174), .out0(new_n176));
  oaoi03aa1n02x5               g081(.a(\a[14] ), .b(\b[13] ), .c(new_n169), .o1(new_n177));
  inv000aa1n02x5               g082(.a(new_n177), .o1(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n176), .c(new_n167), .d(new_n164), .o1(new_n179));
  xorb03aa1n02x5               g084(.a(new_n179), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n09x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n176), .o1(new_n183));
  nand42aa1n04x5               g088(.a(\b[14] ), .b(\a[15] ), .o1(new_n184));
  norb02aa1n02x5               g089(.a(new_n184), .b(new_n181), .out0(new_n185));
  aoai13aa1n02x5               g090(.a(new_n185), .b(new_n177), .c(new_n165), .d(new_n183), .o1(new_n186));
  nor002aa1n06x5               g091(.a(\b[15] ), .b(\a[16] ), .o1(new_n187));
  nanp02aa1n04x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  nanb02aa1n02x5               g093(.a(new_n187), .b(new_n188), .out0(new_n189));
  tech160nm_fiaoi012aa1n04x5   g094(.a(new_n189), .b(new_n186), .c(new_n182), .o1(new_n190));
  inv000aa1d42x5               g095(.a(new_n189), .o1(new_n191));
  aoi112aa1n02x5               g096(.a(new_n181), .b(new_n191), .c(new_n179), .d(new_n184), .o1(new_n192));
  norp02aa1n02x5               g097(.a(new_n190), .b(new_n192), .o1(\s[16] ));
  aoi012aa1n02x5               g098(.a(new_n161), .b(new_n162), .c(new_n163), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n175), .b(new_n174), .out0(new_n195));
  norb02aa1n02x7               g100(.a(new_n195), .b(new_n194), .out0(new_n196));
  nanb03aa1n06x5               g101(.a(new_n187), .b(new_n188), .c(new_n184), .out0(new_n197));
  oai122aa1n02x7               g102(.a(new_n147), .b(\a[15] ), .c(\b[14] ), .d(\a[13] ), .e(\b[12] ), .o1(new_n198));
  norp03aa1n06x5               g103(.a(new_n197), .b(new_n198), .c(new_n171), .o1(new_n199));
  oai112aa1n03x5               g104(.a(new_n175), .b(new_n184), .c(new_n174), .d(new_n168), .o1(new_n200));
  norp02aa1n02x5               g105(.a(new_n187), .b(new_n181), .o1(new_n201));
  nand42aa1n02x5               g106(.a(new_n200), .b(new_n201), .o1(new_n202));
  aoi022aa1n09x5               g107(.a(new_n196), .b(new_n199), .c(new_n188), .d(new_n202), .o1(new_n203));
  nanp03aa1n02x5               g108(.a(new_n141), .b(new_n135), .c(new_n148), .o1(new_n204));
  inv000aa1n02x5               g109(.a(new_n197), .o1(new_n205));
  nona32aa1n03x5               g110(.a(new_n195), .b(new_n171), .c(new_n181), .d(new_n168), .out0(new_n206));
  nano23aa1n06x5               g111(.a(new_n204), .b(new_n206), .c(new_n205), .d(new_n99), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n113), .c(new_n128), .d(new_n132), .o1(new_n208));
  xorc02aa1n12x5               g113(.a(\a[17] ), .b(\b[16] ), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n208), .c(new_n203), .out0(\s[17] ));
  nor002aa1d32x5               g115(.a(\b[16] ), .b(\a[17] ), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  inv000aa1d42x5               g117(.a(new_n114), .o1(new_n213));
  aob012aa1n02x5               g118(.a(new_n213), .b(new_n115), .c(new_n116), .out0(new_n214));
  norb02aa1n02x5               g119(.a(new_n118), .b(new_n119), .out0(new_n215));
  norp02aa1n02x5               g120(.a(\b[2] ), .b(\a[3] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n124), .b(new_n216), .out0(new_n217));
  nanp03aa1n02x5               g122(.a(new_n214), .b(new_n215), .c(new_n217), .o1(new_n218));
  nano23aa1n02x4               g123(.a(new_n129), .b(new_n104), .c(new_n130), .d(new_n103), .out0(new_n219));
  nona22aa1n02x4               g124(.a(new_n219), .b(new_n108), .c(new_n111), .out0(new_n220));
  aoai13aa1n04x5               g125(.a(new_n155), .b(new_n220), .c(new_n218), .d(new_n127), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(new_n202), .b(new_n188), .o1(new_n222));
  aob012aa1n02x5               g127(.a(new_n222), .b(new_n196), .c(new_n199), .out0(new_n223));
  aoai13aa1n02x5               g128(.a(new_n209), .b(new_n223), .c(new_n221), .d(new_n207), .o1(new_n224));
  xnrc02aa1n02x5               g129(.a(\b[17] ), .b(\a[18] ), .out0(new_n225));
  xobna2aa1n03x5               g130(.a(new_n225), .b(new_n224), .c(new_n212), .out0(\s[18] ));
  inv000aa1d42x5               g131(.a(\a[17] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\a[18] ), .o1(new_n228));
  xroi22aa1d04x5               g133(.a(new_n227), .b(\b[16] ), .c(new_n228), .d(\b[17] ), .out0(new_n229));
  inv000aa1n02x5               g134(.a(new_n229), .o1(new_n230));
  oaoi03aa1n12x5               g135(.a(\a[18] ), .b(\b[17] ), .c(new_n212), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n231), .o1(new_n232));
  aoai13aa1n04x5               g137(.a(new_n232), .b(new_n230), .c(new_n208), .d(new_n203), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g139(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1d32x5               g140(.a(\b[18] ), .b(\a[19] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  nona32aa1n09x5               g142(.a(new_n159), .b(new_n197), .c(new_n181), .d(new_n176), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n203), .b(new_n238), .c(new_n157), .d(new_n155), .o1(new_n239));
  nand02aa1d06x5               g144(.a(\b[18] ), .b(\a[19] ), .o1(new_n240));
  nanb02aa1d24x5               g145(.a(new_n236), .b(new_n240), .out0(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n231), .c(new_n239), .d(new_n229), .o1(new_n243));
  xnrc02aa1n03x5               g148(.a(\b[19] ), .b(\a[20] ), .out0(new_n244));
  aoi012aa1n03x5               g149(.a(new_n244), .b(new_n243), .c(new_n237), .o1(new_n245));
  inv030aa1n02x5               g150(.a(new_n244), .o1(new_n246));
  aoi112aa1n02x5               g151(.a(new_n236), .b(new_n246), .c(new_n233), .d(new_n240), .o1(new_n247));
  nor002aa1n02x5               g152(.a(new_n245), .b(new_n247), .o1(\s[20] ));
  nona23aa1d18x5               g153(.a(new_n246), .b(new_n209), .c(new_n225), .d(new_n241), .out0(new_n249));
  oab012aa1n06x5               g154(.a(new_n236), .b(\a[20] ), .c(\b[19] ), .out0(new_n250));
  norp02aa1n04x5               g155(.a(\b[17] ), .b(\a[18] ), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[17] ), .b(\a[18] ), .o1(new_n252));
  oai112aa1n06x5               g157(.a(new_n252), .b(new_n240), .c(new_n251), .d(new_n211), .o1(new_n253));
  aoi022aa1d18x5               g158(.a(new_n253), .b(new_n250), .c(\a[20] ), .d(\b[19] ), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  aoai13aa1n02x7               g160(.a(new_n255), .b(new_n249), .c(new_n208), .d(new_n203), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g162(.a(\b[20] ), .b(\a[21] ), .o1(new_n258));
  inv000aa1n06x5               g163(.a(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n249), .o1(new_n260));
  nanp02aa1n04x5               g165(.a(\b[20] ), .b(\a[21] ), .o1(new_n261));
  norb02aa1n02x5               g166(.a(new_n261), .b(new_n258), .out0(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n254), .c(new_n239), .d(new_n260), .o1(new_n263));
  inv000aa1d42x5               g168(.a(\a[22] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(\b[21] ), .o1(new_n265));
  nand22aa1n06x5               g170(.a(new_n265), .b(new_n264), .o1(new_n266));
  nand22aa1n04x5               g171(.a(\b[21] ), .b(\a[22] ), .o1(new_n267));
  nand02aa1d10x5               g172(.a(new_n266), .b(new_n267), .o1(new_n268));
  tech160nm_fiaoi012aa1n02p5x5 g173(.a(new_n268), .b(new_n263), .c(new_n259), .o1(new_n269));
  inv000aa1d42x5               g174(.a(new_n268), .o1(new_n270));
  aoi112aa1n02x5               g175(.a(new_n258), .b(new_n270), .c(new_n256), .d(new_n261), .o1(new_n271));
  nor002aa1n02x5               g176(.a(new_n269), .b(new_n271), .o1(\s[22] ));
  nano22aa1n03x7               g177(.a(new_n268), .b(new_n259), .c(new_n261), .out0(new_n273));
  nano32aa1n02x4               g178(.a(new_n230), .b(new_n273), .c(new_n242), .d(new_n246), .out0(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nand02aa1d04x5               g180(.a(new_n253), .b(new_n250), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(\b[19] ), .b(\a[20] ), .o1(new_n277));
  nano32aa1d12x5               g182(.a(new_n268), .b(new_n259), .c(new_n261), .d(new_n277), .out0(new_n278));
  oaoi03aa1n09x5               g183(.a(\a[22] ), .b(\b[21] ), .c(new_n259), .o1(new_n279));
  aoi012aa1n09x5               g184(.a(new_n279), .b(new_n276), .c(new_n278), .o1(new_n280));
  aoai13aa1n06x5               g185(.a(new_n280), .b(new_n275), .c(new_n208), .d(new_n203), .o1(new_n281));
  xorb03aa1n02x5               g186(.a(new_n281), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g187(.a(\b[22] ), .b(\a[23] ), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n283), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n280), .o1(new_n285));
  xorc02aa1n02x5               g190(.a(\a[23] ), .b(\b[22] ), .out0(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n239), .d(new_n274), .o1(new_n287));
  xorc02aa1n12x5               g192(.a(\a[24] ), .b(\b[23] ), .out0(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  tech160nm_fiaoi012aa1n02p5x5 g194(.a(new_n289), .b(new_n287), .c(new_n284), .o1(new_n290));
  aoi112aa1n02x5               g195(.a(new_n283), .b(new_n288), .c(new_n281), .d(new_n286), .o1(new_n291));
  nor002aa1n02x5               g196(.a(new_n290), .b(new_n291), .o1(\s[24] ));
  inv000aa1n02x5               g197(.a(new_n250), .o1(new_n293));
  norp02aa1n02x5               g198(.a(new_n251), .b(new_n211), .o1(new_n294));
  nano22aa1n03x7               g199(.a(new_n294), .b(new_n252), .c(new_n240), .out0(new_n295));
  oai012aa1n06x5               g200(.a(new_n278), .b(new_n295), .c(new_n293), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n279), .o1(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[22] ), .b(\a[23] ), .out0(new_n298));
  norb02aa1n06x5               g203(.a(new_n288), .b(new_n298), .out0(new_n299));
  inv040aa1n03x5               g204(.a(new_n299), .o1(new_n300));
  nanp02aa1n02x5               g205(.a(\b[23] ), .b(\a[24] ), .o1(new_n301));
  oai022aa1n02x5               g206(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n302));
  nanp02aa1n02x5               g207(.a(new_n302), .b(new_n301), .o1(new_n303));
  aoai13aa1n12x5               g208(.a(new_n303), .b(new_n300), .c(new_n296), .d(new_n297), .o1(new_n304));
  inv000aa1n02x5               g209(.a(new_n304), .o1(new_n305));
  nano32aa1n02x5               g210(.a(new_n249), .b(new_n288), .c(new_n273), .d(new_n286), .out0(new_n306));
  inv000aa1n02x5               g211(.a(new_n306), .o1(new_n307));
  aoai13aa1n02x7               g212(.a(new_n305), .b(new_n307), .c(new_n208), .d(new_n203), .o1(new_n308));
  xorb03aa1n02x5               g213(.a(new_n308), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g214(.a(\b[24] ), .b(\a[25] ), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n310), .o1(new_n311));
  tech160nm_fixorc02aa1n02p5x5 g216(.a(\a[25] ), .b(\b[24] ), .out0(new_n312));
  aoai13aa1n02x5               g217(.a(new_n312), .b(new_n304), .c(new_n239), .d(new_n306), .o1(new_n313));
  xorc02aa1n12x5               g218(.a(\a[26] ), .b(\b[25] ), .out0(new_n314));
  inv000aa1d42x5               g219(.a(new_n314), .o1(new_n315));
  aoi012aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n311), .o1(new_n316));
  aoi112aa1n02x5               g221(.a(new_n310), .b(new_n314), .c(new_n308), .d(new_n312), .o1(new_n317));
  nor002aa1n02x5               g222(.a(new_n316), .b(new_n317), .o1(\s[26] ));
  and002aa1n12x5               g223(.a(new_n314), .b(new_n312), .o(new_n319));
  nano32aa1n03x7               g224(.a(new_n249), .b(new_n319), .c(new_n273), .d(new_n299), .out0(new_n320));
  aoai13aa1n06x5               g225(.a(new_n320), .b(new_n223), .c(new_n221), .d(new_n207), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[26] ), .b(\b[25] ), .c(new_n311), .carry(new_n322));
  aobi12aa1n12x5               g227(.a(new_n322), .b(new_n304), .c(new_n319), .out0(new_n323));
  xorc02aa1n12x5               g228(.a(\a[27] ), .b(\b[26] ), .out0(new_n324));
  xnbna2aa1n06x5               g229(.a(new_n324), .b(new_n323), .c(new_n321), .out0(\s[27] ));
  norp02aa1n02x5               g230(.a(\b[26] ), .b(\a[27] ), .o1(new_n326));
  inv040aa1n03x5               g231(.a(new_n326), .o1(new_n327));
  aoai13aa1n02x5               g232(.a(new_n299), .b(new_n279), .c(new_n276), .d(new_n278), .o1(new_n328));
  inv000aa1d42x5               g233(.a(new_n319), .o1(new_n329));
  aoai13aa1n06x5               g234(.a(new_n322), .b(new_n329), .c(new_n328), .d(new_n303), .o1(new_n330));
  aoai13aa1n02x7               g235(.a(new_n324), .b(new_n330), .c(new_n239), .d(new_n320), .o1(new_n331));
  xnrc02aa1n12x5               g236(.a(\b[27] ), .b(\a[28] ), .out0(new_n332));
  tech160nm_fiaoi012aa1n02p5x5 g237(.a(new_n332), .b(new_n331), .c(new_n327), .o1(new_n333));
  inv000aa1d42x5               g238(.a(new_n324), .o1(new_n334));
  tech160nm_fiaoi012aa1n03p5x5 g239(.a(new_n334), .b(new_n323), .c(new_n321), .o1(new_n335));
  nano22aa1n03x5               g240(.a(new_n335), .b(new_n327), .c(new_n332), .out0(new_n336));
  norp02aa1n03x5               g241(.a(new_n333), .b(new_n336), .o1(\s[28] ));
  norb02aa1n09x5               g242(.a(new_n324), .b(new_n332), .out0(new_n338));
  aoai13aa1n03x5               g243(.a(new_n338), .b(new_n330), .c(new_n239), .d(new_n320), .o1(new_n339));
  oao003aa1n02x5               g244(.a(\a[28] ), .b(\b[27] ), .c(new_n327), .carry(new_n340));
  xnrc02aa1n12x5               g245(.a(\b[28] ), .b(\a[29] ), .out0(new_n341));
  aoi012aa1n03x5               g246(.a(new_n341), .b(new_n339), .c(new_n340), .o1(new_n342));
  inv000aa1d42x5               g247(.a(new_n338), .o1(new_n343));
  tech160nm_fiaoi012aa1n03p5x5 g248(.a(new_n343), .b(new_n323), .c(new_n321), .o1(new_n344));
  nano22aa1n03x5               g249(.a(new_n344), .b(new_n340), .c(new_n341), .out0(new_n345));
  norp02aa1n03x5               g250(.a(new_n342), .b(new_n345), .o1(\s[29] ));
  xorb03aa1n02x5               g251(.a(new_n115), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1d15x5               g252(.a(new_n324), .b(new_n341), .c(new_n332), .out0(new_n348));
  aoai13aa1n02x5               g253(.a(new_n348), .b(new_n330), .c(new_n239), .d(new_n320), .o1(new_n349));
  oao003aa1n02x5               g254(.a(\a[29] ), .b(\b[28] ), .c(new_n340), .carry(new_n350));
  xnrc02aa1n02x5               g255(.a(\b[29] ), .b(\a[30] ), .out0(new_n351));
  tech160nm_fiaoi012aa1n02p5x5 g256(.a(new_n351), .b(new_n349), .c(new_n350), .o1(new_n352));
  inv000aa1d42x5               g257(.a(new_n348), .o1(new_n353));
  tech160nm_fiaoi012aa1n03p5x5 g258(.a(new_n353), .b(new_n323), .c(new_n321), .o1(new_n354));
  nano22aa1n03x5               g259(.a(new_n354), .b(new_n350), .c(new_n351), .out0(new_n355));
  norp02aa1n03x5               g260(.a(new_n352), .b(new_n355), .o1(\s[30] ));
  xnrc02aa1n02x5               g261(.a(\b[30] ), .b(\a[31] ), .out0(new_n357));
  nona32aa1n02x4               g262(.a(new_n324), .b(new_n351), .c(new_n341), .d(new_n332), .out0(new_n358));
  inv000aa1n02x5               g263(.a(new_n358), .o1(new_n359));
  aoai13aa1n02x5               g264(.a(new_n359), .b(new_n330), .c(new_n239), .d(new_n320), .o1(new_n360));
  oao003aa1n02x5               g265(.a(\a[30] ), .b(\b[29] ), .c(new_n350), .carry(new_n361));
  aoi012aa1n03x5               g266(.a(new_n357), .b(new_n360), .c(new_n361), .o1(new_n362));
  tech160nm_fiaoi012aa1n03p5x5 g267(.a(new_n358), .b(new_n323), .c(new_n321), .o1(new_n363));
  nano22aa1n03x5               g268(.a(new_n363), .b(new_n357), .c(new_n361), .out0(new_n364));
  norp02aa1n03x5               g269(.a(new_n362), .b(new_n364), .o1(\s[31] ));
  xnbna2aa1n03x5               g270(.a(new_n117), .b(new_n124), .c(new_n123), .out0(\s[3] ));
  aoi112aa1n02x5               g271(.a(new_n216), .b(new_n215), .c(new_n214), .d(new_n217), .o1(new_n367));
  aoib12aa1n02x5               g272(.a(new_n367), .b(new_n128), .c(new_n119), .out0(\s[4] ));
  xorb03aa1n02x5               g273(.a(new_n128), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norb02aa1n02x5               g274(.a(new_n103), .b(new_n104), .out0(new_n370));
  oaoi03aa1n02x5               g275(.a(new_n101), .b(new_n102), .c(new_n128), .o1(new_n371));
  xnrc02aa1n02x5               g276(.a(new_n371), .b(new_n370), .out0(\s[6] ));
  inv000aa1d42x5               g277(.a(new_n111), .o1(new_n373));
  nano22aa1n02x4               g278(.a(new_n129), .b(new_n128), .c(new_n130), .out0(new_n374));
  aoai13aa1n06x5               g279(.a(new_n373), .b(new_n153), .c(new_n374), .d(new_n370), .o1(new_n375));
  aoi112aa1n02x5               g280(.a(new_n153), .b(new_n373), .c(new_n374), .d(new_n370), .o1(new_n376));
  norb02aa1n02x5               g281(.a(new_n375), .b(new_n376), .out0(\s[7] ));
  inv000aa1d42x5               g282(.a(new_n110), .o1(new_n378));
  xobna2aa1n03x5               g283(.a(new_n108), .b(new_n375), .c(new_n378), .out0(\s[8] ));
  xorb03aa1n02x5               g284(.a(new_n221), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


