// Benchmark "adder" written by ABC on Thu Jul 18 08:54:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n332, new_n334, new_n335, new_n338, new_n339, new_n341,
    new_n343, new_n344, new_n345;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  orn002aa1n24x5               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nand42aa1n20x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand02aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aob012aa1n12x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .out0(new_n102));
  nor042aa1n03x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norb02aa1n06x4               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  xorc02aa1n12x5               g010(.a(\a[3] ), .b(\b[2] ), .out0(new_n106));
  nanp03aa1d12x5               g011(.a(new_n102), .b(new_n106), .c(new_n105), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[3] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[2] ), .o1(new_n109));
  aoai13aa1n04x5               g014(.a(new_n104), .b(new_n103), .c(new_n108), .d(new_n109), .o1(new_n110));
  nanp02aa1n04x5               g015(.a(new_n107), .b(new_n110), .o1(new_n111));
  xnrc02aa1n12x5               g016(.a(\b[7] ), .b(\a[8] ), .out0(new_n112));
  xorc02aa1n12x5               g017(.a(\a[7] ), .b(\b[6] ), .out0(new_n113));
  xorc02aa1n12x5               g018(.a(\a[6] ), .b(\b[5] ), .out0(new_n114));
  xorc02aa1n12x5               g019(.a(\a[5] ), .b(\b[4] ), .out0(new_n115));
  nano32aa1n03x7               g020(.a(new_n112), .b(new_n115), .c(new_n113), .d(new_n114), .out0(new_n116));
  nor042aa1d18x5               g021(.a(\b[4] ), .b(\a[5] ), .o1(new_n117));
  inv040aa1n02x5               g022(.a(new_n117), .o1(new_n118));
  oaoi03aa1n09x5               g023(.a(\a[6] ), .b(\b[5] ), .c(new_n118), .o1(new_n119));
  nanb03aa1n02x5               g024(.a(new_n112), .b(new_n119), .c(new_n113), .out0(new_n120));
  nanp02aa1n02x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  oai022aa1n02x5               g026(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n122));
  and002aa1n02x5               g027(.a(new_n122), .b(new_n121), .o(new_n123));
  nanb02aa1n02x5               g028(.a(new_n123), .b(new_n120), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n116), .d(new_n111), .o1(new_n126));
  xorc02aa1n12x5               g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n127), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  inv030aa1d32x5               g033(.a(\a[10] ), .o1(new_n129));
  inv030aa1d32x5               g034(.a(\b[9] ), .o1(new_n130));
  aboi22aa1d24x5               g035(.a(\b[8] ), .b(new_n97), .c(new_n130), .d(new_n129), .out0(new_n131));
  nand02aa1n08x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  inv040aa1d32x5               g037(.a(\a[11] ), .o1(new_n133));
  inv040aa1n16x5               g038(.a(\b[10] ), .o1(new_n134));
  nand02aa1d28x5               g039(.a(new_n134), .b(new_n133), .o1(new_n135));
  oai112aa1n02x5               g040(.a(new_n135), .b(new_n132), .c(new_n130), .d(new_n129), .o1(new_n136));
  tech160nm_fiaoi012aa1n02p5x5 g041(.a(new_n136), .b(new_n126), .c(new_n131), .o1(new_n137));
  nanp02aa1n03x5               g042(.a(new_n135), .b(new_n132), .o1(new_n138));
  aoi022aa1n02x5               g043(.a(new_n126), .b(new_n131), .c(\b[9] ), .d(\a[10] ), .o1(new_n139));
  aoib12aa1n02x5               g044(.a(new_n137), .b(new_n138), .c(new_n139), .out0(\s[11] ));
  aoai13aa1n02x5               g045(.a(new_n135), .b(new_n136), .c(new_n126), .d(new_n131), .o1(new_n141));
  xorc02aa1n02x5               g046(.a(\a[12] ), .b(\b[11] ), .out0(new_n142));
  inv000aa1d42x5               g047(.a(\b[11] ), .o1(new_n143));
  nanb02aa1d24x5               g048(.a(\a[12] ), .b(new_n143), .out0(new_n144));
  nand42aa1n16x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  aoi022aa1n02x5               g050(.a(new_n144), .b(new_n145), .c(new_n134), .d(new_n133), .o1(new_n146));
  aboi22aa1n03x5               g051(.a(new_n137), .b(new_n146), .c(new_n141), .d(new_n142), .out0(\s[12] ));
  nano22aa1n03x7               g052(.a(new_n138), .b(new_n144), .c(new_n145), .out0(new_n148));
  nand23aa1d12x5               g053(.a(new_n148), .b(new_n125), .c(new_n127), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n03x5               g055(.a(new_n150), .b(new_n124), .c(new_n116), .d(new_n111), .o1(new_n151));
  oai022aa1d24x5               g056(.a(new_n129), .b(new_n130), .c(\b[10] ), .d(\a[11] ), .o1(new_n152));
  nanp03aa1d12x5               g057(.a(new_n144), .b(new_n132), .c(new_n145), .o1(new_n153));
  aob012aa1d18x5               g058(.a(new_n145), .b(new_n144), .c(new_n135), .out0(new_n154));
  oai013aa1d12x5               g059(.a(new_n154), .b(new_n153), .c(new_n131), .d(new_n152), .o1(new_n155));
  inv000aa1d42x5               g060(.a(new_n155), .o1(new_n156));
  xorc02aa1n02x5               g061(.a(\a[13] ), .b(\b[12] ), .out0(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n151), .c(new_n156), .out0(\s[13] ));
  inv030aa1d32x5               g063(.a(\a[13] ), .o1(new_n159));
  nanb02aa1n12x5               g064(.a(\b[12] ), .b(new_n159), .out0(new_n160));
  xnrc02aa1n02x5               g065(.a(\b[6] ), .b(\a[7] ), .out0(new_n161));
  nona23aa1n09x5               g066(.a(new_n114), .b(new_n115), .c(new_n161), .d(new_n112), .out0(new_n162));
  inv000aa1n02x5               g067(.a(new_n112), .o1(new_n163));
  aoi013aa1n06x4               g068(.a(new_n123), .b(new_n163), .c(new_n119), .d(new_n113), .o1(new_n164));
  aoai13aa1n12x5               g069(.a(new_n164), .b(new_n162), .c(new_n107), .d(new_n110), .o1(new_n165));
  aoai13aa1n03x5               g070(.a(new_n157), .b(new_n155), .c(new_n165), .d(new_n150), .o1(new_n166));
  xorc02aa1n02x5               g071(.a(\a[14] ), .b(\b[13] ), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n166), .c(new_n160), .out0(\s[14] ));
  inv020aa1n04x5               g073(.a(\a[14] ), .o1(new_n169));
  xroi22aa1d06x4               g074(.a(new_n159), .b(\b[12] ), .c(new_n169), .d(\b[13] ), .out0(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n155), .c(new_n165), .d(new_n150), .o1(new_n171));
  oaoi03aa1n09x5               g076(.a(\a[14] ), .b(\b[13] ), .c(new_n160), .o1(new_n172));
  inv000aa1n02x5               g077(.a(new_n172), .o1(new_n173));
  xorc02aa1n12x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n171), .c(new_n173), .out0(\s[15] ));
  nand42aa1n02x5               g080(.a(new_n151), .b(new_n156), .o1(new_n176));
  aoai13aa1n03x5               g081(.a(new_n174), .b(new_n172), .c(new_n176), .d(new_n170), .o1(new_n177));
  nor042aa1d18x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  inv040aa1d28x5               g083(.a(new_n178), .o1(new_n179));
  inv000aa1n02x5               g084(.a(new_n174), .o1(new_n180));
  aoai13aa1n03x5               g085(.a(new_n179), .b(new_n180), .c(new_n171), .d(new_n173), .o1(new_n181));
  xorc02aa1n02x5               g086(.a(\a[16] ), .b(\b[15] ), .out0(new_n182));
  norp02aa1n02x5               g087(.a(new_n182), .b(new_n178), .o1(new_n183));
  aoi022aa1n03x5               g088(.a(new_n181), .b(new_n182), .c(new_n177), .d(new_n183), .o1(\s[16] ));
  nanp02aa1n02x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  xnrc02aa1n12x5               g090(.a(\b[15] ), .b(\a[16] ), .out0(new_n186));
  nano22aa1n09x5               g091(.a(new_n186), .b(new_n179), .c(new_n185), .out0(new_n187));
  nano22aa1d15x5               g092(.a(new_n149), .b(new_n170), .c(new_n187), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n124), .c(new_n116), .d(new_n111), .o1(new_n189));
  oao003aa1n02x5               g094(.a(\a[16] ), .b(\b[15] ), .c(new_n179), .carry(new_n190));
  oai013aa1n03x4               g095(.a(new_n190), .b(new_n173), .c(new_n180), .d(new_n186), .o1(new_n191));
  aoi013aa1n06x4               g096(.a(new_n191), .b(new_n155), .c(new_n170), .d(new_n187), .o1(new_n192));
  xorc02aa1n12x5               g097(.a(\a[17] ), .b(\b[16] ), .out0(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n193), .b(new_n189), .c(new_n192), .out0(\s[17] ));
  inv040aa1d32x5               g099(.a(\a[17] ), .o1(new_n195));
  inv040aa1d28x5               g100(.a(\b[16] ), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n196), .b(new_n195), .o1(new_n197));
  nand03aa1n02x5               g102(.a(new_n155), .b(new_n170), .c(new_n187), .o1(new_n198));
  aobi12aa1n03x7               g103(.a(new_n190), .b(new_n187), .c(new_n172), .out0(new_n199));
  nanp02aa1n06x5               g104(.a(new_n198), .b(new_n199), .o1(new_n200));
  aoai13aa1n04x5               g105(.a(new_n193), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n201));
  nor042aa1n04x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand02aa1d28x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norb02aa1n09x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n201), .c(new_n197), .out0(\s[18] ));
  and002aa1n02x5               g110(.a(new_n193), .b(new_n204), .o(new_n206));
  aoai13aa1n06x5               g111(.a(new_n206), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n207));
  aoi013aa1n09x5               g112(.a(new_n202), .b(new_n203), .c(new_n195), .d(new_n196), .o1(new_n208));
  nor002aa1d32x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand42aa1d28x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  norb02aa1n06x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n207), .c(new_n208), .out0(\s[19] ));
  xnrc02aa1n02x5               g117(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n09x5               g118(.a(new_n189), .b(new_n192), .o1(new_n214));
  oaoi03aa1n02x5               g119(.a(\a[18] ), .b(\b[17] ), .c(new_n197), .o1(new_n215));
  aoai13aa1n03x5               g120(.a(new_n211), .b(new_n215), .c(new_n214), .d(new_n206), .o1(new_n216));
  inv040aa1n08x5               g121(.a(new_n209), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n211), .o1(new_n218));
  aoai13aa1n02x7               g123(.a(new_n217), .b(new_n218), .c(new_n207), .d(new_n208), .o1(new_n219));
  nor002aa1d32x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nand42aa1d28x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  inv000aa1d42x5               g127(.a(\a[19] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[18] ), .o1(new_n224));
  aboi22aa1n03x5               g129(.a(new_n220), .b(new_n221), .c(new_n223), .d(new_n224), .out0(new_n225));
  aoi022aa1n03x5               g130(.a(new_n219), .b(new_n222), .c(new_n216), .d(new_n225), .o1(\s[20] ));
  nano23aa1n06x5               g131(.a(new_n209), .b(new_n220), .c(new_n221), .d(new_n210), .out0(new_n227));
  nand23aa1n06x5               g132(.a(new_n227), .b(new_n193), .c(new_n204), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n230));
  nona23aa1d18x5               g135(.a(new_n221), .b(new_n210), .c(new_n209), .d(new_n220), .out0(new_n231));
  oaoi03aa1n09x5               g136(.a(\a[20] ), .b(\b[19] ), .c(new_n217), .o1(new_n232));
  inv040aa1n02x5               g137(.a(new_n232), .o1(new_n233));
  oai012aa1d24x5               g138(.a(new_n233), .b(new_n231), .c(new_n208), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  xnbna2aa1n03x5               g142(.a(new_n237), .b(new_n230), .c(new_n235), .out0(\s[21] ));
  aoai13aa1n03x5               g143(.a(new_n237), .b(new_n234), .c(new_n214), .d(new_n229), .o1(new_n239));
  nor002aa1d32x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  inv000aa1d42x5               g145(.a(new_n240), .o1(new_n241));
  aoai13aa1n02x7               g146(.a(new_n241), .b(new_n236), .c(new_n230), .d(new_n235), .o1(new_n242));
  xnrc02aa1n12x5               g147(.a(\b[21] ), .b(\a[22] ), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n243), .b(new_n240), .out0(new_n245));
  aoi022aa1n03x5               g150(.a(new_n242), .b(new_n244), .c(new_n239), .d(new_n245), .o1(\s[22] ));
  nor042aa1n06x5               g151(.a(new_n243), .b(new_n236), .o1(new_n247));
  norb02aa1n09x5               g152(.a(new_n247), .b(new_n228), .out0(new_n248));
  aoai13aa1n03x5               g153(.a(new_n248), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n249));
  oao003aa1n12x5               g154(.a(\a[22] ), .b(\b[21] ), .c(new_n241), .carry(new_n250));
  inv000aa1d42x5               g155(.a(new_n250), .o1(new_n251));
  aoi012aa1d18x5               g156(.a(new_n251), .b(new_n234), .c(new_n247), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  xorc02aa1n12x5               g158(.a(\a[23] ), .b(\b[22] ), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n253), .c(new_n214), .d(new_n248), .o1(new_n255));
  aoi112aa1n02x5               g160(.a(new_n254), .b(new_n251), .c(new_n234), .d(new_n247), .o1(new_n256));
  aobi12aa1n02x7               g161(.a(new_n255), .b(new_n256), .c(new_n249), .out0(\s[23] ));
  nor042aa1n09x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n254), .o1(new_n260));
  aoai13aa1n02x7               g165(.a(new_n259), .b(new_n260), .c(new_n249), .d(new_n252), .o1(new_n261));
  tech160nm_fixorc02aa1n03p5x5 g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  norp02aa1n02x5               g167(.a(new_n262), .b(new_n258), .o1(new_n263));
  aoi022aa1n02x7               g168(.a(new_n261), .b(new_n262), .c(new_n255), .d(new_n263), .o1(\s[24] ));
  nano32aa1n03x7               g169(.a(new_n228), .b(new_n262), .c(new_n247), .d(new_n254), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n247), .b(new_n232), .c(new_n227), .d(new_n215), .o1(new_n267));
  and002aa1n06x5               g172(.a(new_n262), .b(new_n254), .o(new_n268));
  inv030aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[24] ), .b(\b[23] ), .c(new_n259), .carry(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n267), .d(new_n250), .o1(new_n271));
  inv000aa1n02x5               g176(.a(new_n271), .o1(new_n272));
  xorc02aa1n12x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  xnbna2aa1n03x5               g178(.a(new_n273), .b(new_n266), .c(new_n272), .out0(\s[25] ));
  aoai13aa1n03x5               g179(.a(new_n273), .b(new_n271), .c(new_n214), .d(new_n265), .o1(new_n275));
  norp02aa1n02x5               g180(.a(\b[24] ), .b(\a[25] ), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n273), .o1(new_n278));
  aoai13aa1n02x7               g183(.a(new_n277), .b(new_n278), .c(new_n266), .d(new_n272), .o1(new_n279));
  xorc02aa1n02x5               g184(.a(\a[26] ), .b(\b[25] ), .out0(new_n280));
  norp02aa1n02x5               g185(.a(new_n280), .b(new_n276), .o1(new_n281));
  aoi022aa1n02x7               g186(.a(new_n279), .b(new_n280), .c(new_n275), .d(new_n281), .o1(\s[26] ));
  and002aa1n03x5               g187(.a(new_n280), .b(new_n273), .o(new_n283));
  inv020aa1n03x5               g188(.a(new_n283), .o1(new_n284));
  nano23aa1n06x5               g189(.a(new_n284), .b(new_n228), .c(new_n268), .d(new_n247), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n200), .c(new_n165), .d(new_n188), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n268), .b(new_n251), .c(new_n234), .d(new_n247), .o1(new_n287));
  nanp02aa1n02x5               g192(.a(\b[25] ), .b(\a[26] ), .o1(new_n288));
  oai022aa1n02x5               g193(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n289));
  nanp02aa1n02x5               g194(.a(new_n289), .b(new_n288), .o1(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n284), .c(new_n287), .d(new_n270), .o1(new_n291));
  xorc02aa1n12x5               g196(.a(\a[27] ), .b(\b[26] ), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n291), .c(new_n214), .d(new_n285), .o1(new_n293));
  aoi122aa1n02x5               g198(.a(new_n292), .b(new_n288), .c(new_n289), .d(new_n271), .e(new_n283), .o1(new_n294));
  aobi12aa1n02x7               g199(.a(new_n293), .b(new_n294), .c(new_n286), .out0(\s[27] ));
  aoi022aa1n02x7               g200(.a(new_n271), .b(new_n283), .c(new_n288), .d(new_n289), .o1(new_n296));
  norp02aa1n02x5               g201(.a(\b[26] ), .b(\a[27] ), .o1(new_n297));
  inv000aa1n03x5               g202(.a(new_n297), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n292), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n298), .b(new_n299), .c(new_n296), .d(new_n286), .o1(new_n300));
  xorc02aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .out0(new_n301));
  norp02aa1n02x5               g206(.a(new_n301), .b(new_n297), .o1(new_n302));
  aoi022aa1n02x7               g207(.a(new_n300), .b(new_n301), .c(new_n293), .d(new_n302), .o1(\s[28] ));
  and002aa1n02x5               g208(.a(new_n301), .b(new_n292), .o(new_n304));
  aoai13aa1n02x5               g209(.a(new_n304), .b(new_n291), .c(new_n214), .d(new_n285), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[28] ), .b(\b[27] ), .c(new_n298), .carry(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n306), .c(new_n296), .d(new_n286), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  norb02aa1n02x5               g214(.a(new_n307), .b(new_n309), .out0(new_n310));
  aoi022aa1n03x5               g215(.a(new_n308), .b(new_n309), .c(new_n305), .d(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g216(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g217(.a(new_n299), .b(new_n301), .c(new_n309), .out0(new_n313));
  aoai13aa1n02x5               g218(.a(new_n313), .b(new_n291), .c(new_n214), .d(new_n285), .o1(new_n314));
  inv000aa1d42x5               g219(.a(new_n313), .o1(new_n315));
  oaoi03aa1n02x5               g220(.a(\a[29] ), .b(\b[28] ), .c(new_n307), .o1(new_n316));
  inv000aa1n03x5               g221(.a(new_n316), .o1(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n315), .c(new_n296), .d(new_n286), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[30] ), .b(\b[29] ), .out0(new_n319));
  and002aa1n02x5               g224(.a(\b[28] ), .b(\a[29] ), .o(new_n320));
  oabi12aa1n02x5               g225(.a(new_n319), .b(\a[29] ), .c(\b[28] ), .out0(new_n321));
  oab012aa1n02x4               g226(.a(new_n321), .b(new_n307), .c(new_n320), .out0(new_n322));
  aoi022aa1n03x5               g227(.a(new_n318), .b(new_n319), .c(new_n314), .d(new_n322), .o1(\s[30] ));
  nano32aa1n03x7               g228(.a(new_n299), .b(new_n319), .c(new_n301), .d(new_n309), .out0(new_n324));
  aoai13aa1n02x5               g229(.a(new_n324), .b(new_n291), .c(new_n214), .d(new_n285), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[31] ), .b(\b[30] ), .out0(new_n326));
  oao003aa1n02x5               g231(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n327));
  norb02aa1n02x5               g232(.a(new_n327), .b(new_n326), .out0(new_n328));
  inv000aa1d42x5               g233(.a(new_n324), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n327), .b(new_n329), .c(new_n296), .d(new_n286), .o1(new_n330));
  aoi022aa1n03x5               g235(.a(new_n330), .b(new_n326), .c(new_n325), .d(new_n328), .o1(\s[31] ));
  nanp03aa1n02x5               g236(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n332));
  xnbna2aa1n03x5               g237(.a(new_n106), .b(new_n332), .c(new_n99), .out0(\s[3] ));
  obai22aa1n02x7               g238(.a(new_n104), .b(new_n103), .c(\a[3] ), .d(\b[2] ), .out0(new_n334));
  aoi012aa1n02x5               g239(.a(new_n334), .b(new_n102), .c(new_n106), .o1(new_n335));
  oaoi13aa1n02x5               g240(.a(new_n335), .b(new_n111), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g241(.a(new_n115), .b(new_n107), .c(new_n110), .out0(\s[5] ));
  aoai13aa1n03x5               g242(.a(new_n114), .b(new_n117), .c(new_n111), .d(new_n115), .o1(new_n338));
  aoi112aa1n02x5               g243(.a(new_n117), .b(new_n114), .c(new_n111), .d(new_n115), .o1(new_n339));
  norb02aa1n02x5               g244(.a(new_n338), .b(new_n339), .out0(\s[6] ));
  orn002aa1n02x5               g245(.a(\a[6] ), .b(\b[5] ), .o(new_n341));
  xnbna2aa1n03x5               g246(.a(new_n113), .b(new_n338), .c(new_n341), .out0(\s[7] ));
  aob012aa1n03x5               g247(.a(new_n113), .b(new_n338), .c(new_n341), .out0(new_n343));
  tech160nm_fioai012aa1n03p5x5 g248(.a(new_n343), .b(\b[6] ), .c(\a[7] ), .o1(new_n344));
  oa0012aa1n02x5               g249(.a(new_n112), .b(\b[6] ), .c(\a[7] ), .o(new_n345));
  aoi022aa1n02x5               g250(.a(new_n344), .b(new_n163), .c(new_n343), .d(new_n345), .o1(\s[8] ));
  xorb03aa1n02x5               g251(.a(new_n165), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


