// Benchmark "adder" written by ABC on Thu Jul 18 10:32:35 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n317, new_n319, new_n321;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor042aa1n06x5               g003(.a(\b[7] ), .b(\a[8] ), .o1(new_n99));
  nand22aa1n04x5               g004(.a(\b[7] ), .b(\a[8] ), .o1(new_n100));
  nor042aa1n12x5               g005(.a(\b[6] ), .b(\a[7] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[6] ), .b(\a[7] ), .o1(new_n102));
  nona23aa1n09x5               g007(.a(new_n102), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n103));
  nand22aa1n03x5               g008(.a(\b[5] ), .b(\a[6] ), .o1(new_n104));
  nor022aa1n06x5               g009(.a(\b[5] ), .b(\a[6] ), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[4] ), .b(\a[5] ), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[4] ), .b(\a[5] ), .o1(new_n107));
  nano23aa1n06x5               g012(.a(new_n106), .b(new_n105), .c(new_n107), .d(new_n104), .out0(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n103), .out0(new_n109));
  nor042aa1n02x5               g014(.a(\b[1] ), .b(\a[2] ), .o1(new_n110));
  nand02aa1d04x5               g015(.a(\b[0] ), .b(\a[1] ), .o1(new_n111));
  nand02aa1d04x5               g016(.a(\b[1] ), .b(\a[2] ), .o1(new_n112));
  aoi012aa1n12x5               g017(.a(new_n110), .b(new_n111), .c(new_n112), .o1(new_n113));
  xnrc02aa1n12x5               g018(.a(\b[3] ), .b(\a[4] ), .out0(new_n114));
  nor002aa1n02x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  tech160nm_finand02aa1n03p5x5 g020(.a(\b[2] ), .b(\a[3] ), .o1(new_n116));
  nanb02aa1n06x5               g021(.a(new_n115), .b(new_n116), .out0(new_n117));
  inv000aa1d42x5               g022(.a(\a[3] ), .o1(new_n118));
  nanb02aa1n03x5               g023(.a(\b[2] ), .b(new_n118), .out0(new_n119));
  oao003aa1n03x5               g024(.a(\a[4] ), .b(\b[3] ), .c(new_n119), .carry(new_n120));
  oai013aa1d12x5               g025(.a(new_n120), .b(new_n114), .c(new_n113), .d(new_n117), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(new_n101), .b(new_n100), .o1(new_n122));
  inv000aa1d42x5               g027(.a(\a[5] ), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\b[4] ), .o1(new_n124));
  aoai13aa1n04x5               g029(.a(new_n104), .b(new_n105), .c(new_n124), .d(new_n123), .o1(new_n125));
  oai122aa1n02x7               g030(.a(new_n122), .b(new_n103), .c(new_n125), .d(\b[7] ), .e(\a[8] ), .o1(new_n126));
  nanp02aa1n04x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n97), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n126), .c(new_n109), .d(new_n121), .o1(new_n129));
  nor022aa1n12x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand02aa1n08x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  nand22aa1n03x5               g038(.a(new_n109), .b(new_n121), .o1(new_n134));
  norp02aa1n03x5               g039(.a(new_n103), .b(new_n125), .o1(new_n135));
  aoi112aa1n03x5               g040(.a(new_n135), .b(new_n99), .c(new_n100), .d(new_n101), .o1(new_n136));
  oai012aa1n12x5               g041(.a(new_n131), .b(new_n130), .c(new_n97), .o1(new_n137));
  nona23aa1d16x5               g042(.a(new_n131), .b(new_n127), .c(new_n97), .d(new_n130), .out0(new_n138));
  aoai13aa1n02x5               g043(.a(new_n137), .b(new_n138), .c(new_n134), .d(new_n136), .o1(new_n139));
  xorb03aa1n02x5               g044(.a(new_n139), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  nand02aa1d08x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  aoi012aa1n02x5               g047(.a(new_n141), .b(new_n139), .c(new_n142), .o1(new_n143));
  xnrb03aa1n02x5               g048(.a(new_n143), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norp02aa1n04x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand02aa1n08x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nona23aa1n12x5               g051(.a(new_n146), .b(new_n142), .c(new_n141), .d(new_n145), .out0(new_n147));
  tech160nm_fiao0012aa1n02p5x5 g052(.a(new_n145), .b(new_n141), .c(new_n146), .o(new_n148));
  oabi12aa1n06x5               g053(.a(new_n148), .b(new_n147), .c(new_n137), .out0(new_n149));
  aoi012aa1n06x5               g054(.a(new_n126), .b(new_n109), .c(new_n121), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n138), .o1(new_n151));
  nano23aa1n06x5               g056(.a(new_n141), .b(new_n145), .c(new_n146), .d(new_n142), .out0(new_n152));
  nano22aa1n03x7               g057(.a(new_n150), .b(new_n151), .c(new_n152), .out0(new_n153));
  tech160nm_fixnrc02aa1n05x5   g058(.a(\b[12] ), .b(\a[13] ), .out0(new_n154));
  oabi12aa1n02x5               g059(.a(new_n154), .b(new_n153), .c(new_n149), .out0(new_n155));
  norb03aa1n02x5               g060(.a(new_n154), .b(new_n153), .c(new_n149), .out0(new_n156));
  norb02aa1n02x5               g061(.a(new_n155), .b(new_n156), .out0(\s[13] ));
  nor042aa1n03x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  inv040aa1n03x5               g063(.a(new_n158), .o1(new_n159));
  xnrc02aa1n12x5               g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  xobna2aa1n03x5               g065(.a(new_n160), .b(new_n155), .c(new_n159), .out0(\s[14] ));
  nor042aa1n06x5               g066(.a(new_n160), .b(new_n154), .o1(new_n162));
  nano32aa1n03x7               g067(.a(new_n150), .b(new_n162), .c(new_n151), .d(new_n152), .out0(new_n163));
  inv040aa1n03x5               g068(.a(new_n137), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n162), .b(new_n148), .c(new_n152), .d(new_n164), .o1(new_n165));
  oao003aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .c(new_n159), .carry(new_n166));
  nano22aa1n03x7               g071(.a(new_n163), .b(new_n165), .c(new_n166), .out0(new_n167));
  xnrb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  oaoi03aa1n03x5               g073(.a(\a[15] ), .b(\b[14] ), .c(new_n167), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  nand03aa1n02x5               g075(.a(new_n152), .b(new_n128), .c(new_n132), .o1(new_n171));
  tech160nm_fixnrc02aa1n04x5   g076(.a(\b[14] ), .b(\a[15] ), .out0(new_n172));
  xnrc02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .out0(new_n173));
  nor042aa1n06x5               g078(.a(new_n173), .b(new_n172), .o1(new_n174));
  nano22aa1n02x5               g079(.a(new_n171), .b(new_n162), .c(new_n174), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n126), .c(new_n109), .d(new_n121), .o1(new_n176));
  inv000aa1n02x5               g081(.a(new_n166), .o1(new_n177));
  aoai13aa1n06x5               g082(.a(new_n174), .b(new_n177), .c(new_n149), .d(new_n162), .o1(new_n178));
  aoi112aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n179));
  oab012aa1n09x5               g084(.a(new_n179), .b(\a[16] ), .c(\b[15] ), .out0(new_n180));
  nand23aa1n06x5               g085(.a(new_n176), .b(new_n178), .c(new_n180), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g087(.a(\a[18] ), .o1(new_n183));
  inv040aa1d32x5               g088(.a(\a[17] ), .o1(new_n184));
  inv030aa1d32x5               g089(.a(\b[16] ), .o1(new_n185));
  oaoi03aa1n02x5               g090(.a(new_n184), .b(new_n185), .c(new_n181), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[17] ), .c(new_n183), .out0(\s[18] ));
  nona23aa1n09x5               g092(.a(new_n174), .b(new_n162), .c(new_n138), .d(new_n147), .out0(new_n188));
  aoi012aa1n12x5               g093(.a(new_n188), .b(new_n134), .c(new_n136), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n174), .o1(new_n190));
  aoai13aa1n12x5               g095(.a(new_n180), .b(new_n190), .c(new_n165), .d(new_n166), .o1(new_n191));
  xroi22aa1d06x4               g096(.a(new_n184), .b(\b[16] ), .c(new_n183), .d(\b[17] ), .out0(new_n192));
  tech160nm_fioai012aa1n05x5   g097(.a(new_n192), .b(new_n189), .c(new_n191), .o1(new_n193));
  oai022aa1n04x5               g098(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n194));
  oaib12aa1n09x5               g099(.a(new_n194), .b(new_n183), .c(\b[17] ), .out0(new_n195));
  nor002aa1d32x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  nand02aa1n16x5               g101(.a(\b[18] ), .b(\a[19] ), .o1(new_n197));
  nanb02aa1n02x5               g102(.a(new_n196), .b(new_n197), .out0(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  xnbna2aa1n03x5               g104(.a(new_n199), .b(new_n193), .c(new_n195), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g106(.a(new_n196), .o1(new_n202));
  tech160nm_fiaoi012aa1n05x5   g107(.a(new_n198), .b(new_n193), .c(new_n195), .o1(new_n203));
  nor042aa1n06x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  nand02aa1d24x5               g109(.a(\b[19] ), .b(\a[20] ), .o1(new_n205));
  nanb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(new_n206));
  nano22aa1n03x7               g111(.a(new_n203), .b(new_n202), .c(new_n206), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(new_n185), .b(new_n184), .o1(new_n208));
  oaoi03aa1n03x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n208), .o1(new_n209));
  aoai13aa1n02x5               g114(.a(new_n199), .b(new_n209), .c(new_n181), .d(new_n192), .o1(new_n210));
  aoi012aa1n03x5               g115(.a(new_n206), .b(new_n210), .c(new_n202), .o1(new_n211));
  norp02aa1n02x5               g116(.a(new_n211), .b(new_n207), .o1(\s[20] ));
  nano23aa1n09x5               g117(.a(new_n196), .b(new_n204), .c(new_n205), .d(new_n197), .out0(new_n213));
  nand22aa1n03x5               g118(.a(new_n192), .b(new_n213), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  tech160nm_fioai012aa1n05x5   g120(.a(new_n215), .b(new_n189), .c(new_n191), .o1(new_n216));
  nona23aa1n09x5               g121(.a(new_n205), .b(new_n197), .c(new_n196), .d(new_n204), .out0(new_n217));
  aoi012aa1n12x5               g122(.a(new_n204), .b(new_n196), .c(new_n205), .o1(new_n218));
  oai012aa1n18x5               g123(.a(new_n218), .b(new_n217), .c(new_n195), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  nor002aa1d32x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  norb02aa1n02x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n216), .c(new_n220), .out0(\s[21] ));
  inv000aa1d42x5               g129(.a(new_n221), .o1(new_n225));
  aobi12aa1n03x5               g130(.a(new_n223), .b(new_n216), .c(new_n220), .out0(new_n226));
  xnrc02aa1n12x5               g131(.a(\b[21] ), .b(\a[22] ), .out0(new_n227));
  nano22aa1n02x4               g132(.a(new_n226), .b(new_n225), .c(new_n227), .out0(new_n228));
  aoai13aa1n02x5               g133(.a(new_n223), .b(new_n219), .c(new_n181), .d(new_n215), .o1(new_n229));
  tech160nm_fiaoi012aa1n02p5x5 g134(.a(new_n227), .b(new_n229), .c(new_n225), .o1(new_n230));
  norp02aa1n02x5               g135(.a(new_n230), .b(new_n228), .o1(\s[22] ));
  nano22aa1n03x7               g136(.a(new_n227), .b(new_n225), .c(new_n222), .out0(new_n232));
  and003aa1n02x5               g137(.a(new_n192), .b(new_n232), .c(new_n213), .o(new_n233));
  tech160nm_fioai012aa1n05x5   g138(.a(new_n233), .b(new_n189), .c(new_n191), .o1(new_n234));
  oao003aa1n12x5               g139(.a(\a[22] ), .b(\b[21] ), .c(new_n225), .carry(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n219), .c(new_n232), .o1(new_n237));
  xnrc02aa1n12x5               g142(.a(\b[22] ), .b(\a[23] ), .out0(new_n238));
  inv000aa1d42x5               g143(.a(new_n238), .o1(new_n239));
  xnbna2aa1n03x5               g144(.a(new_n239), .b(new_n234), .c(new_n237), .out0(\s[23] ));
  nor042aa1n06x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  inv000aa1d42x5               g146(.a(new_n241), .o1(new_n242));
  aoi012aa1n03x5               g147(.a(new_n238), .b(new_n234), .c(new_n237), .o1(new_n243));
  tech160nm_fixnrc02aa1n02p5x5 g148(.a(\b[23] ), .b(\a[24] ), .out0(new_n244));
  nano22aa1n02x4               g149(.a(new_n243), .b(new_n242), .c(new_n244), .out0(new_n245));
  inv000aa1n03x5               g150(.a(new_n237), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n239), .b(new_n246), .c(new_n181), .d(new_n233), .o1(new_n247));
  aoi012aa1n02x5               g152(.a(new_n244), .b(new_n247), .c(new_n242), .o1(new_n248));
  nor002aa1n02x5               g153(.a(new_n248), .b(new_n245), .o1(\s[24] ));
  nor002aa1n04x5               g154(.a(new_n244), .b(new_n238), .o1(new_n250));
  nano22aa1n06x5               g155(.a(new_n214), .b(new_n232), .c(new_n250), .out0(new_n251));
  oai012aa1n06x5               g156(.a(new_n251), .b(new_n189), .c(new_n191), .o1(new_n252));
  inv000aa1n02x5               g157(.a(new_n218), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n232), .b(new_n253), .c(new_n213), .d(new_n209), .o1(new_n254));
  inv000aa1n03x5               g159(.a(new_n250), .o1(new_n255));
  oao003aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n242), .carry(new_n256));
  aoai13aa1n12x5               g161(.a(new_n256), .b(new_n255), .c(new_n254), .d(new_n235), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  xnrc02aa1n12x5               g163(.a(\b[24] ), .b(\a[25] ), .out0(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n252), .c(new_n258), .out0(\s[25] ));
  nor042aa1n03x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  tech160nm_fiaoi012aa1n05x5   g168(.a(new_n259), .b(new_n252), .c(new_n258), .o1(new_n264));
  xnrc02aa1n02x5               g169(.a(\b[25] ), .b(\a[26] ), .out0(new_n265));
  nano22aa1n03x5               g170(.a(new_n264), .b(new_n263), .c(new_n265), .out0(new_n266));
  aoai13aa1n03x5               g171(.a(new_n260), .b(new_n257), .c(new_n181), .d(new_n251), .o1(new_n267));
  aoi012aa1n03x5               g172(.a(new_n265), .b(new_n267), .c(new_n263), .o1(new_n268));
  norp02aa1n03x5               g173(.a(new_n268), .b(new_n266), .o1(\s[26] ));
  nor042aa1n06x5               g174(.a(new_n265), .b(new_n259), .o1(new_n270));
  nano32aa1n03x7               g175(.a(new_n214), .b(new_n270), .c(new_n232), .d(new_n250), .out0(new_n271));
  oai012aa1n12x5               g176(.a(new_n271), .b(new_n189), .c(new_n191), .o1(new_n272));
  oao003aa1n02x5               g177(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n273));
  aobi12aa1n18x5               g178(.a(new_n273), .b(new_n257), .c(new_n270), .out0(new_n274));
  xorc02aa1n12x5               g179(.a(\a[27] ), .b(\b[26] ), .out0(new_n275));
  xnbna2aa1n03x5               g180(.a(new_n275), .b(new_n272), .c(new_n274), .out0(\s[27] ));
  norp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  inv040aa1n03x5               g182(.a(new_n277), .o1(new_n278));
  aobi12aa1n06x5               g183(.a(new_n275), .b(new_n272), .c(new_n274), .out0(new_n279));
  xnrc02aa1n02x5               g184(.a(\b[27] ), .b(\a[28] ), .out0(new_n280));
  nano22aa1n03x7               g185(.a(new_n279), .b(new_n278), .c(new_n280), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n250), .b(new_n236), .c(new_n219), .d(new_n232), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n270), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n273), .b(new_n283), .c(new_n282), .d(new_n256), .o1(new_n284));
  aoai13aa1n02x5               g189(.a(new_n275), .b(new_n284), .c(new_n181), .d(new_n271), .o1(new_n285));
  tech160nm_fiaoi012aa1n02p5x5 g190(.a(new_n280), .b(new_n285), .c(new_n278), .o1(new_n286));
  norp02aa1n03x5               g191(.a(new_n286), .b(new_n281), .o1(\s[28] ));
  norb02aa1n02x5               g192(.a(new_n275), .b(new_n280), .out0(new_n288));
  aobi12aa1n06x5               g193(.a(new_n288), .b(new_n272), .c(new_n274), .out0(new_n289));
  oao003aa1n02x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n278), .carry(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[28] ), .b(\a[29] ), .out0(new_n291));
  nano22aa1n03x7               g196(.a(new_n289), .b(new_n290), .c(new_n291), .out0(new_n292));
  aoai13aa1n02x5               g197(.a(new_n288), .b(new_n284), .c(new_n181), .d(new_n271), .o1(new_n293));
  tech160nm_fiaoi012aa1n02p5x5 g198(.a(new_n291), .b(new_n293), .c(new_n290), .o1(new_n294));
  norp02aa1n03x5               g199(.a(new_n294), .b(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g200(.a(new_n111), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g201(.a(new_n275), .b(new_n291), .c(new_n280), .out0(new_n297));
  aobi12aa1n06x5               g202(.a(new_n297), .b(new_n272), .c(new_n274), .out0(new_n298));
  oao003aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n299));
  xnrc02aa1n02x5               g204(.a(\b[29] ), .b(\a[30] ), .out0(new_n300));
  nano22aa1n03x7               g205(.a(new_n298), .b(new_n299), .c(new_n300), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n297), .b(new_n284), .c(new_n181), .d(new_n271), .o1(new_n302));
  tech160nm_fiaoi012aa1n02p5x5 g207(.a(new_n300), .b(new_n302), .c(new_n299), .o1(new_n303));
  norp02aa1n03x5               g208(.a(new_n303), .b(new_n301), .o1(\s[30] ));
  norb02aa1n02x7               g209(.a(new_n297), .b(new_n300), .out0(new_n305));
  aobi12aa1n06x5               g210(.a(new_n305), .b(new_n272), .c(new_n274), .out0(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n299), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[30] ), .b(\a[31] ), .out0(new_n308));
  nano22aa1n03x7               g213(.a(new_n306), .b(new_n307), .c(new_n308), .out0(new_n309));
  aoai13aa1n02x5               g214(.a(new_n305), .b(new_n284), .c(new_n181), .d(new_n271), .o1(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n308), .b(new_n310), .c(new_n307), .o1(new_n311));
  norp02aa1n03x5               g216(.a(new_n311), .b(new_n309), .o1(\s[31] ));
  xnbna2aa1n03x5               g217(.a(new_n113), .b(new_n116), .c(new_n119), .out0(\s[3] ));
  oaoi03aa1n02x5               g218(.a(\a[3] ), .b(\b[2] ), .c(new_n113), .o1(new_n314));
  xorb03aa1n02x5               g219(.a(new_n314), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g220(.a(new_n121), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g221(.a(new_n123), .b(new_n124), .c(new_n121), .o1(new_n317));
  xnrb03aa1n02x5               g222(.a(new_n317), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aobi12aa1n02x5               g223(.a(new_n125), .b(new_n121), .c(new_n108), .out0(new_n319));
  xnrb03aa1n02x5               g224(.a(new_n319), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g225(.a(\a[7] ), .b(\b[6] ), .c(new_n319), .o1(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g227(.a(new_n150), .b(new_n127), .c(new_n98), .out0(\s[9] ));
endmodule


