// Benchmark "adder" written by ABC on Thu Jul 18 14:51:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n347, new_n349, new_n350, new_n353, new_n354,
    new_n355, new_n356, new_n358, new_n360, new_n361, new_n363;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nor022aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n09x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand22aa1n03x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norb03aa1n12x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  oai012aa1n12x5               g007(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .o1(new_n103));
  nand42aa1n04x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  tech160nm_finand02aa1n03p5x5 g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nor002aa1n12x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nanb03aa1n09x5               g011(.a(new_n106), .b(new_n104), .c(new_n105), .out0(new_n107));
  nor002aa1n02x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  aoi012aa1n06x5               g013(.a(new_n106), .b(new_n108), .c(new_n104), .o1(new_n109));
  oai013aa1d12x5               g014(.a(new_n109), .b(new_n102), .c(new_n107), .d(new_n103), .o1(new_n110));
  xorc02aa1n06x5               g015(.a(\a[5] ), .b(\b[4] ), .out0(new_n111));
  xorc02aa1n02x5               g016(.a(\a[8] ), .b(\b[7] ), .out0(new_n112));
  norp02aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  and002aa1n03x5               g018(.a(\b[5] ), .b(\a[6] ), .o(new_n114));
  norp02aa1n06x5               g019(.a(new_n114), .b(new_n113), .o1(new_n115));
  nor042aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  and002aa1n12x5               g021(.a(\b[6] ), .b(\a[7] ), .o(new_n117));
  nona22aa1n02x4               g022(.a(new_n115), .b(new_n116), .c(new_n117), .out0(new_n118));
  nano22aa1n06x5               g023(.a(new_n118), .b(new_n111), .c(new_n112), .out0(new_n119));
  nanp02aa1n02x5               g024(.a(\b[7] ), .b(\a[8] ), .o1(new_n120));
  oai022aa1n04x7               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  aoi112aa1n09x5               g026(.a(new_n117), .b(new_n116), .c(\a[6] ), .d(\b[5] ), .o1(new_n122));
  oai022aa1n02x5               g027(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n120), .b(new_n123), .c(new_n122), .d(new_n121), .o1(new_n124));
  inv000aa1n04x5               g029(.a(new_n124), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoai13aa1n06x5               g031(.a(new_n126), .b(new_n125), .c(new_n110), .d(new_n119), .o1(new_n127));
  nor042aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand42aa1n06x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  norb02aa1n06x5               g034(.a(new_n129), .b(new_n128), .out0(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n130), .b(new_n127), .c(new_n98), .out0(\s[10] ));
  nona22aa1n06x5               g036(.a(new_n127), .b(new_n128), .c(new_n97), .out0(new_n132));
  nand42aa1n16x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor042aa1n04x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nanb03aa1n02x5               g039(.a(new_n134), .b(new_n129), .c(new_n133), .out0(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n133), .out0(new_n136));
  inv040aa1n02x5               g041(.a(new_n102), .o1(new_n137));
  nona22aa1n09x5               g042(.a(new_n137), .b(new_n107), .c(new_n103), .out0(new_n138));
  xnrc02aa1n02x5               g043(.a(\b[7] ), .b(\a[8] ), .out0(new_n139));
  xnrc02aa1n02x5               g044(.a(\b[6] ), .b(\a[7] ), .out0(new_n140));
  nona23aa1n06x5               g045(.a(new_n115), .b(new_n111), .c(new_n140), .d(new_n139), .out0(new_n141));
  aoai13aa1n12x5               g046(.a(new_n124), .b(new_n141), .c(new_n138), .d(new_n109), .o1(new_n142));
  oai022aa1n02x5               g047(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n129), .b(new_n143), .c(new_n142), .d(new_n126), .o1(new_n144));
  aboi22aa1n03x5               g049(.a(new_n135), .b(new_n132), .c(new_n144), .d(new_n136), .out0(\s[11] ));
  obai22aa1n02x7               g050(.a(new_n132), .b(new_n135), .c(\a[11] ), .d(\b[10] ), .out0(new_n146));
  norp02aa1n04x5               g051(.a(\b[11] ), .b(\a[12] ), .o1(new_n147));
  nand42aa1n08x5               g052(.a(\b[11] ), .b(\a[12] ), .o1(new_n148));
  norb02aa1n02x5               g053(.a(new_n148), .b(new_n147), .out0(new_n149));
  aoi113aa1n02x5               g054(.a(new_n149), .b(new_n134), .c(new_n132), .d(new_n133), .e(new_n129), .o1(new_n150));
  aoi012aa1n03x5               g055(.a(new_n150), .b(new_n146), .c(new_n149), .o1(\s[12] ));
  nano23aa1n06x5               g056(.a(new_n147), .b(new_n134), .c(new_n148), .d(new_n133), .out0(new_n152));
  nand23aa1d12x5               g057(.a(new_n152), .b(new_n126), .c(new_n130), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n125), .c(new_n110), .d(new_n119), .o1(new_n155));
  nano22aa1n03x5               g060(.a(new_n147), .b(new_n133), .c(new_n148), .out0(new_n156));
  tech160nm_fioai012aa1n03p5x5 g061(.a(new_n129), .b(\b[10] ), .c(\a[11] ), .o1(new_n157));
  oab012aa1n06x5               g062(.a(new_n157), .b(new_n97), .c(new_n128), .out0(new_n158));
  tech160nm_fiaoi012aa1n05x5   g063(.a(new_n147), .b(new_n134), .c(new_n148), .o1(new_n159));
  aob012aa1n02x5               g064(.a(new_n159), .b(new_n158), .c(new_n156), .out0(new_n160));
  nanb02aa1n03x5               g065(.a(new_n160), .b(new_n155), .out0(new_n161));
  nor022aa1n08x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand42aa1n04x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  inv030aa1n02x5               g069(.a(new_n159), .o1(new_n165));
  aoi112aa1n02x5               g070(.a(new_n165), .b(new_n164), .c(new_n158), .d(new_n156), .o1(new_n166));
  aoi022aa1n02x5               g071(.a(new_n161), .b(new_n164), .c(new_n155), .d(new_n166), .o1(\s[13] ));
  nor042aa1n04x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  nand42aa1n08x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  norb02aa1n02x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  aoai13aa1n04x5               g075(.a(new_n170), .b(new_n162), .c(new_n161), .d(new_n163), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n162), .b(new_n170), .c(new_n161), .d(new_n164), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[14] ));
  nano23aa1n09x5               g078(.a(new_n162), .b(new_n168), .c(new_n169), .d(new_n163), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n160), .c(new_n142), .d(new_n154), .o1(new_n175));
  oai012aa1n18x5               g080(.a(new_n169), .b(new_n168), .c(new_n162), .o1(new_n176));
  xorc02aa1n12x5               g081(.a(\a[15] ), .b(\b[14] ), .out0(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n175), .c(new_n176), .out0(\s[15] ));
  inv000aa1d42x5               g083(.a(new_n176), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n177), .b(new_n179), .c(new_n161), .d(new_n174), .o1(new_n180));
  nor042aa1n03x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n177), .o1(new_n183));
  aoai13aa1n02x5               g088(.a(new_n182), .b(new_n183), .c(new_n175), .d(new_n176), .o1(new_n184));
  tech160nm_fixorc02aa1n03p5x5 g089(.a(\a[16] ), .b(\b[15] ), .out0(new_n185));
  norp02aa1n02x5               g090(.a(new_n185), .b(new_n181), .o1(new_n186));
  aoi022aa1n02x5               g091(.a(new_n184), .b(new_n185), .c(new_n180), .d(new_n186), .o1(\s[16] ));
  nano32aa1d15x5               g092(.a(new_n153), .b(new_n185), .c(new_n174), .d(new_n177), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n125), .c(new_n110), .d(new_n119), .o1(new_n189));
  and002aa1n02x5               g094(.a(new_n185), .b(new_n177), .o(new_n190));
  aoai13aa1n06x5               g095(.a(new_n174), .b(new_n165), .c(new_n158), .d(new_n156), .o1(new_n191));
  aob012aa1n06x5               g096(.a(new_n190), .b(new_n191), .c(new_n176), .out0(new_n192));
  oao003aa1n02x5               g097(.a(\a[16] ), .b(\b[15] ), .c(new_n182), .carry(new_n193));
  nanp03aa1d12x5               g098(.a(new_n189), .b(new_n192), .c(new_n193), .o1(new_n194));
  xorc02aa1n03x5               g099(.a(\a[17] ), .b(\b[16] ), .out0(new_n195));
  nano22aa1n02x4               g100(.a(new_n195), .b(new_n192), .c(new_n193), .out0(new_n196));
  aoi022aa1n02x5               g101(.a(new_n196), .b(new_n189), .c(new_n194), .d(new_n195), .o1(\s[17] ));
  nor042aa1d18x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(new_n185), .b(new_n177), .o1(new_n200));
  aoai13aa1n06x5               g105(.a(new_n193), .b(new_n200), .c(new_n191), .d(new_n176), .o1(new_n201));
  aoai13aa1n03x5               g106(.a(new_n195), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n202));
  nor042aa1n09x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand02aa1n16x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  norb02aa1n06x4               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n202), .c(new_n199), .out0(\s[18] ));
  and002aa1n02x5               g111(.a(new_n195), .b(new_n205), .o(new_n207));
  aoai13aa1n03x5               g112(.a(new_n207), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n199), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor002aa1d32x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand02aa1n06x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n12x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n208), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g120(.a(new_n213), .b(new_n209), .c(new_n194), .d(new_n207), .o1(new_n216));
  inv000aa1d42x5               g121(.a(new_n211), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n213), .o1(new_n218));
  aoai13aa1n02x5               g123(.a(new_n217), .b(new_n218), .c(new_n208), .d(new_n210), .o1(new_n219));
  nor002aa1n16x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nand22aa1n12x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  norb02aa1n02x5               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  inv000aa1d42x5               g127(.a(\a[19] ), .o1(new_n223));
  inv000aa1d42x5               g128(.a(\b[18] ), .o1(new_n224));
  aboi22aa1n03x5               g129(.a(new_n220), .b(new_n221), .c(new_n223), .d(new_n224), .out0(new_n225));
  aoi022aa1n03x5               g130(.a(new_n219), .b(new_n222), .c(new_n216), .d(new_n225), .o1(\s[20] ));
  nano32aa1n03x7               g131(.a(new_n218), .b(new_n195), .c(new_n222), .d(new_n205), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n228));
  nanb03aa1n06x5               g133(.a(new_n220), .b(new_n221), .c(new_n212), .out0(new_n229));
  oai112aa1n06x5               g134(.a(new_n217), .b(new_n204), .c(new_n203), .d(new_n198), .o1(new_n230));
  aoi012aa1d18x5               g135(.a(new_n220), .b(new_n211), .c(new_n221), .o1(new_n231));
  oaih12aa1n12x5               g136(.a(new_n231), .b(new_n230), .c(new_n229), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  nanp02aa1n02x5               g138(.a(new_n228), .b(new_n233), .o1(new_n234));
  nor042aa1n12x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  nand42aa1n04x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n06x4               g141(.a(new_n236), .b(new_n235), .out0(new_n237));
  nano22aa1n03x7               g142(.a(new_n220), .b(new_n212), .c(new_n221), .out0(new_n238));
  oaih12aa1n02x5               g143(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .o1(new_n239));
  oab012aa1n03x5               g144(.a(new_n239), .b(new_n198), .c(new_n203), .out0(new_n240));
  inv000aa1n02x5               g145(.a(new_n231), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(new_n241), .b(new_n237), .c(new_n240), .d(new_n238), .o1(new_n242));
  aoi022aa1n02x5               g147(.a(new_n234), .b(new_n237), .c(new_n228), .d(new_n242), .o1(\s[21] ));
  aoai13aa1n03x5               g148(.a(new_n237), .b(new_n232), .c(new_n194), .d(new_n227), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n235), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n237), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n246), .c(new_n228), .d(new_n233), .o1(new_n247));
  nor042aa1n04x5               g152(.a(\b[21] ), .b(\a[22] ), .o1(new_n248));
  nand42aa1n16x5               g153(.a(\b[21] ), .b(\a[22] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  aoib12aa1n02x5               g155(.a(new_n235), .b(new_n249), .c(new_n248), .out0(new_n251));
  aoi022aa1n03x5               g156(.a(new_n247), .b(new_n250), .c(new_n244), .d(new_n251), .o1(\s[22] ));
  inv020aa1n02x5               g157(.a(new_n227), .o1(new_n253));
  nano22aa1n02x5               g158(.a(new_n253), .b(new_n237), .c(new_n250), .out0(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n255));
  nano23aa1d12x5               g160(.a(new_n235), .b(new_n248), .c(new_n249), .d(new_n236), .out0(new_n256));
  aoi012aa1d18x5               g161(.a(new_n248), .b(new_n235), .c(new_n249), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  tech160nm_fiaoi012aa1n03p5x5 g163(.a(new_n258), .b(new_n232), .c(new_n256), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(new_n255), .b(new_n259), .o1(new_n260));
  xorc02aa1n12x5               g165(.a(\a[23] ), .b(\b[22] ), .out0(new_n261));
  aoi112aa1n02x5               g166(.a(new_n261), .b(new_n258), .c(new_n232), .d(new_n256), .o1(new_n262));
  aoi022aa1n02x5               g167(.a(new_n260), .b(new_n261), .c(new_n255), .d(new_n262), .o1(\s[23] ));
  inv000aa1n02x5               g168(.a(new_n259), .o1(new_n264));
  aoai13aa1n03x5               g169(.a(new_n261), .b(new_n264), .c(new_n194), .d(new_n254), .o1(new_n265));
  nor042aa1n06x5               g170(.a(\b[22] ), .b(\a[23] ), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n266), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n261), .o1(new_n268));
  aoai13aa1n03x5               g173(.a(new_n267), .b(new_n268), .c(new_n255), .d(new_n259), .o1(new_n269));
  tech160nm_fixorc02aa1n02p5x5 g174(.a(\a[24] ), .b(\b[23] ), .out0(new_n270));
  norp02aa1n02x5               g175(.a(new_n270), .b(new_n266), .o1(new_n271));
  aoi022aa1n02x7               g176(.a(new_n269), .b(new_n270), .c(new_n265), .d(new_n271), .o1(\s[24] ));
  and002aa1n12x5               g177(.a(new_n270), .b(new_n261), .o(new_n273));
  nano22aa1n02x4               g178(.a(new_n253), .b(new_n273), .c(new_n256), .out0(new_n274));
  aoai13aa1n03x5               g179(.a(new_n274), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n256), .b(new_n241), .c(new_n240), .d(new_n238), .o1(new_n276));
  inv000aa1n06x5               g181(.a(new_n273), .o1(new_n277));
  oao003aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .carry(new_n278));
  aoai13aa1n12x5               g183(.a(new_n278), .b(new_n277), .c(new_n276), .d(new_n257), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(new_n275), .b(new_n280), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[25] ), .b(\b[24] ), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n273), .b(new_n258), .c(new_n232), .d(new_n256), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n282), .o1(new_n284));
  and003aa1n02x5               g189(.a(new_n283), .b(new_n284), .c(new_n278), .o(new_n285));
  aoi022aa1n02x5               g190(.a(new_n281), .b(new_n282), .c(new_n275), .d(new_n285), .o1(\s[25] ));
  aoai13aa1n03x5               g191(.a(new_n282), .b(new_n279), .c(new_n194), .d(new_n274), .o1(new_n287));
  nor042aa1n03x5               g192(.a(\b[24] ), .b(\a[25] ), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n289), .b(new_n284), .c(new_n275), .d(new_n280), .o1(new_n290));
  tech160nm_fixorc02aa1n02p5x5 g195(.a(\a[26] ), .b(\b[25] ), .out0(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n288), .o1(new_n292));
  aoi022aa1n02x7               g197(.a(new_n290), .b(new_n291), .c(new_n287), .d(new_n292), .o1(\s[26] ));
  and002aa1n12x5               g198(.a(new_n291), .b(new_n282), .o(new_n294));
  nano32aa1n03x7               g199(.a(new_n253), .b(new_n294), .c(new_n256), .d(new_n273), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n201), .c(new_n142), .d(new_n188), .o1(new_n296));
  oao003aa1n02x5               g201(.a(\a[26] ), .b(\b[25] ), .c(new_n289), .carry(new_n297));
  inv000aa1d42x5               g202(.a(new_n297), .o1(new_n298));
  aoi012aa1d18x5               g203(.a(new_n298), .b(new_n279), .c(new_n294), .o1(new_n299));
  nanp02aa1n02x5               g204(.a(new_n296), .b(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  aoi112aa1n02x5               g206(.a(new_n301), .b(new_n298), .c(new_n279), .d(new_n294), .o1(new_n302));
  aoi022aa1n02x5               g207(.a(new_n300), .b(new_n301), .c(new_n296), .d(new_n302), .o1(\s[27] ));
  inv000aa1d42x5               g208(.a(new_n294), .o1(new_n304));
  aoai13aa1n04x5               g209(.a(new_n297), .b(new_n304), .c(new_n283), .d(new_n278), .o1(new_n305));
  aoai13aa1n03x5               g210(.a(new_n301), .b(new_n305), .c(new_n194), .d(new_n295), .o1(new_n306));
  norp02aa1n02x5               g211(.a(\b[26] ), .b(\a[27] ), .o1(new_n307));
  inv000aa1n03x5               g212(.a(new_n307), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n301), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n308), .b(new_n309), .c(new_n296), .d(new_n299), .o1(new_n310));
  tech160nm_fixorc02aa1n03p5x5 g215(.a(\a[28] ), .b(\b[27] ), .out0(new_n311));
  norp02aa1n02x5               g216(.a(new_n311), .b(new_n307), .o1(new_n312));
  aoi022aa1n03x5               g217(.a(new_n310), .b(new_n311), .c(new_n306), .d(new_n312), .o1(\s[28] ));
  and002aa1n02x5               g218(.a(new_n311), .b(new_n301), .o(new_n314));
  aoai13aa1n03x5               g219(.a(new_n314), .b(new_n305), .c(new_n194), .d(new_n295), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n314), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[28] ), .b(\b[27] ), .c(new_n308), .carry(new_n317));
  aoai13aa1n03x5               g222(.a(new_n317), .b(new_n316), .c(new_n296), .d(new_n299), .o1(new_n318));
  tech160nm_fixorc02aa1n03p5x5 g223(.a(\a[29] ), .b(\b[28] ), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n317), .b(new_n319), .out0(new_n320));
  aoi022aa1n03x5               g225(.a(new_n318), .b(new_n319), .c(new_n315), .d(new_n320), .o1(\s[29] ));
  xorb03aa1n02x5               g226(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g227(.a(new_n309), .b(new_n311), .c(new_n319), .out0(new_n323));
  aoai13aa1n02x5               g228(.a(new_n323), .b(new_n305), .c(new_n194), .d(new_n295), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  inv000aa1d42x5               g230(.a(\b[28] ), .o1(new_n326));
  inv000aa1d42x5               g231(.a(\a[29] ), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n317), .b(\b[28] ), .c(new_n327), .out0(new_n328));
  oaib12aa1n02x5               g233(.a(new_n328), .b(new_n326), .c(\a[29] ), .out0(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n325), .c(new_n296), .d(new_n299), .o1(new_n330));
  tech160nm_fixorc02aa1n02p5x5 g235(.a(\a[30] ), .b(\b[29] ), .out0(new_n331));
  oaoi13aa1n02x5               g236(.a(new_n331), .b(new_n328), .c(new_n327), .d(new_n326), .o1(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n324), .d(new_n332), .o1(\s[30] ));
  nanb02aa1n02x5               g238(.a(\a[31] ), .b(\b[30] ), .out0(new_n334));
  nanb02aa1n02x5               g239(.a(\b[30] ), .b(\a[31] ), .out0(new_n335));
  nanp02aa1n02x5               g240(.a(new_n335), .b(new_n334), .o1(new_n336));
  nano32aa1n02x5               g241(.a(new_n309), .b(new_n331), .c(new_n311), .d(new_n319), .out0(new_n337));
  aoai13aa1n02x5               g242(.a(new_n337), .b(new_n305), .c(new_n194), .d(new_n295), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n337), .o1(new_n339));
  norp02aa1n02x5               g244(.a(\b[29] ), .b(\a[30] ), .o1(new_n340));
  aoi022aa1n02x5               g245(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n341));
  aoi012aa1n02x5               g246(.a(new_n340), .b(new_n328), .c(new_n341), .o1(new_n342));
  aoai13aa1n03x5               g247(.a(new_n342), .b(new_n339), .c(new_n296), .d(new_n299), .o1(new_n343));
  oai112aa1n02x5               g248(.a(new_n334), .b(new_n335), .c(\b[29] ), .d(\a[30] ), .o1(new_n344));
  aoi012aa1n02x5               g249(.a(new_n344), .b(new_n328), .c(new_n341), .o1(new_n345));
  aoi022aa1n03x5               g250(.a(new_n343), .b(new_n336), .c(new_n338), .d(new_n345), .o1(\s[31] ));
  norb02aa1n02x5               g251(.a(new_n105), .b(new_n108), .out0(new_n347));
  xobna2aa1n03x5               g252(.a(new_n347), .b(new_n137), .c(new_n100), .out0(\s[3] ));
  aoai13aa1n02x5               g253(.a(new_n347), .b(new_n102), .c(\a[2] ), .d(\b[1] ), .o1(new_n349));
  nanb02aa1n02x5               g254(.a(new_n106), .b(new_n104), .out0(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n350), .b(new_n349), .c(new_n105), .out0(\s[4] ));
  xnbna2aa1n03x5               g256(.a(new_n111), .b(new_n138), .c(new_n109), .out0(\s[5] ));
  norp02aa1n02x5               g257(.a(\b[4] ), .b(\a[5] ), .o1(new_n353));
  aoi012aa1n02x5               g258(.a(new_n353), .b(new_n110), .c(new_n111), .o1(new_n354));
  nanp02aa1n02x5               g259(.a(new_n110), .b(new_n111), .o1(new_n355));
  nona32aa1n02x4               g260(.a(new_n355), .b(new_n114), .c(new_n113), .d(new_n353), .out0(new_n356));
  oai012aa1n02x5               g261(.a(new_n356), .b(new_n354), .c(new_n115), .o1(\s[6] ));
  nanb02aa1n02x5               g262(.a(new_n114), .b(new_n356), .out0(new_n358));
  aoi022aa1n02x5               g263(.a(new_n358), .b(new_n140), .c(new_n122), .d(new_n356), .o1(\s[7] ));
  aoi012aa1n02x5               g264(.a(new_n116), .b(new_n356), .c(new_n122), .o1(new_n360));
  aoi112aa1n02x5               g265(.a(new_n112), .b(new_n116), .c(new_n356), .d(new_n122), .o1(new_n361));
  oab012aa1n02x4               g266(.a(new_n361), .b(new_n360), .c(new_n139), .out0(\s[8] ));
  aoi112aa1n02x5               g267(.a(new_n125), .b(new_n126), .c(new_n110), .d(new_n119), .o1(new_n363));
  aoi012aa1n02x5               g268(.a(new_n363), .b(new_n142), .c(new_n126), .o1(\s[9] ));
endmodule


