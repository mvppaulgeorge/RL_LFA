// Benchmark "adder" written by ABC on Thu Jul 18 03:05:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n339, new_n340, new_n342, new_n344, new_n346, new_n347, new_n349,
    new_n351, new_n352;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d48x5               g002(.a(\b[8] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv040aa1d32x5               g004(.a(\b[1] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oao003aa1n03x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .carry(new_n102));
  nand42aa1n20x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n06x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand42aa1n08x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano23aa1n02x5               g011(.a(new_n105), .b(new_n104), .c(new_n106), .d(new_n103), .out0(new_n107));
  nanp02aa1n03x5               g012(.a(new_n107), .b(new_n102), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\a[3] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(\b[2] ), .o1(new_n110));
  aoai13aa1n12x5               g015(.a(new_n103), .b(new_n104), .c(new_n110), .d(new_n109), .o1(new_n111));
  nor002aa1n20x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand22aa1n09x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nand22aa1n06x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nano23aa1n06x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nor002aa1d32x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nand02aa1n06x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nanb02aa1n12x5               g023(.a(new_n117), .b(new_n118), .out0(new_n119));
  nand42aa1n08x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nor022aa1n16x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nanb02aa1n12x5               g026(.a(new_n121), .b(new_n120), .out0(new_n122));
  nona22aa1n03x5               g027(.a(new_n116), .b(new_n119), .c(new_n122), .out0(new_n123));
  nona22aa1n09x5               g028(.a(new_n118), .b(new_n121), .c(new_n117), .out0(new_n124));
  oai112aa1n06x5               g029(.a(new_n120), .b(new_n113), .c(new_n114), .d(new_n112), .o1(new_n125));
  oa0012aa1n03x5               g030(.a(new_n118), .b(new_n121), .c(new_n117), .o(new_n126));
  oab012aa1n06x5               g031(.a(new_n126), .b(new_n125), .c(new_n124), .out0(new_n127));
  aoai13aa1n12x5               g032(.a(new_n127), .b(new_n123), .c(new_n108), .d(new_n111), .o1(new_n128));
  oaoi03aa1n02x5               g033(.a(new_n97), .b(new_n98), .c(new_n128), .o1(new_n129));
  xnrb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  tech160nm_fioaoi03aa1n04x5   g035(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n131));
  nona23aa1n09x5               g036(.a(new_n103), .b(new_n106), .c(new_n105), .d(new_n104), .out0(new_n132));
  oai012aa1n12x5               g037(.a(new_n111), .b(new_n132), .c(new_n131), .o1(new_n133));
  nona23aa1n09x5               g038(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n134));
  nor043aa1n06x5               g039(.a(new_n134), .b(new_n119), .c(new_n122), .o1(new_n135));
  oabi12aa1n06x5               g040(.a(new_n126), .b(new_n124), .c(new_n125), .out0(new_n136));
  nor002aa1d32x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  nanp02aa1n06x5               g042(.a(\b[9] ), .b(\a[10] ), .o1(new_n138));
  nor042aa1n03x5               g043(.a(\b[8] ), .b(\a[9] ), .o1(new_n139));
  nanp02aa1n04x5               g044(.a(\b[8] ), .b(\a[9] ), .o1(new_n140));
  nano23aa1n06x5               g045(.a(new_n137), .b(new_n139), .c(new_n140), .d(new_n138), .out0(new_n141));
  aoai13aa1n02x5               g046(.a(new_n141), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n142));
  aoai13aa1n06x5               g047(.a(new_n138), .b(new_n137), .c(new_n97), .d(new_n98), .o1(new_n143));
  nor042aa1n04x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nand02aa1d24x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n142), .c(new_n143), .out0(\s[11] ));
  inv000aa1n03x5               g052(.a(new_n144), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n145), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n148), .b(new_n149), .c(new_n142), .d(new_n143), .o1(new_n150));
  xorb03aa1n02x5               g055(.a(new_n150), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n09x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  nand02aa1n10x5               g057(.a(\b[11] ), .b(\a[12] ), .o1(new_n153));
  nano23aa1n06x5               g058(.a(new_n144), .b(new_n152), .c(new_n153), .d(new_n145), .out0(new_n154));
  and002aa1n02x5               g059(.a(new_n154), .b(new_n141), .o(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n152), .o1(new_n157));
  aoai13aa1n12x5               g062(.a(new_n157), .b(new_n149), .c(new_n143), .d(new_n148), .o1(new_n158));
  and002aa1n02x5               g063(.a(new_n158), .b(new_n153), .o(new_n159));
  inv040aa1n03x5               g064(.a(new_n159), .o1(new_n160));
  nor042aa1n06x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nand22aa1n09x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n160), .c(new_n156), .out0(\s[13] ));
  inv000aa1d42x5               g069(.a(\a[13] ), .o1(new_n165));
  inv000aa1d42x5               g070(.a(\b[12] ), .o1(new_n166));
  nanp02aa1n02x5               g071(.a(new_n160), .b(new_n156), .o1(new_n167));
  oaoi03aa1n03x5               g072(.a(new_n165), .b(new_n166), .c(new_n167), .o1(new_n168));
  xnrb03aa1n03x5               g073(.a(new_n168), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n20x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand22aa1n12x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  nona23aa1n09x5               g076(.a(new_n171), .b(new_n162), .c(new_n161), .d(new_n170), .out0(new_n172));
  aoai13aa1n02x5               g077(.a(new_n171), .b(new_n170), .c(new_n165), .d(new_n166), .o1(new_n173));
  aoai13aa1n06x5               g078(.a(new_n173), .b(new_n172), .c(new_n160), .d(new_n156), .o1(new_n174));
  norp02aa1n24x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  nand02aa1n10x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  nano23aa1n06x5               g082(.a(new_n161), .b(new_n170), .c(new_n171), .d(new_n162), .out0(new_n178));
  oai022aa1d18x5               g083(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n179));
  aoi122aa1n02x5               g084(.a(new_n177), .b(new_n171), .c(new_n179), .d(new_n167), .e(new_n178), .o1(new_n180));
  aoi012aa1n02x5               g085(.a(new_n180), .b(new_n174), .c(new_n177), .o1(\s[15] ));
  nor002aa1n16x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nanp02aa1n04x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nanb02aa1n02x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  aoai13aa1n02x5               g089(.a(new_n184), .b(new_n175), .c(new_n174), .d(new_n176), .o1(new_n185));
  aoi112aa1n03x4               g090(.a(new_n175), .b(new_n184), .c(new_n174), .d(new_n176), .o1(new_n186));
  nanb02aa1n03x5               g091(.a(new_n186), .b(new_n185), .out0(\s[16] ));
  nano23aa1n03x7               g092(.a(new_n175), .b(new_n182), .c(new_n183), .d(new_n176), .out0(new_n188));
  nand02aa1d04x5               g093(.a(new_n188), .b(new_n178), .o1(new_n189));
  nano22aa1d15x5               g094(.a(new_n189), .b(new_n141), .c(new_n154), .out0(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n191));
  nona23aa1n03x5               g096(.a(new_n183), .b(new_n176), .c(new_n175), .d(new_n182), .out0(new_n192));
  nor042aa1n06x5               g097(.a(new_n192), .b(new_n172), .o1(new_n193));
  aoai13aa1n03x5               g098(.a(new_n176), .b(new_n175), .c(new_n179), .d(new_n171), .o1(new_n194));
  tech160nm_fioaoi03aa1n04x5   g099(.a(\a[16] ), .b(\b[15] ), .c(new_n194), .o1(new_n195));
  aoi013aa1n06x4               g100(.a(new_n195), .b(new_n158), .c(new_n193), .d(new_n153), .o1(new_n196));
  nanp02aa1n06x5               g101(.a(new_n191), .b(new_n196), .o1(new_n197));
  nor042aa1n06x5               g102(.a(\b[16] ), .b(\a[17] ), .o1(new_n198));
  nand42aa1n06x5               g103(.a(\b[16] ), .b(\a[17] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  aoi113aa1n02x5               g105(.a(new_n200), .b(new_n195), .c(new_n158), .d(new_n193), .e(new_n153), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n197), .b(new_n200), .c(new_n191), .d(new_n201), .o1(\s[17] ));
  tech160nm_fiaoi012aa1n05x5   g107(.a(new_n198), .b(new_n197), .c(new_n200), .o1(new_n203));
  xnrb03aa1n03x5               g108(.a(new_n203), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp03aa1n06x5               g109(.a(new_n158), .b(new_n193), .c(new_n153), .o1(new_n205));
  nanb02aa1n12x5               g110(.a(new_n195), .b(new_n205), .out0(new_n206));
  nor042aa1n06x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  nand42aa1n10x5               g112(.a(\b[17] ), .b(\a[18] ), .o1(new_n208));
  nano23aa1d15x5               g113(.a(new_n198), .b(new_n207), .c(new_n208), .d(new_n199), .out0(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n206), .c(new_n128), .d(new_n190), .o1(new_n210));
  oa0012aa1n06x5               g115(.a(new_n208), .b(new_n207), .c(new_n198), .o(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor042aa1n04x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand42aa1n06x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n06x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n210), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp02aa1n02x5               g122(.a(new_n210), .b(new_n212), .o1(new_n218));
  nor022aa1n16x5               g123(.a(\b[19] ), .b(\a[20] ), .o1(new_n219));
  nand22aa1n12x5               g124(.a(\b[19] ), .b(\a[20] ), .o1(new_n220));
  nanb02aa1n06x5               g125(.a(new_n219), .b(new_n220), .out0(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n213), .c(new_n218), .d(new_n214), .o1(new_n222));
  aoai13aa1n03x5               g127(.a(new_n215), .b(new_n211), .c(new_n197), .d(new_n209), .o1(new_n223));
  nona22aa1n02x4               g128(.a(new_n223), .b(new_n221), .c(new_n213), .out0(new_n224));
  nanp02aa1n02x5               g129(.a(new_n222), .b(new_n224), .o1(\s[20] ));
  nanb03aa1d24x5               g130(.a(new_n219), .b(new_n220), .c(new_n214), .out0(new_n226));
  oaih22aa1d12x5               g131(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\b[18] ), .o1(new_n228));
  nanb02aa1n12x5               g133(.a(\a[19] ), .b(new_n228), .out0(new_n229));
  nand23aa1n09x5               g134(.a(new_n227), .b(new_n229), .c(new_n208), .o1(new_n230));
  aoi012aa1n09x5               g135(.a(new_n219), .b(new_n213), .c(new_n220), .o1(new_n231));
  oai012aa1d24x5               g136(.a(new_n231), .b(new_n230), .c(new_n226), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  nanb03aa1d18x5               g138(.a(new_n221), .b(new_n209), .c(new_n215), .out0(new_n234));
  aoai13aa1n06x5               g139(.a(new_n233), .b(new_n234), .c(new_n191), .d(new_n196), .o1(new_n235));
  xnrc02aa1n12x5               g140(.a(\b[20] ), .b(\a[21] ), .out0(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  inv040aa1n06x5               g142(.a(new_n234), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n237), .b(new_n197), .c(new_n238), .o1(new_n239));
  aoi022aa1n02x5               g144(.a(new_n239), .b(new_n233), .c(new_n235), .d(new_n237), .o1(\s[21] ));
  nor042aa1n03x5               g145(.a(\b[20] ), .b(\a[21] ), .o1(new_n241));
  tech160nm_fixnrc02aa1n04x5   g146(.a(\b[21] ), .b(\a[22] ), .out0(new_n242));
  aoai13aa1n02x5               g147(.a(new_n242), .b(new_n241), .c(new_n235), .d(new_n237), .o1(new_n243));
  aoi112aa1n03x5               g148(.a(new_n241), .b(new_n242), .c(new_n235), .d(new_n237), .o1(new_n244));
  nanb02aa1n03x5               g149(.a(new_n244), .b(new_n243), .out0(\s[22] ));
  nor042aa1n06x5               g150(.a(new_n242), .b(new_n236), .o1(new_n246));
  inv020aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  nor042aa1n02x5               g152(.a(new_n234), .b(new_n247), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n206), .c(new_n128), .d(new_n190), .o1(new_n249));
  inv000aa1d42x5               g154(.a(\a[22] ), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[21] ), .o1(new_n251));
  oaoi03aa1n09x5               g156(.a(new_n250), .b(new_n251), .c(new_n241), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  aoi012aa1n02x5               g158(.a(new_n253), .b(new_n232), .c(new_n246), .o1(new_n254));
  nand02aa1d04x5               g159(.a(new_n249), .b(new_n254), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[23] ), .b(\b[22] ), .out0(new_n256));
  aoi112aa1n02x5               g161(.a(new_n256), .b(new_n253), .c(new_n232), .d(new_n246), .o1(new_n257));
  aoi022aa1n02x5               g162(.a(new_n255), .b(new_n256), .c(new_n249), .d(new_n257), .o1(\s[23] ));
  norp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  xnrc02aa1n12x5               g164(.a(\b[23] ), .b(\a[24] ), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n259), .c(new_n255), .d(new_n256), .o1(new_n261));
  nand02aa1d04x5               g166(.a(new_n255), .b(new_n256), .o1(new_n262));
  nona22aa1n03x5               g167(.a(new_n262), .b(new_n260), .c(new_n259), .out0(new_n263));
  nanp02aa1n03x5               g168(.a(new_n263), .b(new_n261), .o1(\s[24] ));
  nanb02aa1n09x5               g169(.a(new_n260), .b(new_n256), .out0(new_n265));
  nor043aa1n03x5               g170(.a(new_n234), .b(new_n247), .c(new_n265), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n266), .b(new_n206), .c(new_n128), .d(new_n190), .o1(new_n267));
  nano22aa1n03x5               g172(.a(new_n219), .b(new_n214), .c(new_n220), .out0(new_n268));
  oai012aa1n02x5               g173(.a(new_n208), .b(\b[18] ), .c(\a[19] ), .o1(new_n269));
  oab012aa1n02x5               g174(.a(new_n269), .b(new_n198), .c(new_n207), .out0(new_n270));
  inv040aa1n02x5               g175(.a(new_n231), .o1(new_n271));
  aoai13aa1n06x5               g176(.a(new_n246), .b(new_n271), .c(new_n270), .d(new_n268), .o1(new_n272));
  aoi112aa1n02x5               g177(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n273));
  oab012aa1n02x4               g178(.a(new_n273), .b(\a[24] ), .c(\b[23] ), .out0(new_n274));
  aoai13aa1n04x5               g179(.a(new_n274), .b(new_n265), .c(new_n272), .d(new_n252), .o1(new_n275));
  nanb02aa1n06x5               g180(.a(new_n275), .b(new_n267), .out0(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  inv000aa1n02x5               g182(.a(new_n265), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n253), .c(new_n232), .d(new_n246), .o1(new_n279));
  nano22aa1n02x4               g184(.a(new_n277), .b(new_n279), .c(new_n274), .out0(new_n280));
  aoi022aa1n02x5               g185(.a(new_n276), .b(new_n277), .c(new_n267), .d(new_n280), .o1(\s[25] ));
  nor002aa1n02x5               g186(.a(\b[24] ), .b(\a[25] ), .o1(new_n282));
  tech160nm_fixnrc02aa1n04x5   g187(.a(\b[25] ), .b(\a[26] ), .out0(new_n283));
  aoai13aa1n02x5               g188(.a(new_n283), .b(new_n282), .c(new_n276), .d(new_n277), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n277), .b(new_n275), .c(new_n197), .d(new_n266), .o1(new_n285));
  nona22aa1n02x4               g190(.a(new_n285), .b(new_n283), .c(new_n282), .out0(new_n286));
  nanp02aa1n03x5               g191(.a(new_n284), .b(new_n286), .o1(\s[26] ));
  norb02aa1n12x5               g192(.a(new_n277), .b(new_n283), .out0(new_n288));
  nano23aa1n03x7               g193(.a(new_n234), .b(new_n265), .c(new_n288), .d(new_n246), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n206), .c(new_n128), .d(new_n190), .o1(new_n290));
  inv000aa1d42x5               g195(.a(\a[26] ), .o1(new_n291));
  inv000aa1d42x5               g196(.a(\b[25] ), .o1(new_n292));
  oaoi03aa1n02x5               g197(.a(new_n291), .b(new_n292), .c(new_n282), .o1(new_n293));
  inv000aa1n02x5               g198(.a(new_n293), .o1(new_n294));
  tech160nm_fiaoi012aa1n05x5   g199(.a(new_n294), .b(new_n275), .c(new_n288), .o1(new_n295));
  nand42aa1n02x5               g200(.a(new_n295), .b(new_n290), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[27] ), .b(\b[26] ), .out0(new_n297));
  aoi112aa1n02x5               g202(.a(new_n297), .b(new_n294), .c(new_n275), .d(new_n288), .o1(new_n298));
  aoi022aa1n02x5               g203(.a(new_n296), .b(new_n297), .c(new_n290), .d(new_n298), .o1(\s[27] ));
  norp02aa1n02x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  norp02aa1n02x5               g205(.a(\b[27] ), .b(\a[28] ), .o1(new_n301));
  nanp02aa1n02x5               g206(.a(\b[27] ), .b(\a[28] ), .o1(new_n302));
  norb02aa1n09x5               g207(.a(new_n302), .b(new_n301), .out0(new_n303));
  inv000aa1d42x5               g208(.a(new_n303), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n300), .c(new_n296), .d(new_n297), .o1(new_n305));
  nona23aa1n03x5               g210(.a(new_n238), .b(new_n288), .c(new_n265), .d(new_n247), .out0(new_n306));
  aoi012aa1n06x5               g211(.a(new_n306), .b(new_n191), .c(new_n196), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n288), .o1(new_n308));
  aoai13aa1n06x5               g213(.a(new_n293), .b(new_n308), .c(new_n279), .d(new_n274), .o1(new_n309));
  oaih12aa1n02x5               g214(.a(new_n297), .b(new_n309), .c(new_n307), .o1(new_n310));
  nona22aa1n02x5               g215(.a(new_n310), .b(new_n304), .c(new_n300), .out0(new_n311));
  nanp02aa1n03x5               g216(.a(new_n305), .b(new_n311), .o1(\s[28] ));
  xnrc02aa1n02x5               g217(.a(\b[28] ), .b(\a[29] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n297), .b(new_n304), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n314), .b(new_n309), .c(new_n307), .o1(new_n315));
  oai012aa1n02x5               g220(.a(new_n302), .b(new_n301), .c(new_n300), .o1(new_n316));
  aoi012aa1n03x5               g221(.a(new_n313), .b(new_n315), .c(new_n316), .o1(new_n317));
  aobi12aa1n03x5               g222(.a(new_n314), .b(new_n295), .c(new_n290), .out0(new_n318));
  nano22aa1n02x4               g223(.a(new_n318), .b(new_n313), .c(new_n316), .out0(new_n319));
  norp02aa1n03x5               g224(.a(new_n317), .b(new_n319), .o1(\s[29] ));
  xorb03aa1n02x5               g225(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g226(.a(new_n313), .b(new_n297), .c(new_n303), .out0(new_n322));
  oaih12aa1n02x5               g227(.a(new_n322), .b(new_n309), .c(new_n307), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[29] ), .b(\b[28] ), .c(new_n316), .carry(new_n324));
  nanp02aa1n03x5               g229(.a(new_n323), .b(new_n324), .o1(new_n325));
  xorc02aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .out0(new_n326));
  norb02aa1n02x5               g231(.a(new_n324), .b(new_n326), .out0(new_n327));
  aoi022aa1n02x7               g232(.a(new_n325), .b(new_n326), .c(new_n323), .d(new_n327), .o1(\s[30] ));
  nona23aa1n02x4               g233(.a(new_n326), .b(new_n297), .c(new_n304), .d(new_n313), .out0(new_n329));
  oabi12aa1n02x5               g234(.a(new_n329), .b(new_n309), .c(new_n307), .out0(new_n330));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  and002aa1n02x5               g236(.a(\b[29] ), .b(\a[30] ), .o(new_n332));
  oabi12aa1n02x5               g237(.a(new_n331), .b(\a[30] ), .c(\b[29] ), .out0(new_n333));
  oab012aa1n02x4               g238(.a(new_n333), .b(new_n324), .c(new_n332), .out0(new_n334));
  oao003aa1n02x5               g239(.a(\a[30] ), .b(\b[29] ), .c(new_n324), .carry(new_n335));
  aoai13aa1n03x5               g240(.a(new_n335), .b(new_n329), .c(new_n295), .d(new_n290), .o1(new_n336));
  aoi022aa1n02x5               g241(.a(new_n336), .b(new_n331), .c(new_n330), .d(new_n334), .o1(\s[31] ));
  xorb03aa1n02x5               g242(.a(new_n131), .b(\b[2] ), .c(new_n109), .out0(\s[3] ));
  norb02aa1n02x5               g243(.a(new_n103), .b(new_n104), .out0(new_n339));
  aoi112aa1n02x5               g244(.a(new_n105), .b(new_n339), .c(new_n102), .d(new_n106), .o1(new_n340));
  aoib12aa1n02x5               g245(.a(new_n340), .b(new_n133), .c(new_n104), .out0(\s[4] ));
  nanb02aa1n02x5               g246(.a(new_n114), .b(new_n115), .out0(new_n342));
  xobna2aa1n03x5               g247(.a(new_n342), .b(new_n108), .c(new_n111), .out0(\s[5] ));
  aoi012aa1n02x5               g248(.a(new_n114), .b(new_n133), .c(new_n115), .o1(new_n344));
  xnrb03aa1n02x5               g249(.a(new_n344), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oa0012aa1n02x5               g250(.a(new_n113), .b(new_n114), .c(new_n112), .o(new_n346));
  tech160nm_fiao0012aa1n02p5x5 g251(.a(new_n346), .b(new_n133), .c(new_n116), .o(new_n347));
  xorb03aa1n02x5               g252(.a(new_n347), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g253(.a(new_n121), .b(new_n347), .c(new_n120), .o1(new_n349));
  xnrb03aa1n02x5               g254(.a(new_n349), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  norb02aa1n02x5               g255(.a(new_n140), .b(new_n139), .out0(new_n351));
  aoi112aa1n02x5               g256(.a(new_n351), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n352));
  aoi012aa1n02x5               g257(.a(new_n352), .b(new_n128), .c(new_n351), .o1(\s[9] ));
endmodule


