// Benchmark "adder" written by ABC on Wed Jul 17 22:04:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n141, new_n142, new_n143, new_n144, new_n145, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n342, new_n343, new_n345, new_n347,
    new_n348, new_n350, new_n351, new_n353, new_n354, new_n355, new_n357;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  nor002aa1n04x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nand42aa1n08x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nand02aa1d06x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norb03aa1d15x5               g006(.a(new_n100), .b(new_n99), .c(new_n101), .out0(new_n102));
  inv040aa1n02x5               g007(.a(new_n102), .o1(new_n103));
  oai012aa1n04x7               g008(.a(new_n100), .b(\b[3] ), .c(\a[4] ), .o1(new_n104));
  tech160nm_finand02aa1n05x5   g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1n08x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nor042aa1n04x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nanb03aa1d18x5               g012(.a(new_n107), .b(new_n105), .c(new_n106), .out0(new_n108));
  nona22aa1n09x5               g013(.a(new_n103), .b(new_n108), .c(new_n104), .out0(new_n109));
  norp02aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  aoi012aa1n06x5               g015(.a(new_n110), .b(new_n107), .c(new_n106), .o1(new_n111));
  nand42aa1n06x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nor002aa1d32x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  norb02aa1n03x5               g018(.a(new_n112), .b(new_n113), .out0(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .out0(new_n115));
  xorc02aa1n12x5               g020(.a(\a[7] ), .b(\b[6] ), .out0(new_n116));
  xnrc02aa1n12x5               g021(.a(\b[4] ), .b(\a[5] ), .out0(new_n117));
  nona23aa1n09x5               g022(.a(new_n116), .b(new_n114), .c(new_n117), .d(new_n115), .out0(new_n118));
  inv000aa1d42x5               g023(.a(\a[8] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[7] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\a[7] ), .o1(new_n121));
  inv000aa1d42x5               g026(.a(\b[6] ), .o1(new_n122));
  nand22aa1n03x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  inv000aa1d42x5               g028(.a(\a[5] ), .o1(new_n124));
  inv000aa1d42x5               g029(.a(\b[4] ), .o1(new_n125));
  aoai13aa1n06x5               g030(.a(new_n112), .b(new_n113), .c(new_n125), .d(new_n124), .o1(new_n126));
  oai022aa1n06x5               g031(.a(new_n121), .b(new_n122), .c(new_n120), .d(new_n119), .o1(new_n127));
  tech160nm_fiaoi012aa1n05x5   g032(.a(new_n127), .b(new_n126), .c(new_n123), .o1(new_n128));
  aoi012aa1n12x5               g033(.a(new_n128), .b(new_n119), .c(new_n120), .o1(new_n129));
  aoai13aa1n12x5               g034(.a(new_n129), .b(new_n118), .c(new_n109), .d(new_n111), .o1(new_n130));
  xorc02aa1n12x5               g035(.a(\a[9] ), .b(\b[8] ), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n97), .b(new_n98), .c(new_n130), .d(new_n131), .o1(new_n132));
  oai013aa1n09x5               g037(.a(new_n111), .b(new_n102), .c(new_n108), .d(new_n104), .o1(new_n133));
  xorc02aa1n02x5               g038(.a(\a[8] ), .b(\b[7] ), .out0(new_n134));
  nano32aa1n03x7               g039(.a(new_n117), .b(new_n116), .c(new_n134), .d(new_n114), .out0(new_n135));
  inv040aa1n02x5               g040(.a(new_n129), .o1(new_n136));
  aoai13aa1n02x5               g041(.a(new_n131), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n137));
  norp02aa1n02x5               g042(.a(new_n97), .b(new_n98), .o1(new_n138));
  nanp02aa1n03x5               g043(.a(new_n137), .b(new_n138), .o1(new_n139));
  nanp02aa1n02x5               g044(.a(new_n132), .b(new_n139), .o1(\s[10] ));
  xnrc02aa1n12x5               g045(.a(\b[10] ), .b(\a[11] ), .out0(new_n141));
  aob012aa1n02x5               g046(.a(new_n139), .b(\b[9] ), .c(\a[10] ), .out0(new_n142));
  orn002aa1n02x5               g047(.a(\a[11] ), .b(\b[10] ), .o(new_n143));
  aoi022aa1d24x5               g048(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n144));
  and002aa1n02x5               g049(.a(new_n144), .b(new_n143), .o(new_n145));
  aoi022aa1n02x5               g050(.a(new_n142), .b(new_n141), .c(new_n139), .d(new_n145), .o1(\s[11] ));
  aob012aa1n02x5               g051(.a(new_n143), .b(new_n139), .c(new_n144), .out0(new_n147));
  xorc02aa1n12x5               g052(.a(\a[12] ), .b(\b[11] ), .out0(new_n148));
  nanb02aa1n02x5               g053(.a(new_n148), .b(new_n143), .out0(new_n149));
  aoi012aa1n02x5               g054(.a(new_n149), .b(new_n139), .c(new_n145), .o1(new_n150));
  aoi012aa1n02x5               g055(.a(new_n150), .b(new_n147), .c(new_n148), .o1(\s[12] ));
  nona23aa1d24x5               g056(.a(new_n148), .b(new_n131), .c(new_n97), .d(new_n141), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n02x5               g058(.a(new_n153), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n154));
  nanp02aa1n03x5               g059(.a(new_n135), .b(new_n133), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  oaih22aa1d12x5               g061(.a(\a[11] ), .b(\b[10] ), .c(\b[11] ), .d(\a[12] ), .o1(new_n157));
  oaih22aa1n04x5               g062(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n158));
  aoai13aa1n06x5               g063(.a(new_n156), .b(new_n157), .c(new_n158), .d(new_n144), .o1(new_n159));
  aoai13aa1n03x5               g064(.a(new_n159), .b(new_n152), .c(new_n155), .d(new_n129), .o1(new_n160));
  xnrc02aa1n12x5               g065(.a(\b[12] ), .b(\a[13] ), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  nano32aa1n02x4               g067(.a(new_n157), .b(new_n158), .c(new_n144), .d(new_n156), .out0(new_n163));
  aoi112aa1n02x5               g068(.a(new_n163), .b(new_n162), .c(new_n156), .d(new_n157), .o1(new_n164));
  aoi022aa1n02x5               g069(.a(new_n160), .b(new_n162), .c(new_n154), .d(new_n164), .o1(\s[13] ));
  orn002aa1n24x5               g070(.a(\a[13] ), .b(\b[12] ), .o(new_n166));
  inv000aa1n02x5               g071(.a(new_n157), .o1(new_n167));
  norp02aa1n02x5               g072(.a(\b[9] ), .b(\a[10] ), .o1(new_n168));
  oaih12aa1n02x5               g073(.a(new_n144), .b(new_n98), .c(new_n168), .o1(new_n169));
  aoi022aa1n06x5               g074(.a(new_n169), .b(new_n167), .c(\a[12] ), .d(\b[11] ), .o1(new_n170));
  aoai13aa1n03x5               g075(.a(new_n162), .b(new_n170), .c(new_n130), .d(new_n153), .o1(new_n171));
  tech160nm_fixnrc02aa1n05x5   g076(.a(\b[13] ), .b(\a[14] ), .out0(new_n172));
  xobna2aa1n03x5               g077(.a(new_n172), .b(new_n171), .c(new_n166), .out0(\s[14] ));
  norp02aa1n12x5               g078(.a(new_n172), .b(new_n161), .o1(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n170), .c(new_n130), .d(new_n153), .o1(new_n175));
  oao003aa1n12x5               g080(.a(\a[14] ), .b(\b[13] ), .c(new_n166), .carry(new_n176));
  tech160nm_fixorc02aa1n03p5x5 g081(.a(\a[15] ), .b(\b[14] ), .out0(new_n177));
  xnbna2aa1n03x5               g082(.a(new_n177), .b(new_n175), .c(new_n176), .out0(\s[15] ));
  inv040aa1n02x5               g083(.a(new_n176), .o1(new_n179));
  aoai13aa1n02x5               g084(.a(new_n177), .b(new_n179), .c(new_n160), .d(new_n174), .o1(new_n180));
  nor002aa1d24x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n181), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n177), .o1(new_n183));
  aoai13aa1n02x7               g088(.a(new_n182), .b(new_n183), .c(new_n175), .d(new_n176), .o1(new_n184));
  xorc02aa1n02x5               g089(.a(\a[16] ), .b(\b[15] ), .out0(new_n185));
  norp02aa1n02x5               g090(.a(new_n185), .b(new_n181), .o1(new_n186));
  aoi022aa1n03x5               g091(.a(new_n184), .b(new_n185), .c(new_n180), .d(new_n186), .o1(\s[16] ));
  nanp02aa1n02x5               g092(.a(\b[14] ), .b(\a[15] ), .o1(new_n188));
  xnrc02aa1n02x5               g093(.a(\b[15] ), .b(\a[16] ), .out0(new_n189));
  nano22aa1n03x7               g094(.a(new_n189), .b(new_n182), .c(new_n188), .out0(new_n190));
  nano22aa1d15x5               g095(.a(new_n152), .b(new_n174), .c(new_n190), .out0(new_n191));
  aoai13aa1n06x5               g096(.a(new_n191), .b(new_n136), .c(new_n133), .d(new_n135), .o1(new_n192));
  oai013aa1n02x4               g097(.a(new_n176), .b(new_n159), .c(new_n161), .d(new_n172), .o1(new_n193));
  oao003aa1n02x5               g098(.a(\a[16] ), .b(\b[15] ), .c(new_n182), .carry(new_n194));
  aobi12aa1n06x5               g099(.a(new_n194), .b(new_n193), .c(new_n190), .out0(new_n195));
  nanp02aa1n12x5               g100(.a(new_n192), .b(new_n195), .o1(new_n196));
  tech160nm_fixorc02aa1n05x5   g101(.a(\a[17] ), .b(\b[16] ), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n190), .b(new_n179), .c(new_n170), .d(new_n174), .o1(new_n198));
  nano22aa1n02x4               g103(.a(new_n197), .b(new_n198), .c(new_n194), .out0(new_n199));
  aoi022aa1n02x5               g104(.a(new_n196), .b(new_n197), .c(new_n192), .d(new_n199), .o1(\s[17] ));
  inv040aa1d32x5               g105(.a(\a[17] ), .o1(new_n201));
  inv040aa1d28x5               g106(.a(\b[16] ), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(new_n202), .b(new_n201), .o1(new_n203));
  nand22aa1n04x5               g108(.a(new_n198), .b(new_n194), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n197), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n205));
  nor042aa1n02x5               g110(.a(\b[17] ), .b(\a[18] ), .o1(new_n206));
  nand22aa1n04x5               g111(.a(\b[17] ), .b(\a[18] ), .o1(new_n207));
  norb02aa1n06x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  xnbna2aa1n03x5               g113(.a(new_n208), .b(new_n205), .c(new_n203), .out0(\s[18] ));
  and002aa1n02x5               g114(.a(new_n197), .b(new_n208), .o(new_n210));
  aoai13aa1n06x5               g115(.a(new_n210), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n211));
  aoi013aa1n09x5               g116(.a(new_n206), .b(new_n207), .c(new_n201), .d(new_n202), .o1(new_n212));
  nor002aa1d32x5               g117(.a(\b[18] ), .b(\a[19] ), .o1(new_n213));
  nand42aa1n20x5               g118(.a(\b[18] ), .b(\a[19] ), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n211), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g121(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_fioaoi03aa1n03p5x5 g122(.a(\a[18] ), .b(\b[17] ), .c(new_n203), .o1(new_n218));
  aoai13aa1n03x5               g123(.a(new_n215), .b(new_n218), .c(new_n196), .d(new_n210), .o1(new_n219));
  inv040aa1n08x5               g124(.a(new_n213), .o1(new_n220));
  inv000aa1n02x5               g125(.a(new_n215), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n220), .b(new_n221), .c(new_n211), .d(new_n212), .o1(new_n222));
  nor002aa1d32x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  nand02aa1n06x5               g128(.a(\b[19] ), .b(\a[20] ), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(new_n225));
  inv000aa1d42x5               g130(.a(\a[19] ), .o1(new_n226));
  inv000aa1d42x5               g131(.a(\b[18] ), .o1(new_n227));
  aboi22aa1n03x5               g132(.a(new_n223), .b(new_n224), .c(new_n226), .d(new_n227), .out0(new_n228));
  aoi022aa1n03x5               g133(.a(new_n222), .b(new_n225), .c(new_n219), .d(new_n228), .o1(\s[20] ));
  nona23aa1d18x5               g134(.a(new_n224), .b(new_n214), .c(new_n213), .d(new_n223), .out0(new_n230));
  nano22aa1n03x5               g135(.a(new_n230), .b(new_n197), .c(new_n208), .out0(new_n231));
  aoai13aa1n02x5               g136(.a(new_n231), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n232));
  inv000aa1n02x5               g137(.a(new_n231), .o1(new_n233));
  oaoi03aa1n12x5               g138(.a(\a[20] ), .b(\b[19] ), .c(new_n220), .o1(new_n234));
  inv040aa1n02x5               g139(.a(new_n234), .o1(new_n235));
  oai012aa1d24x5               g140(.a(new_n235), .b(new_n230), .c(new_n212), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n233), .c(new_n192), .d(new_n195), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[20] ), .b(\a[21] ), .out0(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  nano23aa1n03x7               g145(.a(new_n213), .b(new_n223), .c(new_n224), .d(new_n214), .out0(new_n241));
  aoi112aa1n02x5               g146(.a(new_n234), .b(new_n240), .c(new_n241), .d(new_n218), .o1(new_n242));
  aoi022aa1n02x5               g147(.a(new_n238), .b(new_n240), .c(new_n232), .d(new_n242), .o1(\s[21] ));
  nanp02aa1n02x5               g148(.a(new_n238), .b(new_n240), .o1(new_n244));
  nor042aa1n06x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  inv000aa1n03x5               g150(.a(new_n245), .o1(new_n246));
  aoai13aa1n02x7               g151(.a(new_n246), .b(new_n239), .c(new_n232), .d(new_n237), .o1(new_n247));
  xnrc02aa1n12x5               g152(.a(\b[21] ), .b(\a[22] ), .out0(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n248), .b(new_n245), .out0(new_n250));
  aoi022aa1n03x5               g155(.a(new_n247), .b(new_n249), .c(new_n244), .d(new_n250), .o1(\s[22] ));
  nor042aa1n06x5               g156(.a(new_n248), .b(new_n239), .o1(new_n252));
  nano32aa1n02x4               g157(.a(new_n230), .b(new_n252), .c(new_n197), .d(new_n208), .out0(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n252), .b(new_n234), .c(new_n241), .d(new_n218), .o1(new_n255));
  oao003aa1n12x5               g160(.a(\a[22] ), .b(\b[21] ), .c(new_n246), .carry(new_n256));
  nanp02aa1n03x5               g161(.a(new_n255), .b(new_n256), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[23] ), .b(\b[22] ), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n257), .c(new_n196), .d(new_n253), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n256), .o1(new_n260));
  aoi112aa1n02x5               g165(.a(new_n258), .b(new_n260), .c(new_n236), .d(new_n252), .o1(new_n261));
  aobi12aa1n02x7               g166(.a(new_n259), .b(new_n261), .c(new_n254), .out0(\s[23] ));
  inv000aa1n02x5               g167(.a(new_n257), .o1(new_n263));
  nor042aa1n09x5               g168(.a(\b[22] ), .b(\a[23] ), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n264), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n258), .o1(new_n266));
  aoai13aa1n03x5               g171(.a(new_n265), .b(new_n266), .c(new_n254), .d(new_n263), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[24] ), .b(\b[23] ), .out0(new_n268));
  norp02aa1n02x5               g173(.a(new_n268), .b(new_n264), .o1(new_n269));
  aoi022aa1n02x7               g174(.a(new_n267), .b(new_n268), .c(new_n259), .d(new_n269), .o1(\s[24] ));
  and002aa1n12x5               g175(.a(new_n268), .b(new_n258), .o(new_n271));
  nano22aa1n02x5               g176(.a(new_n233), .b(new_n271), .c(new_n252), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n273));
  inv000aa1n03x5               g178(.a(new_n271), .o1(new_n274));
  oao003aa1n02x5               g179(.a(\a[24] ), .b(\b[23] ), .c(new_n265), .carry(new_n275));
  aoai13aa1n12x5               g180(.a(new_n275), .b(new_n274), .c(new_n255), .d(new_n256), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[25] ), .b(\b[24] ), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n276), .c(new_n196), .d(new_n272), .o1(new_n278));
  aoai13aa1n04x5               g183(.a(new_n271), .b(new_n260), .c(new_n236), .d(new_n252), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n277), .o1(new_n280));
  and003aa1n02x5               g185(.a(new_n279), .b(new_n280), .c(new_n275), .o(new_n281));
  aobi12aa1n02x7               g186(.a(new_n278), .b(new_n281), .c(new_n273), .out0(\s[25] ));
  inv000aa1n02x5               g187(.a(new_n276), .o1(new_n283));
  nor042aa1n04x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  inv000aa1n03x5               g189(.a(new_n284), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n280), .c(new_n273), .d(new_n283), .o1(new_n286));
  xorc02aa1n02x5               g191(.a(\a[26] ), .b(\b[25] ), .out0(new_n287));
  norp02aa1n02x5               g192(.a(new_n287), .b(new_n284), .o1(new_n288));
  aoi022aa1n03x5               g193(.a(new_n286), .b(new_n287), .c(new_n278), .d(new_n288), .o1(\s[26] ));
  and002aa1n02x5               g194(.a(new_n287), .b(new_n277), .o(new_n290));
  inv000aa1n02x5               g195(.a(new_n290), .o1(new_n291));
  nano32aa1n03x7               g196(.a(new_n291), .b(new_n231), .c(new_n271), .d(new_n252), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n204), .c(new_n130), .d(new_n191), .o1(new_n293));
  tech160nm_fioaoi03aa1n02p5x5 g198(.a(\a[26] ), .b(\b[25] ), .c(new_n285), .o1(new_n294));
  inv000aa1n02x5               g199(.a(new_n294), .o1(new_n295));
  aoai13aa1n04x5               g200(.a(new_n295), .b(new_n291), .c(new_n279), .d(new_n275), .o1(new_n296));
  xorc02aa1n12x5               g201(.a(\a[27] ), .b(\b[26] ), .out0(new_n297));
  aoai13aa1n06x5               g202(.a(new_n297), .b(new_n296), .c(new_n196), .d(new_n292), .o1(new_n298));
  aoi112aa1n02x5               g203(.a(new_n297), .b(new_n294), .c(new_n276), .d(new_n290), .o1(new_n299));
  aobi12aa1n03x7               g204(.a(new_n298), .b(new_n299), .c(new_n293), .out0(\s[27] ));
  tech160nm_fiaoi012aa1n05x5   g205(.a(new_n294), .b(new_n276), .c(new_n290), .o1(new_n301));
  nor042aa1d18x5               g206(.a(\b[26] ), .b(\a[27] ), .o1(new_n302));
  inv040aa1n06x5               g207(.a(new_n302), .o1(new_n303));
  inv020aa1n03x5               g208(.a(new_n297), .o1(new_n304));
  aoai13aa1n06x5               g209(.a(new_n303), .b(new_n304), .c(new_n301), .d(new_n293), .o1(new_n305));
  xorc02aa1n12x5               g210(.a(\a[28] ), .b(\b[27] ), .out0(new_n306));
  norp02aa1n02x5               g211(.a(new_n306), .b(new_n302), .o1(new_n307));
  aoi022aa1n02x7               g212(.a(new_n305), .b(new_n306), .c(new_n298), .d(new_n307), .o1(\s[28] ));
  and002aa1n02x5               g213(.a(new_n306), .b(new_n297), .o(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n296), .c(new_n196), .d(new_n292), .o1(new_n310));
  inv000aa1d42x5               g215(.a(new_n309), .o1(new_n311));
  oao003aa1n03x5               g216(.a(\a[28] ), .b(\b[27] ), .c(new_n303), .carry(new_n312));
  aoai13aa1n02x7               g217(.a(new_n312), .b(new_n311), .c(new_n301), .d(new_n293), .o1(new_n313));
  xorc02aa1n12x5               g218(.a(\a[29] ), .b(\b[28] ), .out0(new_n314));
  norb02aa1n02x5               g219(.a(new_n312), .b(new_n314), .out0(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n310), .d(new_n315), .o1(\s[29] ));
  xorb03aa1n02x5               g221(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g222(.a(new_n304), .b(new_n306), .c(new_n314), .out0(new_n318));
  aoai13aa1n02x5               g223(.a(new_n318), .b(new_n296), .c(new_n196), .d(new_n292), .o1(new_n319));
  inv000aa1n02x5               g224(.a(new_n318), .o1(new_n320));
  tech160nm_fioaoi03aa1n03p5x5 g225(.a(\a[29] ), .b(\b[28] ), .c(new_n312), .o1(new_n321));
  inv000aa1d42x5               g226(.a(new_n321), .o1(new_n322));
  aoai13aa1n02x7               g227(.a(new_n322), .b(new_n320), .c(new_n301), .d(new_n293), .o1(new_n323));
  tech160nm_fixorc02aa1n03p5x5 g228(.a(\a[30] ), .b(\b[29] ), .out0(new_n324));
  and002aa1n02x5               g229(.a(\b[28] ), .b(\a[29] ), .o(new_n325));
  oabi12aa1n02x5               g230(.a(new_n324), .b(\a[29] ), .c(\b[28] ), .out0(new_n326));
  oab012aa1n02x4               g231(.a(new_n326), .b(new_n312), .c(new_n325), .out0(new_n327));
  aoi022aa1n03x5               g232(.a(new_n323), .b(new_n324), .c(new_n319), .d(new_n327), .o1(\s[30] ));
  nano32aa1n02x4               g233(.a(new_n304), .b(new_n324), .c(new_n306), .d(new_n314), .out0(new_n329));
  aoai13aa1n02x5               g234(.a(new_n329), .b(new_n296), .c(new_n196), .d(new_n292), .o1(new_n330));
  inv000aa1n02x5               g235(.a(new_n329), .o1(new_n331));
  inv000aa1d42x5               g236(.a(\a[30] ), .o1(new_n332));
  inv000aa1d42x5               g237(.a(\b[29] ), .o1(new_n333));
  oaoi03aa1n03x5               g238(.a(new_n332), .b(new_n333), .c(new_n321), .o1(new_n334));
  aoai13aa1n03x5               g239(.a(new_n334), .b(new_n331), .c(new_n301), .d(new_n293), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  oabi12aa1n02x5               g241(.a(new_n336), .b(\a[30] ), .c(\b[29] ), .out0(new_n337));
  oaoi13aa1n02x5               g242(.a(new_n337), .b(new_n321), .c(new_n332), .d(new_n333), .o1(new_n338));
  aoi022aa1n03x5               g243(.a(new_n335), .b(new_n336), .c(new_n330), .d(new_n338), .o1(\s[31] ));
  norb02aa1n02x5               g244(.a(new_n105), .b(new_n107), .out0(new_n340));
  xobna2aa1n03x5               g245(.a(new_n340), .b(new_n103), .c(new_n100), .out0(\s[3] ));
  aoai13aa1n02x5               g246(.a(new_n340), .b(new_n102), .c(\a[2] ), .d(\b[1] ), .o1(new_n342));
  nanb02aa1n02x5               g247(.a(new_n110), .b(new_n106), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n342), .c(new_n105), .out0(\s[4] ));
  inv000aa1d42x5               g249(.a(new_n117), .o1(new_n345));
  xnbna2aa1n03x5               g250(.a(new_n345), .b(new_n109), .c(new_n111), .out0(\s[5] ));
  nanp02aa1n02x5               g251(.a(new_n125), .b(new_n124), .o1(new_n347));
  nanp02aa1n03x5               g252(.a(new_n133), .b(new_n345), .o1(new_n348));
  xnbna2aa1n03x5               g253(.a(new_n114), .b(new_n348), .c(new_n347), .out0(\s[6] ));
  inv000aa1d42x5               g254(.a(new_n113), .o1(new_n350));
  aob012aa1n02x5               g255(.a(new_n114), .b(new_n348), .c(new_n347), .out0(new_n351));
  xnbna2aa1n03x5               g256(.a(new_n116), .b(new_n351), .c(new_n350), .out0(\s[7] ));
  aob012aa1n03x5               g257(.a(new_n116), .b(new_n351), .c(new_n350), .out0(new_n353));
  nanp02aa1n02x5               g258(.a(new_n353), .b(new_n123), .o1(new_n354));
  norb02aa1n02x5               g259(.a(new_n123), .b(new_n134), .out0(new_n355));
  aoi022aa1n02x5               g260(.a(new_n354), .b(new_n134), .c(new_n353), .d(new_n355), .o1(\s[8] ));
  aoi112aa1n02x5               g261(.a(new_n128), .b(new_n131), .c(new_n119), .d(new_n120), .o1(new_n357));
  aoi022aa1n02x5               g262(.a(new_n130), .b(new_n131), .c(new_n155), .d(new_n357), .o1(\s[9] ));
endmodule


