// Benchmark "adder" written by ABC on Thu Jul 18 04:57:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n312, new_n315, new_n317, new_n319;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[8] ), .o1(new_n97));
  xnrc02aa1n12x5               g002(.a(\b[5] ), .b(\a[6] ), .out0(new_n98));
  orn002aa1n24x5               g003(.a(\a[5] ), .b(\b[4] ), .o(new_n99));
  nanp02aa1n02x5               g004(.a(\b[4] ), .b(\a[5] ), .o1(new_n100));
  nand02aa1n03x5               g005(.a(new_n99), .b(new_n100), .o1(new_n101));
  nor002aa1n03x5               g006(.a(new_n98), .b(new_n101), .o1(new_n102));
  nanp02aa1n04x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  nand02aa1n06x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  nor022aa1n16x5               g010(.a(\b[6] ), .b(\a[7] ), .o1(new_n106));
  nona23aa1d18x5               g011(.a(new_n105), .b(new_n103), .c(new_n106), .d(new_n104), .out0(new_n107));
  and002aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o(new_n108));
  oa0022aa1n09x5               g013(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n109));
  inv040aa1d32x5               g014(.a(\a[3] ), .o1(new_n110));
  inv040aa1d32x5               g015(.a(\b[2] ), .o1(new_n111));
  nand42aa1n04x5               g016(.a(new_n111), .b(new_n110), .o1(new_n112));
  nanp02aa1n04x5               g017(.a(\b[2] ), .b(\a[3] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(new_n112), .b(new_n113), .o1(new_n114));
  nor042aa1n03x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nand42aa1n10x5               g020(.a(\b[1] ), .b(\a[2] ), .o1(new_n116));
  nand42aa1d28x5               g021(.a(\b[0] ), .b(\a[1] ), .o1(new_n117));
  aoi012aa1n09x5               g022(.a(new_n115), .b(new_n116), .c(new_n117), .o1(new_n118));
  oaih12aa1n02x5               g023(.a(new_n109), .b(new_n118), .c(new_n114), .o1(new_n119));
  nona23aa1n06x5               g024(.a(new_n119), .b(new_n102), .c(new_n107), .d(new_n108), .out0(new_n120));
  nona22aa1n02x4               g025(.a(new_n105), .b(new_n106), .c(new_n104), .out0(new_n121));
  oaoi03aa1n09x5               g026(.a(\a[6] ), .b(\b[5] ), .c(new_n99), .o1(new_n122));
  aboi22aa1n03x5               g027(.a(new_n107), .b(new_n122), .c(new_n105), .d(new_n121), .out0(new_n123));
  nanp02aa1n06x5               g028(.a(new_n120), .b(new_n123), .o1(new_n124));
  oaib12aa1n06x5               g029(.a(new_n124), .b(new_n97), .c(\a[9] ), .out0(new_n125));
  oa0012aa1n02x5               g030(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .o(new_n126));
  xnrb03aa1n02x5               g031(.a(new_n126), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nand02aa1d16x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nand02aa1d28x5               g033(.a(\b[10] ), .b(\a[11] ), .o1(new_n129));
  nor042aa1n06x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n129), .b(new_n130), .out0(new_n131));
  oai122aa1n06x5               g036(.a(new_n125), .b(\b[9] ), .c(\a[10] ), .d(\b[8] ), .e(\a[9] ), .o1(new_n132));
  xobna2aa1n03x5               g037(.a(new_n131), .b(new_n132), .c(new_n128), .out0(\s[11] ));
  inv040aa1n02x5               g038(.a(new_n130), .o1(new_n134));
  nanp03aa1n03x5               g039(.a(new_n132), .b(new_n128), .c(new_n131), .o1(new_n135));
  xnrc02aa1n12x5               g040(.a(\b[11] ), .b(\a[12] ), .out0(new_n136));
  tech160nm_fiaoi012aa1n02p5x5 g041(.a(new_n136), .b(new_n135), .c(new_n134), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n136), .o1(new_n138));
  aoi113aa1n03x5               g043(.a(new_n130), .b(new_n138), .c(new_n132), .d(new_n128), .e(new_n129), .o1(new_n139));
  nor002aa1n02x5               g044(.a(new_n137), .b(new_n139), .o1(\s[12] ));
  tech160nm_fixnrc02aa1n04x5   g045(.a(\b[8] ), .b(\a[9] ), .out0(new_n141));
  norp02aa1n02x5               g046(.a(\b[9] ), .b(\a[10] ), .o1(new_n142));
  nano23aa1n03x7               g047(.a(new_n130), .b(new_n142), .c(new_n128), .d(new_n129), .out0(new_n143));
  nona22aa1n09x5               g048(.a(new_n143), .b(new_n141), .c(new_n136), .out0(new_n144));
  inv000aa1n02x5               g049(.a(new_n144), .o1(new_n145));
  inv000aa1d42x5               g050(.a(\b[11] ), .o1(new_n146));
  nanb02aa1d24x5               g051(.a(\a[12] ), .b(new_n146), .out0(new_n147));
  and002aa1n02x5               g052(.a(\b[11] ), .b(\a[12] ), .o(new_n148));
  oai022aa1d18x5               g053(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n149));
  nand23aa1d12x5               g054(.a(new_n149), .b(new_n128), .c(new_n129), .o1(new_n150));
  aoi013aa1n09x5               g055(.a(new_n148), .b(new_n150), .c(new_n134), .d(new_n147), .o1(new_n151));
  aoi012aa1n02x5               g056(.a(new_n151), .b(new_n124), .c(new_n145), .o1(new_n152));
  xnrb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  oaoi03aa1n03x5               g058(.a(\a[13] ), .b(\b[12] ), .c(new_n152), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp03aa1n06x5               g060(.a(new_n107), .b(new_n101), .c(new_n98), .o1(new_n156));
  oaoi13aa1n09x5               g061(.a(new_n108), .b(new_n109), .c(new_n118), .d(new_n114), .o1(new_n157));
  inv000aa1d42x5               g062(.a(\a[7] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(\b[6] ), .o1(new_n159));
  aoai13aa1n02x5               g064(.a(new_n105), .b(new_n104), .c(new_n158), .d(new_n159), .o1(new_n160));
  oaib12aa1n06x5               g065(.a(new_n160), .b(new_n107), .c(new_n122), .out0(new_n161));
  aoai13aa1n03x5               g066(.a(new_n145), .b(new_n161), .c(new_n157), .d(new_n156), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n151), .o1(new_n163));
  nor042aa1d18x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nor042aa1d18x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nand42aa1n16x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nona23aa1n02x4               g072(.a(new_n167), .b(new_n165), .c(new_n164), .d(new_n166), .out0(new_n168));
  oai012aa1n02x5               g073(.a(new_n167), .b(new_n166), .c(new_n164), .o1(new_n169));
  aoai13aa1n02x7               g074(.a(new_n169), .b(new_n168), .c(new_n162), .d(new_n163), .o1(new_n170));
  xorb03aa1n02x5               g075(.a(new_n170), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  tech160nm_fixorc02aa1n02p5x5 g077(.a(\a[15] ), .b(\b[14] ), .out0(new_n173));
  tech160nm_fixorc02aa1n02p5x5 g078(.a(\a[16] ), .b(\b[15] ), .out0(new_n174));
  aoi112aa1n02x5               g079(.a(new_n172), .b(new_n174), .c(new_n170), .d(new_n173), .o1(new_n175));
  aoai13aa1n03x5               g080(.a(new_n174), .b(new_n172), .c(new_n170), .d(new_n173), .o1(new_n176));
  norb02aa1n02x7               g081(.a(new_n176), .b(new_n175), .out0(\s[16] ));
  nano23aa1n03x7               g082(.a(new_n164), .b(new_n166), .c(new_n167), .d(new_n165), .out0(new_n178));
  nand23aa1n03x5               g083(.a(new_n178), .b(new_n173), .c(new_n174), .o1(new_n179));
  nor042aa1n06x5               g084(.a(new_n144), .b(new_n179), .o1(new_n180));
  aoai13aa1n12x5               g085(.a(new_n180), .b(new_n161), .c(new_n157), .d(new_n156), .o1(new_n181));
  tech160nm_fixnrc02aa1n02p5x5 g086(.a(\b[14] ), .b(\a[15] ), .out0(new_n182));
  xnrc02aa1n03x5               g087(.a(\b[15] ), .b(\a[16] ), .out0(new_n183));
  nor043aa1n02x5               g088(.a(new_n168), .b(new_n182), .c(new_n183), .o1(new_n184));
  aoi112aa1n03x4               g089(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n185));
  nor002aa1n03x5               g090(.a(\b[15] ), .b(\a[16] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(new_n186), .o1(new_n187));
  oai013aa1n02x5               g092(.a(new_n187), .b(new_n182), .c(new_n183), .d(new_n169), .o1(new_n188));
  aoi112aa1n09x5               g093(.a(new_n188), .b(new_n185), .c(new_n151), .d(new_n184), .o1(new_n189));
  nand02aa1d08x5               g094(.a(new_n181), .b(new_n189), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[18] ), .o1(new_n192));
  inv040aa1d32x5               g097(.a(\a[17] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[16] ), .o1(new_n194));
  oaoi03aa1n03x5               g099(.a(new_n193), .b(new_n194), .c(new_n190), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(new_n192), .out0(\s[18] ));
  xroi22aa1d06x4               g101(.a(new_n193), .b(\b[16] ), .c(new_n192), .d(\b[17] ), .out0(new_n197));
  nanp02aa1n02x5               g102(.a(new_n194), .b(new_n193), .o1(new_n198));
  oaoi03aa1n12x5               g103(.a(\a[18] ), .b(\b[17] ), .c(new_n198), .o1(new_n199));
  nor022aa1n16x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand02aa1d06x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  norb02aa1n02x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  aoai13aa1n06x5               g107(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n197), .o1(new_n203));
  aoi112aa1n02x5               g108(.a(new_n202), .b(new_n199), .c(new_n190), .d(new_n197), .o1(new_n204));
  norb02aa1n03x4               g109(.a(new_n203), .b(new_n204), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nand02aa1d06x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  nona22aa1n02x5               g114(.a(new_n203), .b(new_n209), .c(new_n200), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n209), .o1(new_n211));
  oaoi13aa1n06x5               g116(.a(new_n211), .b(new_n203), .c(\a[19] ), .d(\b[18] ), .o1(new_n212));
  norb02aa1n03x4               g117(.a(new_n210), .b(new_n212), .out0(\s[20] ));
  nano23aa1n03x7               g118(.a(new_n200), .b(new_n207), .c(new_n208), .d(new_n201), .out0(new_n214));
  nanp02aa1n02x5               g119(.a(new_n197), .b(new_n214), .o1(new_n215));
  oai022aa1n02x7               g120(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n216));
  oaib12aa1n09x5               g121(.a(new_n216), .b(new_n192), .c(\b[17] ), .out0(new_n217));
  nona23aa1n09x5               g122(.a(new_n208), .b(new_n201), .c(new_n200), .d(new_n207), .out0(new_n218));
  aoi012aa1n06x5               g123(.a(new_n207), .b(new_n200), .c(new_n208), .o1(new_n219));
  oai012aa1n18x5               g124(.a(new_n219), .b(new_n218), .c(new_n217), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  aoai13aa1n06x5               g126(.a(new_n221), .b(new_n215), .c(new_n181), .d(new_n189), .o1(new_n222));
  xorb03aa1n02x5               g127(.a(new_n222), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  xorc02aa1n02x5               g129(.a(\a[21] ), .b(\b[20] ), .out0(new_n225));
  xorc02aa1n02x5               g130(.a(\a[22] ), .b(\b[21] ), .out0(new_n226));
  aoi112aa1n02x7               g131(.a(new_n224), .b(new_n226), .c(new_n222), .d(new_n225), .o1(new_n227));
  aoai13aa1n03x5               g132(.a(new_n226), .b(new_n224), .c(new_n222), .d(new_n225), .o1(new_n228));
  norb02aa1n02x7               g133(.a(new_n228), .b(new_n227), .out0(\s[22] ));
  inv000aa1d42x5               g134(.a(\a[21] ), .o1(new_n230));
  inv000aa1d42x5               g135(.a(\a[22] ), .o1(new_n231));
  xroi22aa1d06x4               g136(.a(new_n230), .b(\b[20] ), .c(new_n231), .d(\b[21] ), .out0(new_n232));
  nanp03aa1n02x5               g137(.a(new_n232), .b(new_n197), .c(new_n214), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\b[21] ), .o1(new_n234));
  oaoi03aa1n12x5               g139(.a(new_n231), .b(new_n234), .c(new_n224), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n220), .c(new_n232), .o1(new_n237));
  aoai13aa1n06x5               g142(.a(new_n237), .b(new_n233), .c(new_n181), .d(new_n189), .o1(new_n238));
  xorb03aa1n03x5               g143(.a(new_n238), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g144(.a(\b[22] ), .b(\a[23] ), .o1(new_n240));
  tech160nm_fixorc02aa1n05x5   g145(.a(\a[23] ), .b(\b[22] ), .out0(new_n241));
  xorc02aa1n03x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  aoi112aa1n02x5               g147(.a(new_n240), .b(new_n242), .c(new_n238), .d(new_n241), .o1(new_n243));
  aoai13aa1n03x5               g148(.a(new_n242), .b(new_n240), .c(new_n238), .d(new_n241), .o1(new_n244));
  norb02aa1n03x4               g149(.a(new_n244), .b(new_n243), .out0(\s[24] ));
  and002aa1n02x5               g150(.a(new_n242), .b(new_n241), .o(new_n246));
  inv000aa1n02x5               g151(.a(new_n246), .o1(new_n247));
  nano32aa1n02x4               g152(.a(new_n247), .b(new_n232), .c(new_n197), .d(new_n214), .out0(new_n248));
  inv000aa1n02x5               g153(.a(new_n219), .o1(new_n249));
  aoai13aa1n03x5               g154(.a(new_n232), .b(new_n249), .c(new_n214), .d(new_n199), .o1(new_n250));
  norp02aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nanp02aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  aoi012aa1n02x5               g157(.a(new_n251), .b(new_n240), .c(new_n252), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n247), .c(new_n250), .d(new_n235), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[25] ), .b(\b[24] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n190), .d(new_n248), .o1(new_n256));
  aoi112aa1n02x5               g161(.a(new_n255), .b(new_n254), .c(new_n190), .d(new_n248), .o1(new_n257));
  norb02aa1n03x4               g162(.a(new_n256), .b(new_n257), .out0(\s[25] ));
  norp02aa1n02x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  tech160nm_fixorc02aa1n05x5   g164(.a(\a[26] ), .b(\b[25] ), .out0(new_n260));
  nona22aa1n02x5               g165(.a(new_n256), .b(new_n260), .c(new_n259), .out0(new_n261));
  inv000aa1n02x5               g166(.a(new_n259), .o1(new_n262));
  aobi12aa1n06x5               g167(.a(new_n260), .b(new_n256), .c(new_n262), .out0(new_n263));
  norb02aa1n03x4               g168(.a(new_n261), .b(new_n263), .out0(\s[26] ));
  nanp02aa1n02x5               g169(.a(new_n151), .b(new_n184), .o1(new_n265));
  nona22aa1n02x4               g170(.a(new_n265), .b(new_n188), .c(new_n185), .out0(new_n266));
  and002aa1n06x5               g171(.a(new_n260), .b(new_n255), .o(new_n267));
  nano22aa1n03x7               g172(.a(new_n233), .b(new_n246), .c(new_n267), .out0(new_n268));
  aoai13aa1n06x5               g173(.a(new_n268), .b(new_n266), .c(new_n124), .d(new_n180), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .c(new_n262), .carry(new_n270));
  aobi12aa1n06x5               g175(.a(new_n270), .b(new_n254), .c(new_n267), .out0(new_n271));
  xorc02aa1n12x5               g176(.a(\a[27] ), .b(\b[26] ), .out0(new_n272));
  xnbna2aa1n03x5               g177(.a(new_n272), .b(new_n271), .c(new_n269), .out0(\s[27] ));
  norp02aa1n02x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  inv040aa1n03x5               g179(.a(new_n274), .o1(new_n275));
  aobi12aa1n02x7               g180(.a(new_n272), .b(new_n271), .c(new_n269), .out0(new_n276));
  xnrc02aa1n02x5               g181(.a(\b[27] ), .b(\a[28] ), .out0(new_n277));
  nano22aa1n02x4               g182(.a(new_n276), .b(new_n275), .c(new_n277), .out0(new_n278));
  aobi12aa1n06x5               g183(.a(new_n268), .b(new_n181), .c(new_n189), .out0(new_n279));
  aoai13aa1n02x5               g184(.a(new_n246), .b(new_n236), .c(new_n220), .d(new_n232), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n267), .o1(new_n281));
  aoai13aa1n06x5               g186(.a(new_n270), .b(new_n281), .c(new_n280), .d(new_n253), .o1(new_n282));
  oaih12aa1n02x5               g187(.a(new_n272), .b(new_n282), .c(new_n279), .o1(new_n283));
  aoi012aa1n03x5               g188(.a(new_n277), .b(new_n283), .c(new_n275), .o1(new_n284));
  norp02aa1n03x5               g189(.a(new_n284), .b(new_n278), .o1(\s[28] ));
  xnrc02aa1n02x5               g190(.a(\b[28] ), .b(\a[29] ), .out0(new_n286));
  norb02aa1n02x5               g191(.a(new_n272), .b(new_n277), .out0(new_n287));
  aobi12aa1n03x5               g192(.a(new_n287), .b(new_n271), .c(new_n269), .out0(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n275), .carry(new_n289));
  nano22aa1n02x4               g194(.a(new_n288), .b(new_n286), .c(new_n289), .out0(new_n290));
  oaih12aa1n02x5               g195(.a(new_n287), .b(new_n282), .c(new_n279), .o1(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n286), .b(new_n291), .c(new_n289), .o1(new_n292));
  nor002aa1n02x5               g197(.a(new_n292), .b(new_n290), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n117), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g199(.a(new_n272), .b(new_n286), .c(new_n277), .out0(new_n295));
  aobi12aa1n02x7               g200(.a(new_n295), .b(new_n271), .c(new_n269), .out0(new_n296));
  oao003aa1n02x5               g201(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n297));
  xnrc02aa1n02x5               g202(.a(\b[29] ), .b(\a[30] ), .out0(new_n298));
  nano22aa1n02x4               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  oaih12aa1n02x5               g204(.a(new_n295), .b(new_n282), .c(new_n279), .o1(new_n300));
  tech160nm_fiaoi012aa1n02p5x5 g205(.a(new_n298), .b(new_n300), .c(new_n297), .o1(new_n301));
  nor002aa1n02x5               g206(.a(new_n301), .b(new_n299), .o1(\s[30] ));
  norb02aa1n02x5               g207(.a(new_n295), .b(new_n298), .out0(new_n303));
  aobi12aa1n02x7               g208(.a(new_n303), .b(new_n271), .c(new_n269), .out0(new_n304));
  oao003aa1n02x5               g209(.a(\a[30] ), .b(\b[29] ), .c(new_n297), .carry(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[30] ), .b(\a[31] ), .out0(new_n306));
  nano22aa1n02x4               g211(.a(new_n304), .b(new_n305), .c(new_n306), .out0(new_n307));
  oaih12aa1n02x5               g212(.a(new_n303), .b(new_n282), .c(new_n279), .o1(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n306), .b(new_n308), .c(new_n305), .o1(new_n309));
  norp02aa1n03x5               g214(.a(new_n309), .b(new_n307), .o1(\s[31] ));
  xnbna2aa1n03x5               g215(.a(new_n118), .b(new_n112), .c(new_n113), .out0(\s[3] ));
  oaoi03aa1n02x5               g216(.a(\a[3] ), .b(\b[2] ), .c(new_n118), .o1(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g218(.a(new_n157), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nona22aa1n02x4               g219(.a(new_n119), .b(new_n108), .c(new_n101), .out0(new_n315));
  xobna2aa1n03x5               g220(.a(new_n98), .b(new_n315), .c(new_n99), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g221(.a(new_n122), .b(new_n157), .c(new_n102), .o(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g223(.a(new_n158), .b(new_n159), .c(new_n317), .o1(new_n319));
  xnrb03aa1n02x5               g224(.a(new_n319), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xobna2aa1n03x5               g225(.a(new_n141), .b(new_n120), .c(new_n123), .out0(\s[9] ));
endmodule


