// Benchmark "adder" written by ABC on Thu Jul 11 12:32:43 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n147, new_n148, new_n149,
    new_n150, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n175, new_n176, new_n177, new_n178, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n308, new_n311, new_n312,
    new_n313, new_n315, new_n317;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  160nm_ficinv00aa1n08x5       g001(.clk(\a[2] ), .clkout(new_n97));
  160nm_ficinv00aa1n08x5       g002(.clk(\b[1] ), .clkout(new_n98));
  nanp02aa1n02x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  oaoi03aa1n02x5               g004(.a(new_n97), .b(new_n98), .c(new_n99), .o1(new_n100));
  norp02aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  nanp02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nona23aa1n02x4               g009(.a(new_n104), .b(new_n102), .c(new_n101), .d(new_n103), .out0(new_n105));
  aoi012aa1n02x5               g010(.a(new_n101), .b(new_n103), .c(new_n102), .o1(new_n106));
  oai012aa1n02x5               g011(.a(new_n106), .b(new_n105), .c(new_n100), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[7] ), .b(\a[8] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  norp02aa1n02x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nona23aa1n02x4               g016(.a(new_n111), .b(new_n109), .c(new_n108), .d(new_n110), .out0(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[5] ), .b(\a[6] ), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  norp03aa1n02x5               g019(.a(new_n112), .b(new_n113), .c(new_n114), .o1(new_n115));
  orn002aa1n02x5               g020(.a(\a[5] ), .b(\b[4] ), .o(new_n116));
  oaoi03aa1n02x5               g021(.a(\a[6] ), .b(\b[5] ), .c(new_n116), .o1(new_n117));
  aoi012aa1n02x5               g022(.a(new_n108), .b(new_n110), .c(new_n109), .o1(new_n118));
  oaib12aa1n02x5               g023(.a(new_n118), .b(new_n112), .c(new_n117), .out0(new_n119));
  aoi012aa1n02x5               g024(.a(new_n119), .b(new_n107), .c(new_n115), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[9] ), .b(\b[8] ), .c(new_n120), .o1(new_n121));
  xorb03aa1n02x5               g026(.a(new_n121), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  norp02aa1n02x5               g027(.a(\b[10] ), .b(\a[11] ), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  norb02aa1n02x5               g029(.a(new_n124), .b(new_n123), .out0(new_n125));
  norp02aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norp02aa1n02x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  oai012aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n126), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nano23aa1n02x4               g035(.a(new_n126), .b(new_n127), .c(new_n128), .d(new_n130), .out0(new_n131));
  aoai13aa1n02x5               g036(.a(new_n131), .b(new_n119), .c(new_n107), .d(new_n115), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n125), .b(new_n132), .c(new_n129), .out0(\s[11] ));
  160nm_ficinv00aa1n08x5       g038(.clk(new_n131), .clkout(new_n134));
  oai012aa1n02x5               g039(.a(new_n129), .b(new_n120), .c(new_n134), .o1(new_n135));
  aoi012aa1n02x5               g040(.a(new_n123), .b(new_n135), .c(new_n124), .o1(new_n136));
  xnrb03aa1n02x5               g041(.a(new_n136), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  norp02aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nano23aa1n02x4               g044(.a(new_n123), .b(new_n138), .c(new_n139), .d(new_n124), .out0(new_n140));
  nanp02aa1n02x5               g045(.a(new_n140), .b(new_n131), .o1(new_n141));
  nona23aa1n02x4               g046(.a(new_n139), .b(new_n124), .c(new_n123), .d(new_n138), .out0(new_n142));
  160nm_fiao0012aa1n02p5x5     g047(.a(new_n138), .b(new_n123), .c(new_n139), .o(new_n143));
  oabi12aa1n02x5               g048(.a(new_n143), .b(new_n142), .c(new_n129), .out0(new_n144));
  oabi12aa1n02x5               g049(.a(new_n144), .b(new_n120), .c(new_n141), .out0(new_n145));
  xorb03aa1n02x5               g050(.a(new_n145), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  orn002aa1n02x5               g051(.a(\a[13] ), .b(\b[12] ), .o(new_n147));
  xnrc02aa1n02x5               g052(.a(\b[12] ), .b(\a[13] ), .out0(new_n148));
  nanb02aa1n02x5               g053(.a(new_n148), .b(new_n145), .out0(new_n149));
  xnrc02aa1n02x5               g054(.a(\b[13] ), .b(\a[14] ), .out0(new_n150));
  xobna2aa1n03x5               g055(.a(new_n150), .b(new_n149), .c(new_n147), .out0(\s[14] ));
  norp02aa1n02x5               g056(.a(\b[14] ), .b(\a[15] ), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(\b[14] ), .b(\a[15] ), .o1(new_n153));
  nanb02aa1n02x5               g058(.a(new_n152), .b(new_n153), .out0(new_n154));
  160nm_ficinv00aa1n08x5       g059(.clk(new_n154), .clkout(new_n155));
  norp02aa1n02x5               g060(.a(new_n150), .b(new_n148), .o1(new_n156));
  oaoi03aa1n02x5               g061(.a(\a[14] ), .b(\b[13] ), .c(new_n147), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n155), .b(new_n157), .c(new_n145), .d(new_n156), .o1(new_n158));
  aoi112aa1n02x5               g063(.a(new_n155), .b(new_n157), .c(new_n145), .d(new_n156), .o1(new_n159));
  norb02aa1n02x5               g064(.a(new_n158), .b(new_n159), .out0(\s[15] ));
  160nm_ficinv00aa1n08x5       g065(.clk(new_n152), .clkout(new_n161));
  norp02aa1n02x5               g066(.a(\b[15] ), .b(\a[16] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[15] ), .b(\a[16] ), .o1(new_n163));
  nanb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  nanp03aa1n02x5               g069(.a(new_n158), .b(new_n161), .c(new_n164), .o1(new_n165));
  aoi012aa1n02x5               g070(.a(new_n164), .b(new_n158), .c(new_n161), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n165), .b(new_n166), .out0(\s[16] ));
  nano23aa1n02x4               g072(.a(new_n152), .b(new_n162), .c(new_n163), .d(new_n153), .out0(new_n168));
  nano22aa1n02x4               g073(.a(new_n141), .b(new_n156), .c(new_n168), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n119), .c(new_n107), .d(new_n115), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n168), .b(new_n157), .c(new_n144), .d(new_n156), .o1(new_n171));
  aoi012aa1n02x5               g076(.a(new_n162), .b(new_n152), .c(new_n163), .o1(new_n172));
  nanp03aa1n02x5               g077(.a(new_n170), .b(new_n171), .c(new_n172), .o1(new_n173));
  xorb03aa1n02x5               g078(.a(new_n173), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g079(.clk(\a[18] ), .clkout(new_n175));
  160nm_ficinv00aa1n08x5       g080(.clk(\a[17] ), .clkout(new_n176));
  160nm_ficinv00aa1n08x5       g081(.clk(\b[16] ), .clkout(new_n177));
  oaoi03aa1n02x5               g082(.a(new_n176), .b(new_n177), .c(new_n173), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[17] ), .c(new_n175), .out0(\s[18] ));
  160nm_ficinv00aa1n08x5       g084(.clk(new_n120), .clkout(new_n180));
  160nm_ficinv00aa1n08x5       g085(.clk(new_n157), .clkout(new_n181));
  160nm_ficinv00aa1n08x5       g086(.clk(new_n168), .clkout(new_n182));
  160nm_ficinv00aa1n08x5       g087(.clk(new_n129), .clkout(new_n183));
  aoai13aa1n02x5               g088(.a(new_n156), .b(new_n143), .c(new_n140), .d(new_n183), .o1(new_n184));
  aoai13aa1n02x5               g089(.a(new_n172), .b(new_n182), .c(new_n184), .d(new_n181), .o1(new_n185));
  xroi22aa1d04x5               g090(.a(new_n176), .b(\b[16] ), .c(new_n175), .d(\b[17] ), .out0(new_n186));
  aoai13aa1n02x5               g091(.a(new_n186), .b(new_n185), .c(new_n180), .d(new_n169), .o1(new_n187));
  oai022aa1n02x5               g092(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n188));
  oaib12aa1n02x5               g093(.a(new_n188), .b(new_n175), .c(\b[17] ), .out0(new_n189));
  norp02aa1n02x5               g094(.a(\b[18] ), .b(\a[19] ), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nanb02aa1n02x5               g096(.a(new_n190), .b(new_n191), .out0(new_n192));
  160nm_ficinv00aa1n08x5       g097(.clk(new_n192), .clkout(new_n193));
  xnbna2aa1n03x5               g098(.a(new_n193), .b(new_n187), .c(new_n189), .out0(\s[19] ));
  xnrc02aa1n02x5               g099(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  160nm_ficinv00aa1n08x5       g100(.clk(new_n190), .clkout(new_n196));
  aoi012aa1n02x5               g101(.a(new_n192), .b(new_n187), .c(new_n189), .o1(new_n197));
  norp02aa1n02x5               g102(.a(\b[19] ), .b(\a[20] ), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  nano22aa1n02x4               g105(.a(new_n197), .b(new_n196), .c(new_n200), .out0(new_n201));
  nanp02aa1n02x5               g106(.a(new_n177), .b(new_n176), .o1(new_n202));
  oaoi03aa1n02x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n202), .o1(new_n203));
  aoai13aa1n02x5               g108(.a(new_n193), .b(new_n203), .c(new_n173), .d(new_n186), .o1(new_n204));
  aoi012aa1n02x5               g109(.a(new_n200), .b(new_n204), .c(new_n196), .o1(new_n205));
  norp02aa1n02x5               g110(.a(new_n205), .b(new_n201), .o1(\s[20] ));
  nano23aa1n02x4               g111(.a(new_n190), .b(new_n198), .c(new_n199), .d(new_n191), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(new_n186), .b(new_n207), .o1(new_n208));
  160nm_ficinv00aa1n08x5       g113(.clk(new_n208), .clkout(new_n209));
  aoai13aa1n02x5               g114(.a(new_n209), .b(new_n185), .c(new_n180), .d(new_n169), .o1(new_n210));
  nona23aa1n02x4               g115(.a(new_n199), .b(new_n191), .c(new_n190), .d(new_n198), .out0(new_n211));
  aoi012aa1n02x5               g116(.a(new_n198), .b(new_n190), .c(new_n199), .o1(new_n212));
  oai012aa1n02x5               g117(.a(new_n212), .b(new_n211), .c(new_n189), .o1(new_n213));
  160nm_ficinv00aa1n08x5       g118(.clk(new_n213), .clkout(new_n214));
  norp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  nanp02aa1n02x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  norb02aa1n02x5               g121(.a(new_n216), .b(new_n215), .out0(new_n217));
  xnbna2aa1n03x5               g122(.a(new_n217), .b(new_n210), .c(new_n214), .out0(\s[21] ));
  160nm_ficinv00aa1n08x5       g123(.clk(new_n215), .clkout(new_n219));
  aobi12aa1n02x5               g124(.a(new_n217), .b(new_n210), .c(new_n214), .out0(new_n220));
  xnrc02aa1n02x5               g125(.a(\b[21] ), .b(\a[22] ), .out0(new_n221));
  nano22aa1n02x4               g126(.a(new_n220), .b(new_n219), .c(new_n221), .out0(new_n222));
  aoai13aa1n02x5               g127(.a(new_n217), .b(new_n213), .c(new_n173), .d(new_n209), .o1(new_n223));
  aoi012aa1n02x5               g128(.a(new_n221), .b(new_n223), .c(new_n219), .o1(new_n224));
  norp02aa1n02x5               g129(.a(new_n224), .b(new_n222), .o1(\s[22] ));
  nano22aa1n02x4               g130(.a(new_n221), .b(new_n219), .c(new_n216), .out0(new_n226));
  and003aa1n02x5               g131(.a(new_n186), .b(new_n226), .c(new_n207), .o(new_n227));
  aoai13aa1n02x5               g132(.a(new_n227), .b(new_n185), .c(new_n180), .d(new_n169), .o1(new_n228));
  oao003aa1n02x5               g133(.a(\a[22] ), .b(\b[21] ), .c(new_n219), .carry(new_n229));
  160nm_ficinv00aa1n08x5       g134(.clk(new_n229), .clkout(new_n230));
  aoi012aa1n02x5               g135(.a(new_n230), .b(new_n213), .c(new_n226), .o1(new_n231));
  xnrc02aa1n02x5               g136(.a(\b[22] ), .b(\a[23] ), .out0(new_n232));
  160nm_ficinv00aa1n08x5       g137(.clk(new_n232), .clkout(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n228), .c(new_n231), .out0(\s[23] ));
  norp02aa1n02x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  160nm_ficinv00aa1n08x5       g140(.clk(new_n235), .clkout(new_n236));
  aoi012aa1n02x5               g141(.a(new_n232), .b(new_n228), .c(new_n231), .o1(new_n237));
  xnrc02aa1n02x5               g142(.a(\b[23] ), .b(\a[24] ), .out0(new_n238));
  nano22aa1n02x4               g143(.a(new_n237), .b(new_n236), .c(new_n238), .out0(new_n239));
  160nm_ficinv00aa1n08x5       g144(.clk(new_n231), .clkout(new_n240));
  aoai13aa1n02x5               g145(.a(new_n233), .b(new_n240), .c(new_n173), .d(new_n227), .o1(new_n241));
  aoi012aa1n02x5               g146(.a(new_n238), .b(new_n241), .c(new_n236), .o1(new_n242));
  norp02aa1n02x5               g147(.a(new_n242), .b(new_n239), .o1(\s[24] ));
  norp02aa1n02x5               g148(.a(new_n238), .b(new_n232), .o1(new_n244));
  nano22aa1n02x4               g149(.a(new_n208), .b(new_n226), .c(new_n244), .out0(new_n245));
  aoai13aa1n02x5               g150(.a(new_n245), .b(new_n185), .c(new_n180), .d(new_n169), .o1(new_n246));
  160nm_ficinv00aa1n08x5       g151(.clk(new_n212), .clkout(new_n247));
  aoai13aa1n02x5               g152(.a(new_n226), .b(new_n247), .c(new_n207), .d(new_n203), .o1(new_n248));
  160nm_ficinv00aa1n08x5       g153(.clk(new_n244), .clkout(new_n249));
  oao003aa1n02x5               g154(.a(\a[24] ), .b(\b[23] ), .c(new_n236), .carry(new_n250));
  aoai13aa1n02x5               g155(.a(new_n250), .b(new_n249), .c(new_n248), .d(new_n229), .o1(new_n251));
  160nm_ficinv00aa1n08x5       g156(.clk(new_n251), .clkout(new_n252));
  xnrc02aa1n02x5               g157(.a(\b[24] ), .b(\a[25] ), .out0(new_n253));
  160nm_ficinv00aa1n08x5       g158(.clk(new_n253), .clkout(new_n254));
  xnbna2aa1n03x5               g159(.a(new_n254), .b(new_n246), .c(new_n252), .out0(\s[25] ));
  norp02aa1n02x5               g160(.a(\b[24] ), .b(\a[25] ), .o1(new_n256));
  160nm_ficinv00aa1n08x5       g161(.clk(new_n256), .clkout(new_n257));
  aoi012aa1n02x5               g162(.a(new_n253), .b(new_n246), .c(new_n252), .o1(new_n258));
  xnrc02aa1n02x5               g163(.a(\b[25] ), .b(\a[26] ), .out0(new_n259));
  nano22aa1n02x4               g164(.a(new_n258), .b(new_n257), .c(new_n259), .out0(new_n260));
  aoai13aa1n02x5               g165(.a(new_n254), .b(new_n251), .c(new_n173), .d(new_n245), .o1(new_n261));
  aoi012aa1n02x5               g166(.a(new_n259), .b(new_n261), .c(new_n257), .o1(new_n262));
  norp02aa1n02x5               g167(.a(new_n262), .b(new_n260), .o1(\s[26] ));
  norp02aa1n02x5               g168(.a(new_n259), .b(new_n253), .o1(new_n264));
  nano32aa1n02x4               g169(.a(new_n208), .b(new_n264), .c(new_n226), .d(new_n244), .out0(new_n265));
  aoai13aa1n02x5               g170(.a(new_n265), .b(new_n185), .c(new_n180), .d(new_n169), .o1(new_n266));
  oao003aa1n02x5               g171(.a(\a[26] ), .b(\b[25] ), .c(new_n257), .carry(new_n267));
  aobi12aa1n02x5               g172(.a(new_n267), .b(new_n251), .c(new_n264), .out0(new_n268));
  xorc02aa1n02x5               g173(.a(\a[27] ), .b(\b[26] ), .out0(new_n269));
  xnbna2aa1n03x5               g174(.a(new_n269), .b(new_n266), .c(new_n268), .out0(\s[27] ));
  norp02aa1n02x5               g175(.a(\b[26] ), .b(\a[27] ), .o1(new_n271));
  160nm_ficinv00aa1n08x5       g176(.clk(new_n271), .clkout(new_n272));
  aobi12aa1n02x5               g177(.a(new_n269), .b(new_n266), .c(new_n268), .out0(new_n273));
  xnrc02aa1n02x5               g178(.a(\b[27] ), .b(\a[28] ), .out0(new_n274));
  nano22aa1n02x4               g179(.a(new_n273), .b(new_n272), .c(new_n274), .out0(new_n275));
  aoai13aa1n02x5               g180(.a(new_n244), .b(new_n230), .c(new_n213), .d(new_n226), .o1(new_n276));
  160nm_ficinv00aa1n08x5       g181(.clk(new_n264), .clkout(new_n277));
  aoai13aa1n02x5               g182(.a(new_n267), .b(new_n277), .c(new_n276), .d(new_n250), .o1(new_n278));
  aoai13aa1n02x5               g183(.a(new_n269), .b(new_n278), .c(new_n173), .d(new_n265), .o1(new_n279));
  aoi012aa1n02x5               g184(.a(new_n274), .b(new_n279), .c(new_n272), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n280), .b(new_n275), .o1(\s[28] ));
  norb02aa1n02x5               g186(.a(new_n269), .b(new_n274), .out0(new_n282));
  aobi12aa1n02x5               g187(.a(new_n282), .b(new_n266), .c(new_n268), .out0(new_n283));
  oao003aa1n02x5               g188(.a(\a[28] ), .b(\b[27] ), .c(new_n272), .carry(new_n284));
  xnrc02aa1n02x5               g189(.a(\b[28] ), .b(\a[29] ), .out0(new_n285));
  nano22aa1n02x4               g190(.a(new_n283), .b(new_n284), .c(new_n285), .out0(new_n286));
  aoai13aa1n02x5               g191(.a(new_n282), .b(new_n278), .c(new_n173), .d(new_n265), .o1(new_n287));
  aoi012aa1n02x5               g192(.a(new_n285), .b(new_n287), .c(new_n284), .o1(new_n288));
  norp02aa1n02x5               g193(.a(new_n288), .b(new_n286), .o1(\s[29] ));
  xorb03aa1n02x5               g194(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g195(.a(new_n269), .b(new_n285), .c(new_n274), .out0(new_n291));
  aobi12aa1n02x5               g196(.a(new_n291), .b(new_n266), .c(new_n268), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .carry(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[29] ), .b(\a[30] ), .out0(new_n294));
  nano22aa1n02x4               g199(.a(new_n292), .b(new_n293), .c(new_n294), .out0(new_n295));
  aoai13aa1n02x5               g200(.a(new_n291), .b(new_n278), .c(new_n173), .d(new_n265), .o1(new_n296));
  aoi012aa1n02x5               g201(.a(new_n294), .b(new_n296), .c(new_n293), .o1(new_n297));
  norp02aa1n02x5               g202(.a(new_n297), .b(new_n295), .o1(\s[30] ));
  xnrc02aa1n02x5               g203(.a(\b[30] ), .b(\a[31] ), .out0(new_n299));
  norb02aa1n02x5               g204(.a(new_n291), .b(new_n294), .out0(new_n300));
  aobi12aa1n02x5               g205(.a(new_n300), .b(new_n266), .c(new_n268), .out0(new_n301));
  oao003aa1n02x5               g206(.a(\a[30] ), .b(\b[29] ), .c(new_n293), .carry(new_n302));
  nano22aa1n02x4               g207(.a(new_n301), .b(new_n299), .c(new_n302), .out0(new_n303));
  aoai13aa1n02x5               g208(.a(new_n300), .b(new_n278), .c(new_n173), .d(new_n265), .o1(new_n304));
  aoi012aa1n02x5               g209(.a(new_n299), .b(new_n304), .c(new_n302), .o1(new_n305));
  norp02aa1n02x5               g210(.a(new_n305), .b(new_n303), .o1(\s[31] ));
  xnrb03aa1n02x5               g211(.a(new_n100), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g212(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n308));
  xorb03aa1n02x5               g213(.a(new_n308), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g214(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  160nm_ficinv00aa1n08x5       g215(.clk(new_n107), .clkout(new_n311));
  oaoi13aa1n02x5               g216(.a(new_n113), .b(new_n116), .c(new_n311), .d(new_n114), .o1(new_n312));
  oai112aa1n02x5               g217(.a(new_n116), .b(new_n113), .c(new_n311), .d(new_n114), .o1(new_n313));
  norb02aa1n02x5               g218(.a(new_n313), .b(new_n312), .out0(\s[6] ));
  norp02aa1n02x5               g219(.a(new_n312), .b(new_n117), .o1(new_n315));
  xnrb03aa1n02x5               g220(.a(new_n315), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi13aa1n02x5               g221(.a(new_n110), .b(new_n111), .c(new_n312), .d(new_n117), .o1(new_n317));
  xnrb03aa1n02x5               g222(.a(new_n317), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g223(.a(new_n120), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


