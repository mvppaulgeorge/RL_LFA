// Benchmark "adder" written by ABC on Thu Jul 18 03:29:09 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n321, new_n324, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xorc02aa1n12x5               g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  nor042aa1n03x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  inv000aa1n02x5               g003(.a(new_n98), .o1(new_n99));
  inv040aa1d32x5               g004(.a(\a[4] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[3] ), .o1(new_n101));
  nor002aa1d32x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  tech160nm_fioaoi03aa1n03p5x5 g007(.a(new_n100), .b(new_n101), .c(new_n102), .o1(new_n103));
  tech160nm_fixnrc02aa1n02p5x5 g008(.a(\b[3] ), .b(\a[4] ), .out0(new_n104));
  nand22aa1n03x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nand02aa1d28x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  nor022aa1n04x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  norb03aa1n03x5               g012(.a(new_n106), .b(new_n105), .c(new_n107), .out0(new_n108));
  tech160nm_finand02aa1n05x5   g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nanb03aa1n03x5               g014(.a(new_n102), .b(new_n109), .c(new_n106), .out0(new_n110));
  oai013aa1n03x5               g015(.a(new_n103), .b(new_n108), .c(new_n110), .d(new_n104), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nand42aa1n08x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  norp02aa1n24x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nanp02aa1n02x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nona23aa1n03x5               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  xorc02aa1n12x5               g021(.a(\a[8] ), .b(\b[7] ), .out0(new_n117));
  xorc02aa1n12x5               g022(.a(\a[7] ), .b(\b[6] ), .out0(new_n118));
  nano22aa1n02x4               g023(.a(new_n116), .b(new_n117), .c(new_n118), .out0(new_n119));
  orn002aa1n03x5               g024(.a(\a[7] ), .b(\b[6] ), .o(new_n120));
  oaoi03aa1n09x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  oai012aa1n02x7               g026(.a(new_n113), .b(new_n114), .c(new_n112), .o1(new_n122));
  nanb03aa1n06x5               g027(.a(new_n122), .b(new_n117), .c(new_n118), .out0(new_n123));
  nanb02aa1n06x5               g028(.a(new_n121), .b(new_n123), .out0(new_n124));
  xorc02aa1n12x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n111), .d(new_n119), .o1(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n99), .out0(\s[10] ));
  inv030aa1n02x5               g032(.a(new_n103), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[4] ), .b(\b[3] ), .out0(new_n129));
  nona22aa1n06x5               g034(.a(new_n106), .b(new_n107), .c(new_n105), .out0(new_n130));
  nano22aa1n03x7               g035(.a(new_n102), .b(new_n106), .c(new_n109), .out0(new_n131));
  aoi013aa1n06x4               g036(.a(new_n128), .b(new_n131), .c(new_n130), .d(new_n129), .o1(new_n132));
  nanb03aa1n03x5               g037(.a(new_n116), .b(new_n118), .c(new_n117), .out0(new_n133));
  norb02aa1n02x5               g038(.a(new_n123), .b(new_n121), .out0(new_n134));
  oai012aa1n06x5               g039(.a(new_n134), .b(new_n133), .c(new_n132), .o1(new_n135));
  aoai13aa1n03x5               g040(.a(new_n97), .b(new_n98), .c(new_n135), .d(new_n125), .o1(new_n136));
  oai022aa1d24x5               g041(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n137));
  aob012aa1d15x5               g042(.a(new_n137), .b(\b[9] ), .c(\a[10] ), .out0(new_n138));
  nor002aa1d32x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  nand42aa1d28x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n136), .c(new_n138), .out0(\s[11] ));
  aob012aa1n03x5               g047(.a(new_n141), .b(new_n136), .c(new_n138), .out0(new_n143));
  nor002aa1d32x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n16x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  aoib12aa1n02x5               g051(.a(new_n139), .b(new_n145), .c(new_n144), .out0(new_n147));
  inv040aa1n09x5               g052(.a(new_n139), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n141), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n148), .b(new_n149), .c(new_n136), .d(new_n138), .o1(new_n150));
  aoi022aa1n03x5               g055(.a(new_n150), .b(new_n146), .c(new_n143), .d(new_n147), .o1(\s[12] ));
  nano23aa1d15x5               g056(.a(new_n139), .b(new_n144), .c(new_n145), .d(new_n140), .out0(new_n152));
  nanp03aa1d24x5               g057(.a(new_n152), .b(new_n97), .c(new_n125), .o1(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  nona23aa1n03x5               g059(.a(new_n145), .b(new_n140), .c(new_n139), .d(new_n144), .out0(new_n155));
  oaoi03aa1n09x5               g060(.a(\a[12] ), .b(\b[11] ), .c(new_n148), .o1(new_n156));
  oabi12aa1n02x7               g061(.a(new_n156), .b(new_n155), .c(new_n138), .out0(new_n157));
  tech160nm_fiao0012aa1n03p5x5 g062(.a(new_n157), .b(new_n135), .c(new_n154), .o(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  xnrc02aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .out0(new_n160));
  nanb02aa1n02x5               g065(.a(new_n160), .b(new_n158), .out0(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[13] ), .b(\a[14] ), .out0(new_n162));
  nor002aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n162), .b(new_n163), .out0(new_n164));
  oai012aa1n02x5               g069(.a(new_n161), .b(\b[12] ), .c(\a[13] ), .o1(new_n165));
  aboi22aa1n03x5               g070(.a(new_n162), .b(new_n165), .c(new_n161), .d(new_n164), .out0(\s[14] ));
  nor002aa1n04x5               g071(.a(new_n162), .b(new_n160), .o1(new_n167));
  aoai13aa1n03x5               g072(.a(new_n167), .b(new_n157), .c(new_n135), .d(new_n154), .o1(new_n168));
  inv000aa1d42x5               g073(.a(\a[14] ), .o1(new_n169));
  inv000aa1d42x5               g074(.a(\b[13] ), .o1(new_n170));
  tech160nm_fioaoi03aa1n03p5x5 g075(.a(new_n169), .b(new_n170), .c(new_n163), .o1(new_n171));
  nor042aa1d18x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nand02aa1d28x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(new_n174));
  xobna2aa1n03x5               g079(.a(new_n174), .b(new_n168), .c(new_n171), .out0(\s[15] ));
  ao0012aa1n03x7               g080(.a(new_n174), .b(new_n168), .c(new_n171), .o(new_n176));
  nor042aa1n06x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nand02aa1d10x5               g082(.a(\b[15] ), .b(\a[16] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  aoib12aa1n02x5               g084(.a(new_n172), .b(new_n178), .c(new_n177), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n172), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n174), .c(new_n168), .d(new_n171), .o1(new_n182));
  aboi22aa1n03x5               g087(.a(new_n179), .b(new_n182), .c(new_n176), .d(new_n180), .out0(\s[16] ));
  nano23aa1d15x5               g088(.a(new_n172), .b(new_n177), .c(new_n178), .d(new_n173), .out0(new_n184));
  nano22aa1n03x7               g089(.a(new_n153), .b(new_n167), .c(new_n184), .out0(new_n185));
  aoai13aa1n06x5               g090(.a(new_n185), .b(new_n124), .c(new_n111), .d(new_n119), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n171), .o1(new_n187));
  aoai13aa1n06x5               g092(.a(new_n184), .b(new_n187), .c(new_n157), .d(new_n167), .o1(new_n188));
  aoi012aa1n02x5               g093(.a(new_n177), .b(new_n172), .c(new_n178), .o1(new_n189));
  nanp03aa1d12x5               g094(.a(new_n186), .b(new_n188), .c(new_n189), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[16] ), .o1(new_n193));
  nanp02aa1n02x5               g098(.a(new_n193), .b(new_n192), .o1(new_n194));
  inv000aa1d42x5               g099(.a(new_n184), .o1(new_n195));
  tech160nm_fioaoi03aa1n03p5x5 g100(.a(\a[10] ), .b(\b[9] ), .c(new_n99), .o1(new_n196));
  aoai13aa1n02x5               g101(.a(new_n167), .b(new_n156), .c(new_n152), .d(new_n196), .o1(new_n197));
  aoai13aa1n03x5               g102(.a(new_n189), .b(new_n195), .c(new_n197), .d(new_n171), .o1(new_n198));
  tech160nm_fixorc02aa1n05x5   g103(.a(\a[17] ), .b(\b[16] ), .out0(new_n199));
  aoai13aa1n02x5               g104(.a(new_n199), .b(new_n198), .c(new_n135), .d(new_n185), .o1(new_n200));
  nor042aa1n12x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nand42aa1n03x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  norb02aa1n06x4               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  xnbna2aa1n03x5               g108(.a(new_n203), .b(new_n200), .c(new_n194), .out0(\s[18] ));
  and002aa1n02x5               g109(.a(new_n199), .b(new_n203), .o(new_n205));
  aoai13aa1n06x5               g110(.a(new_n202), .b(new_n201), .c(new_n192), .d(new_n193), .o1(new_n206));
  inv000aa1n02x5               g111(.a(new_n206), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  tech160nm_finand02aa1n05x5   g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nanb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  inv000aa1d42x5               g115(.a(new_n210), .o1(new_n211));
  aoai13aa1n06x5               g116(.a(new_n211), .b(new_n207), .c(new_n190), .d(new_n205), .o1(new_n212));
  aoi112aa1n02x5               g117(.a(new_n211), .b(new_n207), .c(new_n190), .d(new_n205), .o1(new_n213));
  norb02aa1n03x4               g118(.a(new_n212), .b(new_n213), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand42aa1n06x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  aoib12aa1n02x5               g123(.a(new_n208), .b(new_n217), .c(new_n216), .out0(new_n219));
  tech160nm_fioai012aa1n03p5x5 g124(.a(new_n212), .b(\b[18] ), .c(\a[19] ), .o1(new_n220));
  aoi022aa1n02x7               g125(.a(new_n220), .b(new_n218), .c(new_n212), .d(new_n219), .o1(\s[20] ));
  nano23aa1d15x5               g126(.a(new_n208), .b(new_n216), .c(new_n217), .d(new_n209), .out0(new_n222));
  nand23aa1d12x5               g127(.a(new_n222), .b(new_n199), .c(new_n203), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  nona23aa1n09x5               g129(.a(new_n217), .b(new_n209), .c(new_n208), .d(new_n216), .out0(new_n225));
  aoi012aa1n12x5               g130(.a(new_n216), .b(new_n208), .c(new_n217), .o1(new_n226));
  oai012aa1n09x5               g131(.a(new_n226), .b(new_n225), .c(new_n206), .o1(new_n227));
  xorc02aa1n02x5               g132(.a(\a[21] ), .b(\b[20] ), .out0(new_n228));
  aoai13aa1n06x5               g133(.a(new_n228), .b(new_n227), .c(new_n190), .d(new_n224), .o1(new_n229));
  aoi112aa1n02x5               g134(.a(new_n228), .b(new_n227), .c(new_n190), .d(new_n224), .o1(new_n230));
  norb02aa1n03x4               g135(.a(new_n229), .b(new_n230), .out0(\s[21] ));
  xorc02aa1n02x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  nor042aa1n03x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  norp02aa1n02x5               g138(.a(new_n232), .b(new_n233), .o1(new_n234));
  inv000aa1d42x5               g139(.a(\a[21] ), .o1(new_n235));
  oaib12aa1n06x5               g140(.a(new_n229), .b(\b[20] ), .c(new_n235), .out0(new_n236));
  aoi022aa1n03x5               g141(.a(new_n236), .b(new_n232), .c(new_n229), .d(new_n234), .o1(\s[22] ));
  inv040aa1d32x5               g142(.a(\a[22] ), .o1(new_n238));
  xroi22aa1d04x5               g143(.a(new_n235), .b(\b[20] ), .c(new_n238), .d(\b[21] ), .out0(new_n239));
  norb02aa1n09x5               g144(.a(new_n239), .b(new_n223), .out0(new_n240));
  inv000aa1n02x5               g145(.a(new_n226), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n239), .b(new_n241), .c(new_n222), .d(new_n207), .o1(new_n242));
  inv000aa1d42x5               g147(.a(\b[21] ), .o1(new_n243));
  oaoi03aa1n12x5               g148(.a(new_n238), .b(new_n243), .c(new_n233), .o1(new_n244));
  nanp02aa1n02x5               g149(.a(new_n242), .b(new_n244), .o1(new_n245));
  xorc02aa1n12x5               g150(.a(\a[23] ), .b(\b[22] ), .out0(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n245), .c(new_n190), .d(new_n240), .o1(new_n247));
  aoi112aa1n02x5               g152(.a(new_n246), .b(new_n245), .c(new_n190), .d(new_n240), .o1(new_n248));
  norb02aa1n03x4               g153(.a(new_n247), .b(new_n248), .out0(\s[23] ));
  nor042aa1n03x5               g154(.a(\b[23] ), .b(\a[24] ), .o1(new_n250));
  tech160nm_finand02aa1n05x5   g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  norb02aa1n06x4               g156(.a(new_n251), .b(new_n250), .out0(new_n252));
  norp02aa1n02x5               g157(.a(\b[22] ), .b(\a[23] ), .o1(new_n253));
  aoib12aa1n02x5               g158(.a(new_n253), .b(new_n251), .c(new_n250), .out0(new_n254));
  inv000aa1d42x5               g159(.a(\a[23] ), .o1(new_n255));
  oaib12aa1n06x5               g160(.a(new_n247), .b(\b[22] ), .c(new_n255), .out0(new_n256));
  aoi022aa1n02x7               g161(.a(new_n256), .b(new_n252), .c(new_n247), .d(new_n254), .o1(\s[24] ));
  nano32aa1n02x5               g162(.a(new_n223), .b(new_n252), .c(new_n239), .d(new_n246), .out0(new_n258));
  and002aa1n12x5               g163(.a(new_n246), .b(new_n252), .o(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  aoi012aa1n02x5               g165(.a(new_n250), .b(new_n253), .c(new_n251), .o1(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n260), .c(new_n242), .d(new_n244), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n190), .d(new_n258), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n262), .c(new_n190), .d(new_n258), .o1(new_n265));
  norb02aa1n03x4               g170(.a(new_n264), .b(new_n265), .out0(\s[25] ));
  xorc02aa1n02x5               g171(.a(\a[26] ), .b(\b[25] ), .out0(new_n267));
  norp02aa1n02x5               g172(.a(\b[24] ), .b(\a[25] ), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n267), .b(new_n268), .o1(new_n269));
  inv000aa1d42x5               g174(.a(\a[25] ), .o1(new_n270));
  oaib12aa1n06x5               g175(.a(new_n264), .b(\b[24] ), .c(new_n270), .out0(new_n271));
  aoi022aa1n03x5               g176(.a(new_n271), .b(new_n267), .c(new_n264), .d(new_n269), .o1(\s[26] ));
  inv000aa1d42x5               g177(.a(\a[26] ), .o1(new_n273));
  xroi22aa1d04x5               g178(.a(new_n270), .b(\b[24] ), .c(new_n273), .d(\b[25] ), .out0(new_n274));
  inv000aa1n02x5               g179(.a(new_n274), .o1(new_n275));
  nano23aa1n06x5               g180(.a(new_n223), .b(new_n275), .c(new_n259), .d(new_n239), .out0(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n198), .c(new_n135), .d(new_n185), .o1(new_n277));
  inv000aa1d42x5               g182(.a(\b[25] ), .o1(new_n278));
  oaoi03aa1n02x5               g183(.a(new_n273), .b(new_n278), .c(new_n268), .o1(new_n279));
  aobi12aa1n06x5               g184(.a(new_n279), .b(new_n262), .c(new_n274), .out0(new_n280));
  xorc02aa1n02x5               g185(.a(\a[27] ), .b(\b[26] ), .out0(new_n281));
  xnbna2aa1n03x5               g186(.a(new_n281), .b(new_n277), .c(new_n280), .out0(\s[27] ));
  inv000aa1d42x5               g187(.a(new_n244), .o1(new_n283));
  aoai13aa1n06x5               g188(.a(new_n259), .b(new_n283), .c(new_n227), .d(new_n239), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n279), .b(new_n275), .c(new_n284), .d(new_n261), .o1(new_n285));
  aoai13aa1n06x5               g190(.a(new_n281), .b(new_n285), .c(new_n190), .d(new_n276), .o1(new_n286));
  xorc02aa1n02x5               g191(.a(\a[28] ), .b(\b[27] ), .out0(new_n287));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  norp02aa1n02x5               g193(.a(new_n287), .b(new_n288), .o1(new_n289));
  inv000aa1d42x5               g194(.a(\a[27] ), .o1(new_n290));
  oaib12aa1n06x5               g195(.a(new_n286), .b(\b[26] ), .c(new_n290), .out0(new_n291));
  aoi022aa1n02x7               g196(.a(new_n291), .b(new_n287), .c(new_n286), .d(new_n289), .o1(\s[28] ));
  inv000aa1d42x5               g197(.a(\a[28] ), .o1(new_n293));
  xroi22aa1d04x5               g198(.a(new_n290), .b(\b[26] ), .c(new_n293), .d(\b[27] ), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n285), .c(new_n190), .d(new_n276), .o1(new_n295));
  oai022aa1n02x5               g200(.a(\a[27] ), .b(\b[26] ), .c(\b[27] ), .d(\a[28] ), .o1(new_n296));
  oaib12aa1n02x5               g201(.a(new_n296), .b(new_n293), .c(\b[27] ), .out0(new_n297));
  nanp02aa1n03x5               g202(.a(new_n295), .b(new_n297), .o1(new_n298));
  xorc02aa1n02x5               g203(.a(\a[29] ), .b(\b[28] ), .out0(new_n299));
  norb02aa1n02x5               g204(.a(new_n297), .b(new_n299), .out0(new_n300));
  aoi022aa1n02x7               g205(.a(new_n298), .b(new_n299), .c(new_n295), .d(new_n300), .o1(\s[29] ));
  xorb03aa1n02x5               g206(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g207(.a(new_n281), .b(new_n299), .c(new_n287), .o(new_n303));
  aoai13aa1n03x5               g208(.a(new_n303), .b(new_n285), .c(new_n190), .d(new_n276), .o1(new_n304));
  oao003aa1n02x5               g209(.a(\a[29] ), .b(\b[28] ), .c(new_n297), .carry(new_n305));
  nand42aa1n02x5               g210(.a(new_n304), .b(new_n305), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  norb02aa1n02x5               g212(.a(new_n305), .b(new_n307), .out0(new_n308));
  aoi022aa1n02x7               g213(.a(new_n306), .b(new_n307), .c(new_n304), .d(new_n308), .o1(\s[30] ));
  nanb02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  nanb02aa1n02x5               g215(.a(\a[31] ), .b(\b[30] ), .out0(new_n311));
  and003aa1n02x5               g216(.a(new_n294), .b(new_n307), .c(new_n299), .o(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n285), .c(new_n190), .d(new_n276), .o1(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n314));
  aoi022aa1n03x5               g219(.a(new_n313), .b(new_n314), .c(new_n311), .d(new_n310), .o1(new_n315));
  aobi12aa1n06x5               g220(.a(new_n312), .b(new_n277), .c(new_n280), .out0(new_n316));
  nano32aa1n02x4               g221(.a(new_n316), .b(new_n314), .c(new_n310), .d(new_n311), .out0(new_n317));
  nor002aa1n02x5               g222(.a(new_n315), .b(new_n317), .o1(\s[31] ));
  norb02aa1n02x5               g223(.a(new_n109), .b(new_n102), .out0(new_n319));
  xobna2aa1n03x5               g224(.a(new_n319), .b(new_n130), .c(new_n106), .out0(\s[3] ));
  aoi112aa1n02x5               g225(.a(new_n102), .b(new_n129), .c(new_n131), .d(new_n130), .o1(new_n321));
  oaoi13aa1n02x5               g226(.a(new_n321), .b(new_n111), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g228(.a(\a[5] ), .b(\b[4] ), .c(new_n132), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoi012aa1n02x5               g230(.a(new_n112), .b(new_n324), .c(new_n113), .o1(new_n326));
  xnrc02aa1n02x5               g231(.a(new_n326), .b(new_n118), .out0(\s[7] ));
  aoai13aa1n02x5               g232(.a(new_n118), .b(new_n112), .c(new_n324), .d(new_n113), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n117), .b(new_n328), .c(new_n120), .out0(\s[8] ));
  xorb03aa1n02x5               g234(.a(new_n135), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


