// Benchmark "adder" written by ABC on Wed Jul 17 18:00:18 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n322, new_n323, new_n326,
    new_n328, new_n330;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  oai022aa1d24x5               g003(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n99));
  nor042aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  nand42aa1n10x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  norb02aa1n12x5               g006(.a(new_n101), .b(new_n100), .out0(new_n102));
  nor042aa1n03x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  aoi022aa1n12x5               g008(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n104));
  oaoi13aa1n12x5               g009(.a(new_n99), .b(new_n102), .c(new_n104), .d(new_n103), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nand42aa1d28x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  nor002aa1d24x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  norb02aa1n15x5               g014(.a(new_n108), .b(new_n109), .out0(new_n110));
  nand23aa1n06x5               g015(.a(new_n110), .b(new_n106), .c(new_n107), .o1(new_n111));
  inv040aa1d32x5               g016(.a(\a[8] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\b[7] ), .o1(new_n113));
  nand42aa1n03x5               g018(.a(new_n113), .b(new_n112), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n12x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  norb02aa1n03x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nor042aa1n06x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nand42aa1d28x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  norb02aa1n03x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  nand23aa1n06x5               g025(.a(new_n117), .b(new_n120), .c(new_n114), .o1(new_n121));
  aoi022aa1d18x5               g026(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n122));
  nand02aa1n02x5               g027(.a(new_n109), .b(new_n119), .o1(new_n123));
  nona22aa1n03x5               g028(.a(new_n123), .b(new_n118), .c(new_n115), .out0(new_n124));
  aoi022aa1n09x5               g029(.a(new_n124), .b(new_n122), .c(new_n112), .d(new_n113), .o1(new_n125));
  oai013aa1d12x5               g030(.a(new_n125), .b(new_n105), .c(new_n121), .d(new_n111), .o1(new_n126));
  tech160nm_fioaoi03aa1n03p5x5 g031(.a(new_n97), .b(new_n98), .c(new_n126), .o1(new_n127));
  orn002aa1n02x7               g032(.a(\a[10] ), .b(\b[9] ), .o(new_n128));
  nand42aa1n08x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n127), .b(new_n129), .c(new_n128), .out0(\s[10] ));
  xnrc02aa1n02x5               g035(.a(\b[10] ), .b(\a[11] ), .out0(new_n131));
  nanp02aa1n03x5               g036(.a(new_n127), .b(new_n128), .o1(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n131), .b(new_n132), .c(new_n129), .out0(\s[11] ));
  norp02aa1n02x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  xorc02aa1n12x5               g039(.a(\a[11] ), .b(\b[10] ), .out0(new_n135));
  nor042aa1n02x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanp02aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  aoi113aa1n02x5               g043(.a(new_n134), .b(new_n138), .c(new_n132), .d(new_n135), .e(new_n129), .o1(new_n139));
  aoi013aa1n03x5               g044(.a(new_n134), .b(new_n132), .c(new_n135), .d(new_n129), .o1(new_n140));
  norb02aa1n02x5               g045(.a(new_n138), .b(new_n140), .out0(new_n141));
  norp02aa1n02x5               g046(.a(new_n141), .b(new_n139), .o1(\s[12] ));
  inv000aa1d42x5               g047(.a(new_n99), .o1(new_n143));
  nanb02aa1n02x5               g048(.a(new_n100), .b(new_n101), .out0(new_n144));
  inv000aa1n02x5               g049(.a(new_n103), .o1(new_n145));
  nand42aa1n03x5               g050(.a(\b[0] ), .b(\a[1] ), .o1(new_n146));
  aob012aa1n02x5               g051(.a(new_n146), .b(\b[1] ), .c(\a[2] ), .out0(new_n147));
  aoai13aa1n04x5               g052(.a(new_n143), .b(new_n144), .c(new_n147), .d(new_n145), .o1(new_n148));
  nano32aa1n02x4               g053(.a(new_n109), .b(new_n108), .c(new_n107), .d(new_n106), .out0(new_n149));
  inv000aa1d42x5               g054(.a(new_n115), .o1(new_n150));
  nanb02aa1n02x5               g055(.a(new_n118), .b(new_n119), .out0(new_n151));
  nano32aa1n02x4               g056(.a(new_n151), .b(new_n150), .c(new_n114), .d(new_n116), .out0(new_n152));
  nanp03aa1n03x5               g057(.a(new_n148), .b(new_n149), .c(new_n152), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(new_n98), .b(new_n97), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(\b[8] ), .b(\a[9] ), .o1(new_n155));
  tech160nm_fixorc02aa1n03p5x5 g060(.a(\a[10] ), .b(\b[9] ), .out0(new_n156));
  nano22aa1n03x7               g061(.a(new_n136), .b(new_n129), .c(new_n137), .out0(new_n157));
  nanp02aa1n02x5               g062(.a(new_n157), .b(new_n135), .o1(new_n158));
  nano32aa1n02x5               g063(.a(new_n158), .b(new_n156), .c(new_n155), .d(new_n154), .out0(new_n159));
  inv000aa1n02x5               g064(.a(new_n159), .o1(new_n160));
  aoi112aa1n02x5               g065(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n161));
  oai112aa1n03x5               g066(.a(new_n128), .b(new_n129), .c(\b[8] ), .d(\a[9] ), .o1(new_n162));
  nanp03aa1n03x5               g067(.a(new_n157), .b(new_n162), .c(new_n135), .o1(new_n163));
  nona22aa1n06x5               g068(.a(new_n163), .b(new_n161), .c(new_n136), .out0(new_n164));
  inv040aa1n03x5               g069(.a(new_n164), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n165), .b(new_n160), .c(new_n153), .d(new_n125), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n06x5               g072(.a(\b[13] ), .b(\a[14] ), .o1(new_n168));
  and002aa1n12x5               g073(.a(\b[13] ), .b(\a[14] ), .o(new_n169));
  norp02aa1n02x5               g074(.a(new_n169), .b(new_n168), .o1(new_n170));
  nor042aa1n06x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nanp02aa1n02x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  aoi012aa1n02x5               g077(.a(new_n171), .b(new_n166), .c(new_n172), .o1(new_n173));
  xnrc02aa1n02x5               g078(.a(new_n173), .b(new_n170), .out0(\s[14] ));
  norb02aa1n02x5               g079(.a(new_n172), .b(new_n171), .out0(new_n175));
  oabi12aa1n18x5               g080(.a(new_n169), .b(new_n171), .c(new_n168), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n176), .o1(new_n177));
  aoi013aa1n06x4               g082(.a(new_n177), .b(new_n166), .c(new_n175), .d(new_n170), .o1(new_n178));
  nor002aa1n03x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  inv000aa1n02x5               g084(.a(new_n179), .o1(new_n180));
  nand02aa1d28x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n178), .b(new_n181), .c(new_n180), .out0(\s[15] ));
  nanb02aa1n02x5               g087(.a(new_n179), .b(new_n181), .out0(new_n183));
  nor002aa1n16x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nanp02aa1n12x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nanb02aa1n02x5               g090(.a(new_n184), .b(new_n185), .out0(new_n186));
  oaoi13aa1n09x5               g091(.a(new_n186), .b(new_n180), .c(new_n178), .d(new_n183), .o1(new_n187));
  oai112aa1n03x5               g092(.a(new_n186), .b(new_n180), .c(new_n178), .d(new_n183), .o1(new_n188));
  norb02aa1n03x4               g093(.a(new_n188), .b(new_n187), .out0(\s[16] ));
  nor043aa1n03x5               g094(.a(new_n169), .b(new_n168), .c(new_n171), .o1(new_n190));
  nano23aa1n06x5               g095(.a(new_n179), .b(new_n184), .c(new_n185), .d(new_n181), .out0(new_n191));
  nand23aa1n03x5               g096(.a(new_n191), .b(new_n172), .c(new_n190), .o1(new_n192));
  inv040aa1n02x5               g097(.a(new_n192), .o1(new_n193));
  inv000aa1d42x5               g098(.a(new_n184), .o1(new_n194));
  nanp02aa1n02x5               g099(.a(new_n185), .b(new_n181), .o1(new_n195));
  aoai13aa1n09x5               g100(.a(new_n194), .b(new_n195), .c(new_n176), .d(new_n180), .o1(new_n196));
  aoi012aa1d18x5               g101(.a(new_n196), .b(new_n164), .c(new_n193), .o1(new_n197));
  nanp03aa1n02x5               g102(.a(new_n156), .b(new_n154), .c(new_n155), .o1(new_n198));
  nona32aa1d24x5               g103(.a(new_n126), .b(new_n192), .c(new_n198), .d(new_n158), .out0(new_n199));
  nand22aa1n09x5               g104(.a(new_n199), .b(new_n197), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g106(.a(\a[18] ), .o1(new_n202));
  inv040aa1d32x5               g107(.a(\a[17] ), .o1(new_n203));
  inv000aa1d42x5               g108(.a(\b[16] ), .o1(new_n204));
  oaoi03aa1n03x5               g109(.a(new_n203), .b(new_n204), .c(new_n200), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[17] ), .c(new_n202), .out0(\s[18] ));
  xroi22aa1d06x4               g111(.a(new_n203), .b(\b[16] ), .c(new_n202), .d(\b[17] ), .out0(new_n207));
  nanp02aa1n02x5               g112(.a(new_n204), .b(new_n203), .o1(new_n208));
  oaoi03aa1n12x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n208), .o1(new_n209));
  nor022aa1n08x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nanp02aa1n06x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  norb02aa1n02x5               g116(.a(new_n211), .b(new_n210), .out0(new_n212));
  aoai13aa1n06x5               g117(.a(new_n212), .b(new_n209), .c(new_n200), .d(new_n207), .o1(new_n213));
  aoi112aa1n02x5               g118(.a(new_n212), .b(new_n209), .c(new_n200), .d(new_n207), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n213), .b(new_n214), .out0(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n08x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand42aa1n04x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  nona22aa1n03x5               g124(.a(new_n213), .b(new_n219), .c(new_n210), .out0(new_n220));
  orn002aa1n24x5               g125(.a(\a[19] ), .b(\b[18] ), .o(new_n221));
  aobi12aa1n03x5               g126(.a(new_n219), .b(new_n213), .c(new_n221), .out0(new_n222));
  norb02aa1n03x4               g127(.a(new_n220), .b(new_n222), .out0(\s[20] ));
  nano23aa1n09x5               g128(.a(new_n210), .b(new_n217), .c(new_n218), .d(new_n211), .out0(new_n224));
  nanp02aa1n02x5               g129(.a(new_n207), .b(new_n224), .o1(new_n225));
  oai022aa1n02x7               g130(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n226));
  oaib12aa1n09x5               g131(.a(new_n226), .b(new_n202), .c(\b[17] ), .out0(new_n227));
  nona23aa1n09x5               g132(.a(new_n218), .b(new_n211), .c(new_n210), .d(new_n217), .out0(new_n228));
  oaoi03aa1n09x5               g133(.a(\a[20] ), .b(\b[19] ), .c(new_n221), .o1(new_n229));
  oabi12aa1n18x5               g134(.a(new_n229), .b(new_n228), .c(new_n227), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n225), .c(new_n199), .d(new_n197), .o1(new_n232));
  xorb03aa1n02x5               g137(.a(new_n232), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(\b[20] ), .b(\a[21] ), .o1(new_n235));
  xorc02aa1n02x5               g140(.a(\a[22] ), .b(\b[21] ), .out0(new_n236));
  aoi112aa1n03x5               g141(.a(new_n234), .b(new_n236), .c(new_n232), .d(new_n235), .o1(new_n237));
  aoai13aa1n04x5               g142(.a(new_n236), .b(new_n234), .c(new_n232), .d(new_n235), .o1(new_n238));
  norb02aa1n03x4               g143(.a(new_n238), .b(new_n237), .out0(\s[22] ));
  inv000aa1d42x5               g144(.a(\a[21] ), .o1(new_n240));
  inv040aa1d32x5               g145(.a(\a[22] ), .o1(new_n241));
  xroi22aa1d06x4               g146(.a(new_n240), .b(\b[20] ), .c(new_n241), .d(\b[21] ), .out0(new_n242));
  nand03aa1n06x5               g147(.a(new_n242), .b(new_n207), .c(new_n224), .o1(new_n243));
  inv000aa1d42x5               g148(.a(\b[21] ), .o1(new_n244));
  oao003aa1n02x5               g149(.a(new_n241), .b(new_n244), .c(new_n234), .carry(new_n245));
  aoi012aa1n02x5               g150(.a(new_n245), .b(new_n230), .c(new_n242), .o1(new_n246));
  aoai13aa1n06x5               g151(.a(new_n246), .b(new_n243), .c(new_n199), .d(new_n197), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  xorc02aa1n12x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  xorc02aa1n12x5               g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  aoi112aa1n03x5               g156(.a(new_n249), .b(new_n251), .c(new_n247), .d(new_n250), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n251), .b(new_n249), .c(new_n247), .d(new_n250), .o1(new_n253));
  norb02aa1n03x4               g158(.a(new_n253), .b(new_n252), .out0(\s[24] ));
  and002aa1n02x7               g159(.a(new_n251), .b(new_n250), .o(new_n255));
  inv030aa1n02x5               g160(.a(new_n255), .o1(new_n256));
  nano32aa1n02x5               g161(.a(new_n256), .b(new_n242), .c(new_n207), .d(new_n224), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n242), .b(new_n229), .c(new_n224), .d(new_n209), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n245), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n260));
  oab012aa1n02x4               g165(.a(new_n260), .b(\a[24] ), .c(\b[23] ), .out0(new_n261));
  aoai13aa1n04x5               g166(.a(new_n261), .b(new_n256), .c(new_n258), .d(new_n259), .o1(new_n262));
  xorc02aa1n02x5               g167(.a(\a[25] ), .b(\b[24] ), .out0(new_n263));
  aoai13aa1n06x5               g168(.a(new_n263), .b(new_n262), .c(new_n200), .d(new_n257), .o1(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n262), .c(new_n200), .d(new_n257), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n264), .b(new_n265), .out0(\s[25] ));
  nor042aa1n03x5               g171(.a(\b[24] ), .b(\a[25] ), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  nona22aa1n03x5               g173(.a(new_n264), .b(new_n268), .c(new_n267), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n267), .o1(new_n270));
  aobi12aa1n02x7               g175(.a(new_n268), .b(new_n264), .c(new_n270), .out0(new_n271));
  norb02aa1n03x4               g176(.a(new_n269), .b(new_n271), .out0(\s[26] ));
  norp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  nanp02aa1n02x5               g178(.a(\b[26] ), .b(\a[27] ), .o1(new_n274));
  norb02aa1n02x5               g179(.a(new_n274), .b(new_n273), .out0(new_n275));
  inv040aa1d30x5               g180(.a(\a[25] ), .o1(new_n276));
  inv040aa1d32x5               g181(.a(\a[26] ), .o1(new_n277));
  xroi22aa1d06x4               g182(.a(new_n276), .b(\b[24] ), .c(new_n277), .d(\b[25] ), .out0(new_n278));
  nano22aa1d15x5               g183(.a(new_n243), .b(new_n255), .c(new_n278), .out0(new_n279));
  nanp02aa1n06x5               g184(.a(new_n200), .b(new_n279), .o1(new_n280));
  oao003aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .c(new_n270), .carry(new_n281));
  aobi12aa1n06x5               g186(.a(new_n281), .b(new_n262), .c(new_n278), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n275), .b(new_n280), .c(new_n282), .out0(\s[27] ));
  inv000aa1n06x5               g188(.a(new_n273), .o1(new_n284));
  inv020aa1n03x5               g189(.a(new_n279), .o1(new_n285));
  aoi012aa1n12x5               g190(.a(new_n285), .b(new_n199), .c(new_n197), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n255), .b(new_n245), .c(new_n230), .d(new_n242), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n278), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n281), .b(new_n288), .c(new_n287), .d(new_n261), .o1(new_n289));
  oaih12aa1n02x5               g194(.a(new_n274), .b(new_n289), .c(new_n286), .o1(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  tech160nm_fiaoi012aa1n02p5x5 g196(.a(new_n291), .b(new_n290), .c(new_n284), .o1(new_n292));
  aobi12aa1n02x7               g197(.a(new_n274), .b(new_n280), .c(new_n282), .out0(new_n293));
  nano22aa1n03x5               g198(.a(new_n293), .b(new_n284), .c(new_n291), .out0(new_n294));
  norp02aa1n03x5               g199(.a(new_n292), .b(new_n294), .o1(\s[28] ));
  nano22aa1n02x4               g200(.a(new_n291), .b(new_n284), .c(new_n274), .out0(new_n296));
  oaih12aa1n02x5               g201(.a(new_n296), .b(new_n289), .c(new_n286), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .c(new_n284), .carry(new_n298));
  xnrc02aa1n02x5               g203(.a(\b[28] ), .b(\a[29] ), .out0(new_n299));
  tech160nm_fiaoi012aa1n02p5x5 g204(.a(new_n299), .b(new_n297), .c(new_n298), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n296), .b(new_n280), .c(new_n282), .out0(new_n301));
  nano22aa1n02x4               g206(.a(new_n301), .b(new_n298), .c(new_n299), .out0(new_n302));
  norp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[29] ));
  xorb03aa1n02x5               g208(.a(new_n146), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g209(.a(new_n275), .b(new_n299), .c(new_n291), .out0(new_n305));
  oaih12aa1n02x5               g210(.a(new_n305), .b(new_n289), .c(new_n286), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[29] ), .b(\b[28] ), .c(new_n298), .carry(new_n307));
  xnrc02aa1n02x5               g212(.a(\b[29] ), .b(\a[30] ), .out0(new_n308));
  tech160nm_fiaoi012aa1n02p5x5 g213(.a(new_n308), .b(new_n306), .c(new_n307), .o1(new_n309));
  aobi12aa1n02x7               g214(.a(new_n305), .b(new_n280), .c(new_n282), .out0(new_n310));
  nano22aa1n02x4               g215(.a(new_n310), .b(new_n307), .c(new_n308), .out0(new_n311));
  norp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[30] ));
  xnrc02aa1n02x5               g217(.a(\b[30] ), .b(\a[31] ), .out0(new_n313));
  norb03aa1n02x5               g218(.a(new_n296), .b(new_n308), .c(new_n299), .out0(new_n314));
  oaih12aa1n02x5               g219(.a(new_n314), .b(new_n289), .c(new_n286), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .c(new_n307), .carry(new_n316));
  tech160nm_fiaoi012aa1n02p5x5 g221(.a(new_n313), .b(new_n315), .c(new_n316), .o1(new_n317));
  aobi12aa1n02x7               g222(.a(new_n314), .b(new_n280), .c(new_n282), .out0(new_n318));
  nano22aa1n03x5               g223(.a(new_n318), .b(new_n313), .c(new_n316), .out0(new_n319));
  norp02aa1n03x5               g224(.a(new_n317), .b(new_n319), .o1(\s[31] ));
  xnbna2aa1n03x5               g225(.a(new_n102), .b(new_n147), .c(new_n145), .out0(\s[3] ));
  xorc02aa1n02x5               g226(.a(\a[4] ), .b(\b[3] ), .out0(new_n322));
  oaoi13aa1n02x5               g227(.a(new_n100), .b(new_n101), .c(new_n104), .d(new_n103), .o1(new_n323));
  mtn022aa1n02x5               g228(.a(new_n148), .b(new_n323), .sa(new_n322), .o1(\s[4] ));
  xobna2aa1n03x5               g229(.a(new_n110), .b(new_n148), .c(new_n107), .out0(\s[5] ));
  aoai13aa1n06x5               g230(.a(new_n110), .b(new_n105), .c(\a[4] ), .d(\b[3] ), .o1(new_n326));
  xnbna2aa1n03x5               g231(.a(new_n151), .b(new_n326), .c(new_n108), .out0(\s[6] ));
  aoi013aa1n02x4               g232(.a(new_n118), .b(new_n326), .c(new_n119), .d(new_n108), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n150), .c(new_n116), .out0(\s[7] ));
  oaoi03aa1n03x5               g234(.a(\a[7] ), .b(\b[6] ), .c(new_n328), .o1(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g236(.a(new_n126), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


