// Benchmark "adder" written by ABC on Wed Jul 17 23:26:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n320, new_n321, new_n323, new_n324,
    new_n325, new_n327, new_n328, new_n329, new_n331, new_n332, new_n333,
    new_n335, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n10x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1d24x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nand42aa1n04x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nor022aa1n16x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand42aa1n20x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nanb03aa1n06x5               g008(.a(new_n102), .b(new_n103), .c(new_n101), .out0(new_n104));
  nand22aa1n06x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nor022aa1n08x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  norb03aa1d15x5               g011(.a(new_n103), .b(new_n106), .c(new_n105), .out0(new_n107));
  norp02aa1n03x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  nor002aa1n02x5               g013(.a(new_n108), .b(new_n102), .o1(new_n109));
  oai012aa1n04x7               g014(.a(new_n109), .b(new_n107), .c(new_n104), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand42aa1n04x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand02aa1n03x5               g017(.a(\b[3] ), .b(\a[4] ), .o1(new_n113));
  nanp03aa1n02x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .o1(new_n114));
  xnrc02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .out0(new_n115));
  nor002aa1d24x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  oab012aa1n06x5               g021(.a(new_n116), .b(\a[6] ), .c(\b[5] ), .out0(new_n117));
  norp02aa1n24x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  aoi012aa1n02x5               g023(.a(new_n118), .b(\a[6] ), .c(\b[5] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n117), .b(new_n119), .o1(new_n120));
  nona32aa1n09x5               g025(.a(new_n110), .b(new_n120), .c(new_n115), .d(new_n114), .out0(new_n121));
  xorc02aa1n12x5               g026(.a(\a[8] ), .b(\b[7] ), .out0(new_n122));
  inv000aa1n02x5               g027(.a(new_n117), .o1(new_n123));
  inv000aa1d42x5               g028(.a(new_n118), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  nand22aa1n02x5               g030(.a(\b[5] ), .b(\a[6] ), .o1(new_n126));
  nano22aa1n03x7               g031(.a(new_n118), .b(new_n112), .c(new_n126), .out0(new_n127));
  aoi013aa1n09x5               g032(.a(new_n125), .b(new_n127), .c(new_n122), .d(new_n123), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(new_n121), .b(new_n128), .o1(new_n129));
  xnrc02aa1n12x5               g034(.a(\b[8] ), .b(\a[9] ), .out0(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  aoai13aa1n02x5               g036(.a(new_n99), .b(new_n100), .c(new_n129), .d(new_n131), .o1(new_n132));
  nona22aa1n02x4               g037(.a(new_n98), .b(new_n100), .c(new_n97), .out0(new_n133));
  tech160nm_fiao0012aa1n02p5x5 g038(.a(new_n133), .b(new_n129), .c(new_n131), .o(new_n134));
  nanp02aa1n02x5               g039(.a(new_n134), .b(new_n132), .o1(\s[10] ));
  nor002aa1d32x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  inv040aa1n08x5               g041(.a(new_n136), .o1(new_n137));
  nanp02aa1n06x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  aoi022aa1n02x5               g043(.a(new_n134), .b(new_n98), .c(new_n138), .d(new_n137), .o1(new_n139));
  nano22aa1n02x4               g044(.a(new_n136), .b(new_n98), .c(new_n138), .out0(new_n140));
  aoai13aa1n02x5               g045(.a(new_n140), .b(new_n133), .c(new_n129), .d(new_n131), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n139), .out0(\s[11] ));
  norp02aa1n24x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nanp02aa1n09x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n02x5               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  xnbna2aa1n03x5               g050(.a(new_n145), .b(new_n141), .c(new_n137), .out0(\s[12] ));
  nona23aa1n02x4               g051(.a(new_n144), .b(new_n138), .c(new_n136), .d(new_n143), .out0(new_n147));
  nona22aa1n02x4               g052(.a(new_n131), .b(new_n147), .c(new_n99), .out0(new_n148));
  oaih12aa1n12x5               g053(.a(new_n144), .b(new_n143), .c(new_n136), .o1(new_n149));
  nanb03aa1d18x5               g054(.a(new_n143), .b(new_n144), .c(new_n138), .out0(new_n150));
  oai112aa1n06x5               g055(.a(new_n137), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n151));
  oai012aa1d24x5               g056(.a(new_n149), .b(new_n151), .c(new_n150), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  aoai13aa1n04x5               g058(.a(new_n153), .b(new_n148), .c(new_n121), .d(new_n128), .o1(new_n154));
  xorb03aa1n02x5               g059(.a(new_n154), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  nand02aa1d06x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nanp03aa1n02x5               g063(.a(new_n154), .b(new_n157), .c(new_n158), .o1(new_n159));
  norp02aa1n12x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n08x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnbna2aa1n03x5               g067(.a(new_n162), .b(new_n159), .c(new_n157), .out0(\s[14] ));
  nona23aa1d24x5               g068(.a(new_n161), .b(new_n158), .c(new_n156), .d(new_n160), .out0(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  oaoi03aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n166));
  nor002aa1n04x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n04x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n06x4               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  aoai13aa1n02x5               g074(.a(new_n169), .b(new_n166), .c(new_n154), .d(new_n165), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n169), .b(new_n166), .c(new_n154), .d(new_n165), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(\s[15] ));
  inv000aa1d42x5               g077(.a(\a[15] ), .o1(new_n173));
  oaib12aa1n02x5               g078(.a(new_n170), .b(\b[14] ), .c(new_n173), .out0(new_n174));
  nor002aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand02aa1d06x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  norb02aa1n06x4               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  norp02aa1n02x5               g082(.a(new_n177), .b(new_n167), .o1(new_n178));
  aoi022aa1n02x5               g083(.a(new_n174), .b(new_n177), .c(new_n170), .d(new_n178), .o1(\s[16] ));
  nano22aa1d15x5               g084(.a(new_n164), .b(new_n169), .c(new_n177), .out0(new_n180));
  nona32aa1n09x5               g085(.a(new_n180), .b(new_n147), .c(new_n130), .d(new_n99), .out0(new_n181));
  tech160nm_fiao0012aa1n02p5x5 g086(.a(new_n181), .b(new_n121), .c(new_n128), .o(new_n182));
  nanb03aa1n02x5               g087(.a(new_n175), .b(new_n176), .c(new_n168), .out0(new_n183));
  oai122aa1n02x7               g088(.a(new_n161), .b(new_n160), .c(new_n156), .d(\b[14] ), .e(\a[15] ), .o1(new_n184));
  aoi012aa1n02x5               g089(.a(new_n175), .b(new_n167), .c(new_n176), .o1(new_n185));
  oai012aa1n06x5               g090(.a(new_n185), .b(new_n184), .c(new_n183), .o1(new_n186));
  aoi012aa1d18x5               g091(.a(new_n186), .b(new_n152), .c(new_n180), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n181), .c(new_n121), .d(new_n128), .o1(new_n188));
  xorc02aa1n12x5               g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  aoi112aa1n02x5               g094(.a(new_n189), .b(new_n186), .c(new_n152), .d(new_n180), .o1(new_n190));
  aoi022aa1n02x5               g095(.a(new_n182), .b(new_n190), .c(new_n188), .d(new_n189), .o1(\s[17] ));
  norp02aa1n02x5               g096(.a(\b[16] ), .b(\a[17] ), .o1(new_n192));
  xorc02aa1n12x5               g097(.a(\a[18] ), .b(\b[17] ), .out0(new_n193));
  aoai13aa1n02x5               g098(.a(new_n193), .b(new_n192), .c(new_n188), .d(new_n189), .o1(new_n194));
  aoi112aa1n02x5               g099(.a(new_n192), .b(new_n193), .c(new_n188), .d(new_n189), .o1(new_n195));
  norb02aa1n02x5               g100(.a(new_n194), .b(new_n195), .out0(\s[18] ));
  and002aa1n02x5               g101(.a(new_n193), .b(new_n189), .o(new_n197));
  nand22aa1n03x5               g102(.a(new_n188), .b(new_n197), .o1(new_n198));
  nanp02aa1n02x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  oai022aa1n04x5               g104(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n200));
  nanp02aa1n02x5               g105(.a(new_n200), .b(new_n199), .o1(new_n201));
  xorc02aa1n12x5               g106(.a(\a[19] ), .b(\b[18] ), .out0(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n198), .c(new_n201), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g109(.a(new_n202), .b(new_n198), .c(new_n201), .out0(new_n205));
  inv000aa1d42x5               g110(.a(\a[19] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[18] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(new_n207), .b(new_n206), .o1(new_n208));
  inv040aa1n02x5               g113(.a(new_n202), .o1(new_n209));
  aoai13aa1n02x5               g114(.a(new_n208), .b(new_n209), .c(new_n198), .d(new_n201), .o1(new_n210));
  xorc02aa1n02x5               g115(.a(\a[20] ), .b(\b[19] ), .out0(new_n211));
  inv040aa1d32x5               g116(.a(\a[20] ), .o1(new_n212));
  inv000aa1d42x5               g117(.a(\b[19] ), .o1(new_n213));
  nanp02aa1n04x5               g118(.a(new_n213), .b(new_n212), .o1(new_n214));
  nand42aa1n02x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  aoi022aa1n02x5               g120(.a(new_n214), .b(new_n215), .c(new_n207), .d(new_n206), .o1(new_n216));
  aoi022aa1n03x5               g121(.a(new_n210), .b(new_n211), .c(new_n205), .d(new_n216), .o1(\s[20] ));
  nano32aa1n03x7               g122(.a(new_n209), .b(new_n211), .c(new_n189), .d(new_n193), .out0(new_n218));
  oai112aa1n03x5               g123(.a(new_n214), .b(new_n215), .c(new_n207), .d(new_n206), .o1(new_n219));
  nand23aa1n02x5               g124(.a(new_n200), .b(new_n208), .c(new_n199), .o1(new_n220));
  aoi112aa1n02x7               g125(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n221));
  norb02aa1n06x4               g126(.a(new_n214), .b(new_n221), .out0(new_n222));
  oai012aa1n06x5               g127(.a(new_n222), .b(new_n220), .c(new_n219), .o1(new_n223));
  xorc02aa1n02x5               g128(.a(\a[21] ), .b(\b[20] ), .out0(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n223), .c(new_n188), .d(new_n218), .o1(new_n225));
  aoi112aa1n02x5               g130(.a(new_n224), .b(new_n223), .c(new_n188), .d(new_n218), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n225), .b(new_n226), .out0(\s[21] ));
  inv000aa1d42x5               g132(.a(\a[21] ), .o1(new_n228));
  oaib12aa1n03x5               g133(.a(new_n225), .b(\b[20] ), .c(new_n228), .out0(new_n229));
  xorc02aa1n02x5               g134(.a(\a[22] ), .b(\b[21] ), .out0(new_n230));
  norp02aa1n02x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norp02aa1n02x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  aoi022aa1n02x5               g137(.a(new_n229), .b(new_n230), .c(new_n225), .d(new_n232), .o1(\s[22] ));
  inv040aa1d32x5               g138(.a(\a[22] ), .o1(new_n234));
  xroi22aa1d06x4               g139(.a(new_n228), .b(\b[20] ), .c(new_n234), .d(\b[21] ), .out0(new_n235));
  and002aa1n02x5               g140(.a(new_n218), .b(new_n235), .o(new_n236));
  aob012aa1n02x5               g141(.a(new_n231), .b(\b[21] ), .c(\a[22] ), .out0(new_n237));
  oaib12aa1n02x5               g142(.a(new_n237), .b(\b[21] ), .c(new_n234), .out0(new_n238));
  tech160nm_fiao0012aa1n02p5x5 g143(.a(new_n238), .b(new_n223), .c(new_n235), .o(new_n239));
  xorc02aa1n02x5               g144(.a(\a[23] ), .b(\b[22] ), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n239), .c(new_n188), .d(new_n236), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(new_n240), .b(new_n238), .c(new_n223), .d(new_n235), .o1(new_n242));
  aobi12aa1n02x5               g147(.a(new_n242), .b(new_n188), .c(new_n236), .out0(new_n243));
  norb02aa1n02x5               g148(.a(new_n241), .b(new_n243), .out0(\s[23] ));
  inv000aa1d42x5               g149(.a(\a[23] ), .o1(new_n245));
  oaib12aa1n02x7               g150(.a(new_n241), .b(\b[22] ), .c(new_n245), .out0(new_n246));
  xorc02aa1n02x5               g151(.a(\a[24] ), .b(\b[23] ), .out0(new_n247));
  norp02aa1n02x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  norp02aa1n02x5               g153(.a(new_n247), .b(new_n248), .o1(new_n249));
  aoi022aa1n02x5               g154(.a(new_n246), .b(new_n247), .c(new_n241), .d(new_n249), .o1(\s[24] ));
  inv000aa1n02x5               g155(.a(new_n218), .o1(new_n251));
  inv000aa1d42x5               g156(.a(\a[24] ), .o1(new_n252));
  xroi22aa1d04x5               g157(.a(new_n245), .b(\b[22] ), .c(new_n252), .d(\b[23] ), .out0(new_n253));
  nano22aa1n02x4               g158(.a(new_n251), .b(new_n235), .c(new_n253), .out0(new_n254));
  nand02aa1d04x5               g159(.a(new_n188), .b(new_n254), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n253), .b(new_n238), .c(new_n223), .d(new_n235), .o1(new_n256));
  inv000aa1d42x5               g161(.a(\b[23] ), .o1(new_n257));
  oaoi03aa1n02x5               g162(.a(new_n252), .b(new_n257), .c(new_n248), .o1(new_n258));
  and002aa1n02x5               g163(.a(new_n256), .b(new_n258), .o(new_n259));
  xorc02aa1n12x5               g164(.a(\a[25] ), .b(\b[24] ), .out0(new_n260));
  aob012aa1n03x5               g165(.a(new_n260), .b(new_n255), .c(new_n259), .out0(new_n261));
  inv000aa1d42x5               g166(.a(new_n260), .o1(new_n262));
  and003aa1n02x5               g167(.a(new_n256), .b(new_n262), .c(new_n258), .o(new_n263));
  aobi12aa1n02x7               g168(.a(new_n261), .b(new_n263), .c(new_n255), .out0(\s[25] ));
  nor042aa1n03x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  aoai13aa1n02x5               g171(.a(new_n266), .b(new_n262), .c(new_n255), .d(new_n259), .o1(new_n267));
  xorc02aa1n02x5               g172(.a(\a[26] ), .b(\b[25] ), .out0(new_n268));
  norp02aa1n02x5               g173(.a(new_n268), .b(new_n265), .o1(new_n269));
  aoi022aa1n02x7               g174(.a(new_n267), .b(new_n268), .c(new_n261), .d(new_n269), .o1(\s[26] ));
  and002aa1n02x5               g175(.a(new_n268), .b(new_n260), .o(new_n271));
  aob012aa1n03x5               g176(.a(new_n271), .b(new_n256), .c(new_n258), .out0(new_n272));
  nano32aa1n02x5               g177(.a(new_n251), .b(new_n271), .c(new_n235), .d(new_n253), .out0(new_n273));
  nand02aa1d06x5               g178(.a(new_n188), .b(new_n273), .o1(new_n274));
  oao003aa1n02x5               g179(.a(\a[26] ), .b(\b[25] ), .c(new_n266), .carry(new_n275));
  nand23aa1n06x5               g180(.a(new_n272), .b(new_n274), .c(new_n275), .o1(new_n276));
  xorc02aa1n02x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n275), .o1(new_n278));
  aoi112aa1n02x5               g183(.a(new_n277), .b(new_n278), .c(new_n188), .d(new_n273), .o1(new_n279));
  aoi022aa1n02x5               g184(.a(new_n276), .b(new_n277), .c(new_n272), .d(new_n279), .o1(\s[27] ));
  nanp02aa1n03x5               g185(.a(new_n276), .b(new_n277), .o1(new_n281));
  tech160nm_fiaoi012aa1n05x5   g186(.a(new_n278), .b(new_n188), .c(new_n273), .o1(new_n282));
  orn002aa1n02x5               g187(.a(\a[27] ), .b(\b[26] ), .o(new_n283));
  and002aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .o(new_n284));
  aoai13aa1n03x5               g189(.a(new_n283), .b(new_n284), .c(new_n282), .d(new_n272), .o1(new_n285));
  norp02aa1n02x5               g190(.a(\b[27] ), .b(\a[28] ), .o1(new_n286));
  nanp02aa1n02x5               g191(.a(\b[27] ), .b(\a[28] ), .o1(new_n287));
  norb02aa1n02x5               g192(.a(new_n287), .b(new_n286), .out0(new_n288));
  norp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  aoib12aa1n02x5               g194(.a(new_n289), .b(new_n287), .c(new_n286), .out0(new_n290));
  aoi022aa1n03x5               g195(.a(new_n285), .b(new_n288), .c(new_n281), .d(new_n290), .o1(\s[28] ));
  nano23aa1n02x4               g196(.a(new_n286), .b(new_n284), .c(new_n283), .d(new_n287), .out0(new_n292));
  nand42aa1n02x5               g197(.a(new_n276), .b(new_n292), .o1(new_n293));
  inv000aa1n03x5               g198(.a(new_n292), .o1(new_n294));
  oai012aa1n02x5               g199(.a(new_n287), .b(new_n286), .c(new_n289), .o1(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n294), .c(new_n282), .d(new_n272), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[29] ), .b(\b[28] ), .out0(new_n297));
  norb02aa1n02x5               g202(.a(new_n295), .b(new_n297), .out0(new_n298));
  aoi022aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n293), .d(new_n298), .o1(\s[29] ));
  xorb03aa1n02x5               g204(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g205(.a(new_n277), .b(new_n297), .c(new_n288), .o(new_n301));
  nand22aa1n03x5               g206(.a(new_n276), .b(new_n301), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n301), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[29] ), .b(\b[28] ), .c(new_n295), .carry(new_n304));
  aoai13aa1n03x5               g209(.a(new_n304), .b(new_n303), .c(new_n282), .d(new_n272), .o1(new_n305));
  xorc02aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .out0(new_n306));
  norb02aa1n02x5               g211(.a(new_n304), .b(new_n306), .out0(new_n307));
  aoi022aa1n03x5               g212(.a(new_n305), .b(new_n306), .c(new_n302), .d(new_n307), .o1(\s[30] ));
  nano22aa1n02x4               g213(.a(new_n294), .b(new_n297), .c(new_n306), .out0(new_n309));
  nanp02aa1n03x5               g214(.a(new_n276), .b(new_n309), .o1(new_n310));
  xorc02aa1n02x5               g215(.a(\a[31] ), .b(\b[30] ), .out0(new_n311));
  and002aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .o(new_n312));
  oabi12aa1n02x5               g217(.a(new_n311), .b(\a[30] ), .c(\b[29] ), .out0(new_n313));
  oab012aa1n02x4               g218(.a(new_n313), .b(new_n304), .c(new_n312), .out0(new_n314));
  inv000aa1n02x5               g219(.a(new_n309), .o1(new_n315));
  oao003aa1n02x5               g220(.a(\a[30] ), .b(\b[29] ), .c(new_n304), .carry(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n315), .c(new_n282), .d(new_n272), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n311), .c(new_n310), .d(new_n314), .o1(\s[31] ));
  norp02aa1n02x5               g223(.a(new_n107), .b(new_n104), .o1(new_n319));
  oai012aa1n02x5               g224(.a(new_n103), .b(new_n106), .c(new_n105), .o1(new_n320));
  oaib12aa1n02x5               g225(.a(new_n320), .b(new_n102), .c(new_n101), .out0(new_n321));
  norb02aa1n02x5               g226(.a(new_n321), .b(new_n319), .out0(\s[3] ));
  obai22aa1n02x7               g227(.a(new_n113), .b(new_n108), .c(\a[3] ), .d(\b[2] ), .out0(new_n323));
  and002aa1n02x5               g228(.a(new_n110), .b(new_n113), .o(new_n324));
  inv000aa1d42x5               g229(.a(new_n324), .o1(new_n325));
  oa0022aa1n02x5               g230(.a(new_n325), .b(new_n108), .c(new_n319), .d(new_n323), .o(\s[4] ));
  nanb03aa1n02x5               g231(.a(new_n116), .b(new_n111), .c(new_n113), .out0(new_n327));
  oaoi13aa1n02x5               g232(.a(new_n327), .b(new_n109), .c(new_n107), .d(new_n104), .o1(new_n328));
  aboi22aa1n03x5               g233(.a(new_n116), .b(new_n111), .c(new_n110), .d(new_n113), .out0(new_n329));
  norp02aa1n02x5               g234(.a(new_n329), .b(new_n328), .o1(\s[5] ));
  xorc02aa1n02x5               g235(.a(\a[6] ), .b(\b[5] ), .out0(new_n331));
  oai012aa1n02x5               g236(.a(new_n331), .b(new_n328), .c(new_n116), .o1(new_n332));
  norp03aa1n02x5               g237(.a(new_n328), .b(new_n331), .c(new_n116), .o1(new_n333));
  norb02aa1n02x5               g238(.a(new_n332), .b(new_n333), .out0(\s[6] ));
  oai012aa1n02x5               g239(.a(new_n332), .b(\b[5] ), .c(\a[6] ), .o1(new_n335));
  xorb03aa1n02x5               g240(.a(new_n335), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp03aa1n02x5               g241(.a(new_n335), .b(new_n112), .c(new_n124), .o1(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n122), .b(new_n337), .c(new_n124), .out0(\s[8] ));
  xnbna2aa1n03x5               g243(.a(new_n131), .b(new_n121), .c(new_n128), .out0(\s[9] ));
endmodule


