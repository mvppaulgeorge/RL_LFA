// Benchmark "adder" written by ABC on Wed Jul 17 14:10:19 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n183, new_n184, new_n185, new_n186,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n320, new_n322, new_n323, new_n325, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[9] ), .o1(new_n97));
  nanb02aa1n12x5               g002(.a(\a[10] ), .b(new_n97), .out0(new_n98));
  nand42aa1n10x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  nanp02aa1n03x5               g004(.a(new_n98), .b(new_n99), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nand42aa1n03x5               g006(.a(\b[8] ), .b(\a[9] ), .o1(new_n102));
  nor002aa1n04x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  aoi022aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n104));
  nor002aa1n12x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand02aa1d16x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  norb02aa1n03x5               g011(.a(new_n106), .b(new_n105), .out0(new_n107));
  oai022aa1n09x5               g012(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n108));
  oaoi13aa1n04x5               g013(.a(new_n108), .b(new_n107), .c(new_n104), .d(new_n103), .o1(new_n109));
  nand42aa1n16x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  tech160nm_fioai012aa1n04x5   g015(.a(new_n110), .b(\b[7] ), .c(\a[8] ), .o1(new_n111));
  nor042aa1n09x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand42aa1n16x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  norb02aa1n03x5               g018(.a(new_n113), .b(new_n112), .out0(new_n114));
  nand42aa1d28x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  tech160nm_fioai012aa1n04x5   g020(.a(new_n115), .b(\b[5] ), .c(\a[6] ), .o1(new_n116));
  nand42aa1d28x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nand42aa1n08x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  nor042aa1n02x5               g023(.a(\b[4] ), .b(\a[5] ), .o1(new_n119));
  nano22aa1n03x7               g024(.a(new_n119), .b(new_n117), .c(new_n118), .out0(new_n120));
  nona23aa1n03x5               g025(.a(new_n120), .b(new_n114), .c(new_n111), .d(new_n116), .out0(new_n121));
  nano22aa1n03x7               g026(.a(new_n112), .b(new_n113), .c(new_n117), .out0(new_n122));
  oaih22aa1n04x5               g027(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n123));
  nor042aa1d18x5               g028(.a(\b[7] ), .b(\a[8] ), .o1(new_n124));
  norb02aa1n06x5               g029(.a(new_n115), .b(new_n124), .out0(new_n125));
  inv040aa1n02x5               g030(.a(new_n124), .o1(new_n126));
  aob012aa1n06x5               g031(.a(new_n126), .b(new_n112), .c(new_n115), .out0(new_n127));
  aoi013aa1n09x5               g032(.a(new_n127), .b(new_n122), .c(new_n123), .d(new_n125), .o1(new_n128));
  oai012aa1n06x5               g033(.a(new_n128), .b(new_n121), .c(new_n109), .o1(new_n129));
  aoai13aa1n02x5               g034(.a(new_n100), .b(new_n101), .c(new_n129), .d(new_n102), .o1(new_n130));
  oai112aa1n02x5               g035(.a(new_n98), .b(new_n99), .c(\b[8] ), .d(\a[9] ), .o1(new_n131));
  ao0012aa1n03x7               g036(.a(new_n131), .b(new_n129), .c(new_n102), .o(new_n132));
  nanp02aa1n02x5               g037(.a(new_n132), .b(new_n130), .o1(\s[10] ));
  nand02aa1n20x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n06x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n136), .b(new_n132), .c(new_n99), .out0(\s[11] ));
  inv040aa1n08x5               g042(.a(new_n135), .o1(new_n138));
  nanp03aa1n02x5               g043(.a(new_n132), .b(new_n99), .c(new_n136), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand02aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n12x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n139), .c(new_n138), .out0(\s[12] ));
  inv000aa1n06x5               g048(.a(new_n103), .o1(new_n144));
  nand42aa1n06x5               g049(.a(\b[0] ), .b(\a[1] ), .o1(new_n145));
  aob012aa1n12x5               g050(.a(new_n145), .b(\b[1] ), .c(\a[2] ), .out0(new_n146));
  nanb02aa1n06x5               g051(.a(new_n105), .b(new_n106), .out0(new_n147));
  inv000aa1n02x5               g052(.a(new_n108), .o1(new_n148));
  aoai13aa1n06x5               g053(.a(new_n148), .b(new_n147), .c(new_n146), .d(new_n144), .o1(new_n149));
  nanb02aa1n02x5               g054(.a(new_n112), .b(new_n113), .out0(new_n150));
  nor043aa1n02x5               g055(.a(new_n150), .b(new_n116), .c(new_n111), .o1(new_n151));
  nand03aa1n03x5               g056(.a(new_n149), .b(new_n151), .c(new_n120), .o1(new_n152));
  nano23aa1n02x4               g057(.a(new_n140), .b(new_n135), .c(new_n141), .d(new_n134), .out0(new_n153));
  nanb02aa1n03x5               g058(.a(new_n101), .b(new_n102), .out0(new_n154));
  nona22aa1n03x5               g059(.a(new_n153), .b(new_n154), .c(new_n100), .out0(new_n155));
  nor002aa1d32x5               g060(.a(\b[9] ), .b(\a[10] ), .o1(new_n156));
  oai112aa1n06x5               g061(.a(new_n138), .b(new_n99), .c(new_n101), .d(new_n156), .o1(new_n157));
  nanb03aa1n12x5               g062(.a(new_n140), .b(new_n141), .c(new_n134), .out0(new_n158));
  aoi012aa1d24x5               g063(.a(new_n140), .b(new_n135), .c(new_n141), .o1(new_n159));
  oai012aa1d24x5               g064(.a(new_n159), .b(new_n157), .c(new_n158), .o1(new_n160));
  inv000aa1d42x5               g065(.a(new_n160), .o1(new_n161));
  aoai13aa1n03x5               g066(.a(new_n161), .b(new_n155), .c(new_n152), .d(new_n128), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1d18x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n154), .b(new_n100), .c(new_n136), .d(new_n142), .out0(new_n166));
  nanp02aa1n04x5               g071(.a(\b[12] ), .b(\a[13] ), .o1(new_n167));
  norb02aa1n02x7               g072(.a(new_n167), .b(new_n164), .out0(new_n168));
  aoai13aa1n02x5               g073(.a(new_n168), .b(new_n160), .c(new_n129), .d(new_n166), .o1(new_n169));
  nor042aa1n04x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  nand22aa1n04x5               g075(.a(\b[13] ), .b(\a[14] ), .o1(new_n171));
  norb02aa1n06x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  xnbna2aa1n03x5               g077(.a(new_n172), .b(new_n169), .c(new_n165), .out0(\s[14] ));
  nano23aa1n06x5               g078(.a(new_n164), .b(new_n170), .c(new_n171), .d(new_n167), .out0(new_n174));
  aoi012aa1n12x5               g079(.a(new_n170), .b(new_n164), .c(new_n171), .o1(new_n175));
  inv000aa1n03x5               g080(.a(new_n175), .o1(new_n176));
  nor042aa1d18x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nand02aa1d06x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  norb02aa1n02x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  aoai13aa1n03x5               g084(.a(new_n179), .b(new_n176), .c(new_n162), .d(new_n174), .o1(new_n180));
  aoi112aa1n02x5               g085(.a(new_n179), .b(new_n176), .c(new_n162), .d(new_n174), .o1(new_n181));
  norb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(\s[15] ));
  inv040aa1n03x5               g087(.a(new_n177), .o1(new_n183));
  nor042aa1n06x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand22aa1n04x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  norb02aa1n02x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  xnbna2aa1n03x5               g091(.a(new_n186), .b(new_n180), .c(new_n183), .out0(\s[16] ));
  nona23aa1d18x5               g092(.a(new_n185), .b(new_n178), .c(new_n177), .d(new_n184), .out0(new_n188));
  nano22aa1n03x7               g093(.a(new_n188), .b(new_n168), .c(new_n172), .out0(new_n189));
  nand02aa1n02x5               g094(.a(new_n166), .b(new_n189), .o1(new_n190));
  oaoi03aa1n02x5               g095(.a(\a[16] ), .b(\b[15] ), .c(new_n183), .o1(new_n191));
  oabi12aa1n18x5               g096(.a(new_n191), .b(new_n188), .c(new_n175), .out0(new_n192));
  aoi012aa1n12x5               g097(.a(new_n192), .b(new_n160), .c(new_n189), .o1(new_n193));
  aoai13aa1n12x5               g098(.a(new_n193), .b(new_n190), .c(new_n152), .d(new_n128), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor022aa1n08x5               g100(.a(\b[16] ), .b(\a[17] ), .o1(new_n196));
  nand42aa1n16x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  tech160nm_fiaoi012aa1n05x5   g102(.a(new_n196), .b(new_n194), .c(new_n197), .o1(new_n198));
  xnrb03aa1n03x5               g103(.a(new_n198), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor042aa1n04x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nanp02aa1n04x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nano23aa1n09x5               g106(.a(new_n196), .b(new_n200), .c(new_n201), .d(new_n197), .out0(new_n202));
  aoi012aa1n02x5               g107(.a(new_n200), .b(new_n196), .c(new_n201), .o1(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  nor042aa1d18x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nand02aa1n04x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  norb02aa1n06x5               g111(.a(new_n206), .b(new_n205), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n204), .c(new_n194), .d(new_n202), .o1(new_n208));
  aoi112aa1n02x5               g113(.a(new_n207), .b(new_n204), .c(new_n194), .d(new_n202), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n208), .b(new_n209), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g116(.a(new_n205), .o1(new_n212));
  nor042aa1n04x5               g117(.a(\b[19] ), .b(\a[20] ), .o1(new_n213));
  nand02aa1d10x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  norb02aa1n06x5               g119(.a(new_n214), .b(new_n213), .out0(new_n215));
  xnbna2aa1n03x5               g120(.a(new_n215), .b(new_n208), .c(new_n212), .out0(\s[20] ));
  nano23aa1n02x5               g121(.a(new_n205), .b(new_n213), .c(new_n214), .d(new_n206), .out0(new_n217));
  nand02aa1d04x5               g122(.a(new_n217), .b(new_n202), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n218), .o1(new_n219));
  aoi112aa1n09x5               g124(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n220));
  oai112aa1n03x5               g125(.a(new_n207), .b(new_n215), .c(new_n220), .d(new_n200), .o1(new_n221));
  aoi012aa1n02x7               g126(.a(new_n213), .b(new_n205), .c(new_n214), .o1(new_n222));
  nanp02aa1n02x5               g127(.a(new_n221), .b(new_n222), .o1(new_n223));
  tech160nm_fiaoi012aa1n05x5   g128(.a(new_n223), .b(new_n194), .c(new_n219), .o1(new_n224));
  nor042aa1d18x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  inv040aa1n02x5               g130(.a(new_n225), .o1(new_n226));
  nanp02aa1n09x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  xnbna2aa1n03x5               g132(.a(new_n224), .b(new_n227), .c(new_n226), .out0(\s[21] ));
  norb02aa1n03x5               g133(.a(new_n227), .b(new_n225), .out0(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n223), .c(new_n194), .d(new_n219), .o1(new_n230));
  xnrc02aa1n12x5               g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  xobna2aa1n03x5               g136(.a(new_n231), .b(new_n230), .c(new_n226), .out0(\s[22] ));
  nano22aa1n03x7               g137(.a(new_n231), .b(new_n226), .c(new_n227), .out0(new_n233));
  nanb02aa1n02x5               g138(.a(new_n231), .b(new_n229), .out0(new_n234));
  oao003aa1n02x5               g139(.a(\a[22] ), .b(\b[21] ), .c(new_n226), .carry(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n234), .c(new_n221), .d(new_n222), .o1(new_n236));
  aoi013aa1n06x4               g141(.a(new_n236), .b(new_n194), .c(new_n219), .d(new_n233), .o1(new_n237));
  xnrb03aa1n03x5               g142(.a(new_n237), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g143(.a(\b[22] ), .b(\a[23] ), .o1(new_n239));
  inv000aa1d42x5               g144(.a(new_n239), .o1(new_n240));
  tech160nm_fixnrc02aa1n04x5   g145(.a(\b[22] ), .b(\a[23] ), .out0(new_n241));
  tech160nm_fixnrc02aa1n02p5x5 g146(.a(\b[23] ), .b(\a[24] ), .out0(new_n242));
  oaoi13aa1n03x5               g147(.a(new_n242), .b(new_n240), .c(new_n237), .d(new_n241), .o1(new_n243));
  nor042aa1n04x5               g148(.a(new_n237), .b(new_n241), .o1(new_n244));
  nano22aa1n03x7               g149(.a(new_n244), .b(new_n240), .c(new_n242), .out0(new_n245));
  norp02aa1n03x5               g150(.a(new_n243), .b(new_n245), .o1(\s[24] ));
  nor042aa1n02x5               g151(.a(new_n242), .b(new_n241), .o1(new_n247));
  oaoi03aa1n02x5               g152(.a(\a[24] ), .b(\b[23] ), .c(new_n240), .o1(new_n248));
  tech160nm_fiao0012aa1n02p5x5 g153(.a(new_n248), .b(new_n236), .c(new_n247), .o(new_n249));
  norb02aa1n02x5               g154(.a(new_n247), .b(new_n234), .out0(new_n250));
  aoi013aa1n06x4               g155(.a(new_n249), .b(new_n194), .c(new_n219), .d(new_n250), .o1(new_n251));
  xnrb03aa1n03x5               g156(.a(new_n251), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g157(.a(\b[24] ), .b(\a[25] ), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  tech160nm_fixnrc02aa1n05x5   g159(.a(\b[24] ), .b(\a[25] ), .out0(new_n255));
  xnrc02aa1n02x5               g160(.a(\b[25] ), .b(\a[26] ), .out0(new_n256));
  oaoi13aa1n02x5               g161(.a(new_n256), .b(new_n254), .c(new_n251), .d(new_n255), .o1(new_n257));
  norp02aa1n03x5               g162(.a(new_n251), .b(new_n255), .o1(new_n258));
  nano22aa1n03x5               g163(.a(new_n258), .b(new_n254), .c(new_n256), .out0(new_n259));
  norp02aa1n03x5               g164(.a(new_n257), .b(new_n259), .o1(\s[26] ));
  norp02aa1n02x5               g165(.a(new_n256), .b(new_n255), .o1(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n248), .c(new_n236), .d(new_n247), .o1(new_n262));
  nano23aa1n03x7               g167(.a(new_n177), .b(new_n184), .c(new_n185), .d(new_n178), .out0(new_n263));
  nanp02aa1n02x5               g168(.a(new_n263), .b(new_n174), .o1(new_n264));
  nor042aa1n02x5               g169(.a(new_n155), .b(new_n264), .o1(new_n265));
  aoi012aa1n02x5               g170(.a(new_n135), .b(\a[10] ), .c(\b[9] ), .o1(new_n266));
  nano22aa1n02x4               g171(.a(new_n140), .b(new_n134), .c(new_n141), .out0(new_n267));
  nanp03aa1n02x5               g172(.a(new_n267), .b(new_n131), .c(new_n266), .o1(new_n268));
  aoi012aa1n02x7               g173(.a(new_n191), .b(new_n263), .c(new_n176), .o1(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n264), .c(new_n268), .d(new_n159), .o1(new_n270));
  nano32aa1n03x7               g175(.a(new_n218), .b(new_n261), .c(new_n233), .d(new_n247), .out0(new_n271));
  aoai13aa1n06x5               g176(.a(new_n271), .b(new_n270), .c(new_n129), .d(new_n265), .o1(new_n272));
  oao003aa1n03x5               g177(.a(\a[26] ), .b(\b[25] ), .c(new_n254), .carry(new_n273));
  nanp03aa1d12x5               g178(.a(new_n262), .b(new_n272), .c(new_n273), .o1(new_n274));
  xorb03aa1n03x5               g179(.a(new_n274), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  inv000aa1n06x5               g181(.a(new_n276), .o1(new_n277));
  nanp02aa1n02x5               g182(.a(\b[26] ), .b(\a[27] ), .o1(new_n278));
  nand42aa1n08x5               g183(.a(new_n274), .b(new_n278), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[28] ), .b(\b[27] ), .out0(new_n280));
  inv000aa1n02x5               g185(.a(new_n280), .o1(new_n281));
  aoi012aa1n03x5               g186(.a(new_n281), .b(new_n279), .c(new_n277), .o1(new_n282));
  aoi112aa1n03x5               g187(.a(new_n276), .b(new_n280), .c(new_n274), .d(new_n278), .o1(new_n283));
  norp02aa1n03x5               g188(.a(new_n282), .b(new_n283), .o1(\s[28] ));
  nano22aa1n02x4               g189(.a(new_n281), .b(new_n277), .c(new_n278), .out0(new_n285));
  tech160nm_finand02aa1n03p5x5 g190(.a(new_n274), .b(new_n285), .o1(new_n286));
  oao003aa1n12x5               g191(.a(\a[28] ), .b(\b[27] ), .c(new_n277), .carry(new_n287));
  tech160nm_fixorc02aa1n03p5x5 g192(.a(\a[29] ), .b(\b[28] ), .out0(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  aoi012aa1n03x5               g194(.a(new_n289), .b(new_n286), .c(new_n287), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n287), .o1(new_n291));
  aoi112aa1n03x5               g196(.a(new_n288), .b(new_n291), .c(new_n274), .d(new_n285), .o1(new_n292));
  norp02aa1n03x5               g197(.a(new_n290), .b(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n145), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g199(.a(new_n289), .b(new_n280), .c(new_n278), .d(new_n277), .out0(new_n295));
  tech160nm_finand02aa1n03p5x5 g200(.a(new_n274), .b(new_n295), .o1(new_n296));
  oao003aa1n12x5               g201(.a(\a[29] ), .b(\b[28] ), .c(new_n287), .carry(new_n297));
  xorc02aa1n12x5               g202(.a(\a[30] ), .b(\b[29] ), .out0(new_n298));
  inv000aa1d42x5               g203(.a(new_n298), .o1(new_n299));
  aoi012aa1n03x5               g204(.a(new_n299), .b(new_n296), .c(new_n297), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n297), .o1(new_n301));
  aoi112aa1n03x5               g206(.a(new_n298), .b(new_n301), .c(new_n274), .d(new_n295), .o1(new_n302));
  norp02aa1n03x5               g207(.a(new_n300), .b(new_n302), .o1(\s[30] ));
  xnrc02aa1n02x5               g208(.a(\b[30] ), .b(\a[31] ), .out0(new_n304));
  and003aa1n03x7               g209(.a(new_n285), .b(new_n298), .c(new_n288), .o(new_n305));
  tech160nm_finand02aa1n03p5x5 g210(.a(new_n274), .b(new_n305), .o1(new_n306));
  tech160nm_fioaoi03aa1n03p5x5 g211(.a(\a[30] ), .b(\b[29] ), .c(new_n297), .o1(new_n307));
  inv000aa1n02x5               g212(.a(new_n307), .o1(new_n308));
  aoi012aa1n03x5               g213(.a(new_n304), .b(new_n306), .c(new_n308), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n304), .o1(new_n310));
  aoi112aa1n03x5               g215(.a(new_n310), .b(new_n307), .c(new_n274), .d(new_n305), .o1(new_n311));
  nor042aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[31] ));
  xnbna2aa1n03x5               g217(.a(new_n107), .b(new_n146), .c(new_n144), .out0(\s[3] ));
  inv000aa1d42x5               g218(.a(\a[4] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(\b[3] ), .o1(new_n315));
  nanp02aa1n02x5               g220(.a(new_n315), .b(new_n314), .o1(new_n316));
  aoi012aa1n02x5               g221(.a(new_n147), .b(new_n146), .c(new_n144), .o1(new_n317));
  aoi112aa1n02x5               g222(.a(new_n317), .b(new_n105), .c(new_n316), .d(new_n110), .o1(new_n318));
  aoi013aa1n02x4               g223(.a(new_n318), .b(new_n149), .c(new_n110), .d(new_n316), .o1(\s[4] ));
  nanb02aa1n02x5               g224(.a(new_n119), .b(new_n118), .out0(new_n320));
  xnbna2aa1n03x5               g225(.a(new_n320), .b(new_n149), .c(new_n110), .out0(\s[5] ));
  xorc02aa1n02x5               g226(.a(\a[6] ), .b(\b[5] ), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n118), .b(new_n119), .c(new_n149), .d(new_n110), .o1(new_n323));
  xnrc02aa1n02x5               g228(.a(new_n323), .b(new_n322), .out0(\s[6] ));
  aobi12aa1n02x5               g229(.a(new_n122), .b(new_n323), .c(new_n322), .out0(new_n325));
  oaoi03aa1n02x5               g230(.a(\a[6] ), .b(\b[5] ), .c(new_n323), .o1(new_n326));
  oab012aa1n02x4               g231(.a(new_n325), .b(new_n326), .c(new_n114), .out0(\s[7] ));
  norp02aa1n02x5               g232(.a(new_n325), .b(new_n112), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n328), .b(new_n126), .c(new_n115), .out0(\s[8] ));
  xorb03aa1n02x5               g234(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


