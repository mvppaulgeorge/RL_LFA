// Benchmark "adder" written by ABC on Wed Jul 17 14:10:56 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n283, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n303, new_n304, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n313, new_n315, new_n316, new_n318;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1d28x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  norp02aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[8] ), .b(\a[9] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  aoi022aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n103));
  nor002aa1n03x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  norb02aa1n03x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  oai022aa1n02x5               g011(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n107));
  oaoi13aa1n06x5               g012(.a(new_n107), .b(new_n106), .c(new_n103), .d(new_n102), .o1(new_n108));
  nanp02aa1n04x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  nand42aa1n02x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  norp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nano22aa1n02x4               g016(.a(new_n111), .b(new_n109), .c(new_n110), .out0(new_n112));
  xorc02aa1n02x5               g017(.a(\a[5] ), .b(\b[4] ), .out0(new_n113));
  nor042aa1n02x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand02aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  inv000aa1n02x5               g020(.a(new_n115), .o1(new_n116));
  nand22aa1n04x5               g021(.a(\b[3] ), .b(\a[4] ), .o1(new_n117));
  oai012aa1n02x5               g022(.a(new_n117), .b(\b[7] ), .c(\a[8] ), .o1(new_n118));
  nor003aa1n02x5               g023(.a(new_n118), .b(new_n116), .c(new_n114), .o1(new_n119));
  nanp03aa1n02x5               g024(.a(new_n119), .b(new_n112), .c(new_n113), .o1(new_n120));
  nano22aa1n02x5               g025(.a(new_n114), .b(new_n109), .c(new_n115), .out0(new_n121));
  oai022aa1n02x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  nor002aa1n02x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  norb02aa1n03x4               g028(.a(new_n110), .b(new_n123), .out0(new_n124));
  tech160nm_fiao0012aa1n02p5x5 g029(.a(new_n123), .b(new_n114), .c(new_n110), .o(new_n125));
  aoi013aa1n03x5               g030(.a(new_n125), .b(new_n121), .c(new_n122), .d(new_n124), .o1(new_n126));
  oai012aa1n12x5               g031(.a(new_n126), .b(new_n120), .c(new_n108), .o1(new_n127));
  aoai13aa1n02x5               g032(.a(new_n99), .b(new_n100), .c(new_n127), .d(new_n101), .o1(new_n128));
  inv040aa1n09x5               g033(.a(new_n97), .o1(new_n129));
  oai112aa1n06x5               g034(.a(new_n129), .b(new_n98), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  inv000aa1d42x5               g035(.a(new_n130), .o1(new_n131));
  aob012aa1n02x5               g036(.a(new_n131), .b(new_n127), .c(new_n101), .out0(new_n132));
  nanp02aa1n02x5               g037(.a(new_n128), .b(new_n132), .o1(\s[10] ));
  nand42aa1n03x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nor002aa1n02x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n136), .b(new_n132), .c(new_n98), .out0(\s[11] ));
  norp02aa1n02x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand42aa1n03x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n06x4               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoi013aa1n02x4               g045(.a(new_n135), .b(new_n132), .c(new_n134), .d(new_n98), .o1(new_n141));
  xnrc02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(\s[12] ));
  norb02aa1n02x5               g047(.a(new_n101), .b(new_n100), .out0(new_n143));
  nano32aa1n02x4               g048(.a(new_n99), .b(new_n143), .c(new_n136), .d(new_n140), .out0(new_n144));
  nanp02aa1n02x5               g049(.a(new_n127), .b(new_n144), .o1(new_n145));
  nano22aa1n02x4               g050(.a(new_n135), .b(new_n98), .c(new_n134), .out0(new_n146));
  nand43aa1n04x5               g051(.a(new_n130), .b(new_n146), .c(new_n140), .o1(new_n147));
  aoi012aa1n02x7               g052(.a(new_n138), .b(new_n135), .c(new_n139), .o1(new_n148));
  nanp02aa1n09x5               g053(.a(new_n147), .b(new_n148), .o1(new_n149));
  inv000aa1d42x5               g054(.a(new_n149), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(new_n145), .b(new_n150), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n04x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  aoi012aa1n02x5               g059(.a(new_n153), .b(new_n151), .c(new_n154), .o1(new_n155));
  xnrb03aa1n02x5               g060(.a(new_n155), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n03x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  nand22aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nano23aa1n06x5               g063(.a(new_n153), .b(new_n157), .c(new_n158), .d(new_n154), .out0(new_n159));
  aoai13aa1n06x5               g064(.a(new_n159), .b(new_n149), .c(new_n127), .d(new_n144), .o1(new_n160));
  aoi012aa1d18x5               g065(.a(new_n157), .b(new_n153), .c(new_n158), .o1(new_n161));
  nor002aa1n12x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  nanp02aa1n02x5               g067(.a(\b[14] ), .b(\a[15] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n160), .c(new_n161), .out0(\s[15] ));
  inv000aa1d42x5               g070(.a(new_n162), .o1(new_n166));
  inv000aa1d42x5               g071(.a(new_n164), .o1(new_n167));
  aoai13aa1n03x5               g072(.a(new_n166), .b(new_n167), .c(new_n160), .d(new_n161), .o1(new_n168));
  xorb03aa1n02x5               g073(.a(new_n168), .b(\b[15] ), .c(\a[16] ), .out0(\s[16] ));
  inv000aa1d42x5               g074(.a(\a[17] ), .o1(new_n170));
  nano23aa1n02x4               g075(.a(new_n135), .b(new_n97), .c(new_n98), .d(new_n134), .out0(new_n171));
  nor042aa1n02x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nano23aa1n09x5               g078(.a(new_n162), .b(new_n172), .c(new_n173), .d(new_n163), .out0(new_n174));
  nand02aa1d06x5               g079(.a(new_n174), .b(new_n159), .o1(new_n175));
  nano32aa1d12x5               g080(.a(new_n175), .b(new_n171), .c(new_n143), .d(new_n140), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n161), .o1(new_n177));
  oaoi03aa1n02x5               g082(.a(\a[16] ), .b(\b[15] ), .c(new_n166), .o1(new_n178));
  tech160nm_fiaoi012aa1n03p5x5 g083(.a(new_n178), .b(new_n174), .c(new_n177), .o1(new_n179));
  aoai13aa1n06x5               g084(.a(new_n179), .b(new_n175), .c(new_n147), .d(new_n148), .o1(new_n180));
  aoi012aa1n06x5               g085(.a(new_n180), .b(new_n127), .c(new_n176), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[16] ), .c(new_n170), .out0(\s[17] ));
  oaoi03aa1n02x5               g087(.a(\a[17] ), .b(\b[16] ), .c(new_n181), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nanp02aa1n02x5               g089(.a(new_n127), .b(new_n176), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n175), .o1(new_n186));
  aobi12aa1n06x5               g091(.a(new_n179), .b(new_n149), .c(new_n186), .out0(new_n187));
  nanp02aa1n06x5               g092(.a(new_n185), .b(new_n187), .o1(new_n188));
  inv000aa1d42x5               g093(.a(\a[18] ), .o1(new_n189));
  xroi22aa1d04x5               g094(.a(new_n170), .b(\b[16] ), .c(new_n189), .d(\b[17] ), .out0(new_n190));
  aoi112aa1n09x5               g095(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n191));
  oabi12aa1n02x5               g096(.a(new_n191), .b(\a[18] ), .c(\b[17] ), .out0(new_n192));
  nor042aa1d18x5               g097(.a(\b[18] ), .b(\a[19] ), .o1(new_n193));
  nand22aa1n12x5               g098(.a(\b[18] ), .b(\a[19] ), .o1(new_n194));
  norb02aa1n06x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  aoai13aa1n06x5               g100(.a(new_n195), .b(new_n192), .c(new_n188), .d(new_n190), .o1(new_n196));
  aoi112aa1n02x5               g101(.a(new_n195), .b(new_n192), .c(new_n188), .d(new_n190), .o1(new_n197));
  norb02aa1n02x5               g102(.a(new_n196), .b(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g103(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g104(.a(new_n193), .o1(new_n200));
  nor042aa1n06x5               g105(.a(\b[19] ), .b(\a[20] ), .o1(new_n201));
  nand22aa1n12x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  norb02aa1n06x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  aobi12aa1n03x5               g108(.a(new_n203), .b(new_n196), .c(new_n200), .out0(new_n204));
  nona22aa1n03x5               g109(.a(new_n196), .b(new_n203), .c(new_n193), .out0(new_n205));
  norb02aa1n03x4               g110(.a(new_n205), .b(new_n204), .out0(\s[20] ));
  nano23aa1n02x5               g111(.a(new_n193), .b(new_n201), .c(new_n202), .d(new_n194), .out0(new_n207));
  nand02aa1d04x5               g112(.a(new_n190), .b(new_n207), .o1(new_n208));
  inv000aa1d42x5               g113(.a(new_n208), .o1(new_n209));
  aoai13aa1n06x5               g114(.a(new_n209), .b(new_n180), .c(new_n127), .d(new_n176), .o1(new_n210));
  tech160nm_fiaoi012aa1n03p5x5 g115(.a(new_n201), .b(new_n193), .c(new_n202), .o1(new_n211));
  aobi12aa1n02x5               g116(.a(new_n211), .b(new_n192), .c(new_n207), .out0(new_n212));
  xorc02aa1n12x5               g117(.a(\a[21] ), .b(\b[20] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n210), .c(new_n212), .out0(\s[21] ));
  norp02aa1n02x5               g119(.a(\b[20] ), .b(\a[21] ), .o1(new_n215));
  aobi12aa1n06x5               g120(.a(new_n213), .b(new_n210), .c(new_n212), .out0(new_n216));
  xnrc02aa1n12x5               g121(.a(\b[21] ), .b(\a[22] ), .out0(new_n217));
  oab012aa1n03x5               g122(.a(new_n217), .b(new_n216), .c(new_n215), .out0(new_n218));
  norb03aa1n02x5               g123(.a(new_n217), .b(new_n216), .c(new_n215), .out0(new_n219));
  norp02aa1n02x5               g124(.a(new_n218), .b(new_n219), .o1(\s[22] ));
  nanb02aa1n06x5               g125(.a(new_n217), .b(new_n213), .out0(new_n221));
  nor042aa1n02x5               g126(.a(\b[17] ), .b(\a[18] ), .o1(new_n222));
  oai112aa1n06x5               g127(.a(new_n195), .b(new_n203), .c(new_n191), .d(new_n222), .o1(new_n223));
  aoi112aa1n02x5               g128(.a(\b[20] ), .b(\a[21] ), .c(\a[22] ), .d(\b[21] ), .o1(new_n224));
  oab012aa1n04x5               g129(.a(new_n224), .b(\a[22] ), .c(\b[21] ), .out0(new_n225));
  aoai13aa1n12x5               g130(.a(new_n225), .b(new_n221), .c(new_n223), .d(new_n211), .o1(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[22] ), .b(\a[23] ), .out0(new_n228));
  oaoi13aa1n09x5               g133(.a(new_n228), .b(new_n227), .c(new_n210), .d(new_n221), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n213), .b(new_n217), .out0(new_n230));
  nano22aa1n03x7               g135(.a(new_n181), .b(new_n209), .c(new_n230), .out0(new_n231));
  nano22aa1n02x4               g136(.a(new_n231), .b(new_n227), .c(new_n228), .out0(new_n232));
  norp02aa1n02x5               g137(.a(new_n229), .b(new_n232), .o1(\s[23] ));
  nor042aa1n06x5               g138(.a(\b[22] ), .b(\a[23] ), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  oabi12aa1n02x5               g140(.a(new_n228), .b(new_n231), .c(new_n226), .out0(new_n236));
  tech160nm_fixnrc02aa1n04x5   g141(.a(\b[23] ), .b(\a[24] ), .out0(new_n237));
  aoi012aa1n03x5               g142(.a(new_n237), .b(new_n236), .c(new_n235), .o1(new_n238));
  nano22aa1n02x4               g143(.a(new_n229), .b(new_n235), .c(new_n237), .out0(new_n239));
  norp02aa1n02x5               g144(.a(new_n238), .b(new_n239), .o1(\s[24] ));
  nor042aa1n04x5               g145(.a(new_n237), .b(new_n228), .o1(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[24] ), .b(\b[23] ), .c(new_n235), .o1(new_n242));
  aoi012aa1d18x5               g147(.a(new_n242), .b(new_n226), .c(new_n241), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n241), .o1(new_n244));
  nona32aa1n06x5               g149(.a(new_n188), .b(new_n244), .c(new_n221), .d(new_n208), .out0(new_n245));
  xnrc02aa1n03x5               g150(.a(\b[24] ), .b(\a[25] ), .out0(new_n246));
  xobna2aa1n03x5               g151(.a(new_n246), .b(new_n245), .c(new_n243), .out0(\s[25] ));
  nor042aa1n03x5               g152(.a(\b[24] ), .b(\a[25] ), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n248), .o1(new_n249));
  inv000aa1d42x5               g154(.a(new_n243), .o1(new_n250));
  nano32aa1n03x7               g155(.a(new_n181), .b(new_n241), .c(new_n209), .d(new_n230), .out0(new_n251));
  oabi12aa1n02x7               g156(.a(new_n246), .b(new_n251), .c(new_n250), .out0(new_n252));
  xnrc02aa1n02x5               g157(.a(\b[25] ), .b(\a[26] ), .out0(new_n253));
  tech160nm_fiaoi012aa1n04x5   g158(.a(new_n253), .b(new_n252), .c(new_n249), .o1(new_n254));
  tech160nm_fiaoi012aa1n05x5   g159(.a(new_n246), .b(new_n245), .c(new_n243), .o1(new_n255));
  nano22aa1n03x5               g160(.a(new_n255), .b(new_n249), .c(new_n253), .out0(new_n256));
  norp02aa1n03x5               g161(.a(new_n254), .b(new_n256), .o1(\s[26] ));
  norp02aa1n02x5               g162(.a(new_n253), .b(new_n246), .o1(new_n258));
  nano32aa1n06x5               g163(.a(new_n208), .b(new_n258), .c(new_n230), .d(new_n241), .out0(new_n259));
  aoai13aa1n06x5               g164(.a(new_n259), .b(new_n180), .c(new_n127), .d(new_n176), .o1(new_n260));
  aoai13aa1n09x5               g165(.a(new_n258), .b(new_n242), .c(new_n226), .d(new_n241), .o1(new_n261));
  oao003aa1n02x5               g166(.a(\a[26] ), .b(\b[25] ), .c(new_n249), .carry(new_n262));
  nanp03aa1d12x5               g167(.a(new_n260), .b(new_n261), .c(new_n262), .o1(new_n263));
  xorb03aa1n03x5               g168(.a(new_n263), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1d18x5               g169(.a(\b[26] ), .b(\a[27] ), .o1(new_n265));
  inv040aa1n08x5               g170(.a(new_n265), .o1(new_n266));
  nanp02aa1n02x5               g171(.a(\b[26] ), .b(\a[27] ), .o1(new_n267));
  nanp02aa1n03x5               g172(.a(new_n263), .b(new_n267), .o1(new_n268));
  xorc02aa1n12x5               g173(.a(\a[28] ), .b(\b[27] ), .out0(new_n269));
  inv000aa1d42x5               g174(.a(new_n269), .o1(new_n270));
  aoi012aa1n03x5               g175(.a(new_n270), .b(new_n268), .c(new_n266), .o1(new_n271));
  aoi112aa1n03x4               g176(.a(new_n265), .b(new_n269), .c(new_n263), .d(new_n267), .o1(new_n272));
  norp02aa1n03x5               g177(.a(new_n271), .b(new_n272), .o1(\s[28] ));
  nano22aa1n02x4               g178(.a(new_n270), .b(new_n266), .c(new_n267), .out0(new_n274));
  nanp02aa1n03x5               g179(.a(new_n263), .b(new_n274), .o1(new_n275));
  oao003aa1n12x5               g180(.a(\a[28] ), .b(\b[27] ), .c(new_n266), .carry(new_n276));
  tech160nm_fixorc02aa1n02p5x5 g181(.a(\a[29] ), .b(\b[28] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  aoi012aa1n03x5               g183(.a(new_n278), .b(new_n275), .c(new_n276), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n276), .o1(new_n280));
  aoi112aa1n03x4               g185(.a(new_n277), .b(new_n280), .c(new_n263), .d(new_n274), .o1(new_n281));
  norp02aa1n03x5               g186(.a(new_n279), .b(new_n281), .o1(\s[29] ));
  nanp02aa1n02x5               g187(.a(\b[0] ), .b(\a[1] ), .o1(new_n283));
  xorb03aa1n02x5               g188(.a(new_n283), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g189(.a(new_n278), .b(new_n269), .c(new_n267), .d(new_n266), .out0(new_n285));
  nand42aa1n02x5               g190(.a(new_n263), .b(new_n285), .o1(new_n286));
  oao003aa1n12x5               g191(.a(\a[29] ), .b(\b[28] ), .c(new_n276), .carry(new_n287));
  tech160nm_fixorc02aa1n02p5x5 g192(.a(\a[30] ), .b(\b[29] ), .out0(new_n288));
  inv000aa1d42x5               g193(.a(new_n288), .o1(new_n289));
  aoi012aa1n03x5               g194(.a(new_n289), .b(new_n286), .c(new_n287), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n287), .o1(new_n291));
  aoi112aa1n03x4               g196(.a(new_n288), .b(new_n291), .c(new_n263), .d(new_n285), .o1(new_n292));
  norp02aa1n03x5               g197(.a(new_n290), .b(new_n292), .o1(\s[30] ));
  xnrc02aa1n02x5               g198(.a(\b[30] ), .b(\a[31] ), .out0(new_n294));
  and003aa1n03x7               g199(.a(new_n274), .b(new_n288), .c(new_n277), .o(new_n295));
  nanp02aa1n03x5               g200(.a(new_n263), .b(new_n295), .o1(new_n296));
  oaoi03aa1n12x5               g201(.a(\a[30] ), .b(\b[29] ), .c(new_n287), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n297), .o1(new_n298));
  aoi012aa1n03x5               g203(.a(new_n294), .b(new_n296), .c(new_n298), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n294), .o1(new_n300));
  aoi112aa1n03x5               g205(.a(new_n300), .b(new_n297), .c(new_n263), .d(new_n295), .o1(new_n301));
  nor042aa1n03x5               g206(.a(new_n299), .b(new_n301), .o1(\s[31] ));
  inv000aa1n02x5               g207(.a(new_n102), .o1(new_n303));
  aob012aa1n02x5               g208(.a(new_n283), .b(\b[1] ), .c(\a[2] ), .out0(new_n304));
  xnbna2aa1n03x5               g209(.a(new_n106), .b(new_n304), .c(new_n303), .out0(\s[3] ));
  norp02aa1n02x5               g210(.a(\b[3] ), .b(\a[4] ), .o1(new_n306));
  nanp02aa1n02x5               g211(.a(new_n304), .b(new_n303), .o1(new_n307));
  obai22aa1n02x7               g212(.a(new_n117), .b(new_n306), .c(\a[3] ), .d(\b[2] ), .out0(new_n308));
  aoi012aa1n02x5               g213(.a(new_n308), .b(new_n307), .c(new_n106), .o1(new_n309));
  aoai13aa1n02x5               g214(.a(new_n117), .b(new_n107), .c(new_n307), .d(new_n106), .o1(new_n310));
  oab012aa1n02x4               g215(.a(new_n309), .b(new_n310), .c(new_n306), .out0(\s[4] ));
  xnrc02aa1n02x5               g216(.a(new_n310), .b(new_n113), .out0(\s[5] ));
  oao003aa1n03x5               g217(.a(\a[5] ), .b(\b[4] ), .c(new_n310), .carry(new_n313));
  xnrb03aa1n02x5               g218(.a(new_n313), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g219(.a(new_n115), .b(new_n114), .out0(new_n315));
  nanb03aa1n02x5               g220(.a(new_n111), .b(new_n313), .c(new_n109), .out0(new_n316));
  xobna2aa1n03x5               g221(.a(new_n315), .b(new_n316), .c(new_n109), .out0(\s[7] ));
  tech160nm_fiaoi012aa1n05x5   g222(.a(new_n114), .b(new_n316), .c(new_n121), .o1(new_n318));
  xnrc02aa1n02x5               g223(.a(new_n318), .b(new_n124), .out0(\s[8] ));
  xorb03aa1n02x5               g224(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


