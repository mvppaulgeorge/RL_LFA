// Benchmark "adder" written by ABC on Thu Jul 18 05:01:55 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n311, new_n312, new_n313, new_n316, new_n317, new_n318, new_n320,
    new_n322, new_n323, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n04x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\a[3] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[4] ), .o1(new_n99));
  inv040aa1d32x5               g004(.a(\b[2] ), .o1(new_n100));
  aboi22aa1n12x5               g005(.a(\b[3] ), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n101));
  nand22aa1n12x5               g006(.a(new_n100), .b(new_n98), .o1(new_n102));
  nand22aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand02aa1d04x5               g008(.a(new_n102), .b(new_n103), .o1(new_n104));
  nor042aa1d18x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand02aa1d28x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nand42aa1n08x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  oai012aa1d24x5               g012(.a(new_n107), .b(new_n105), .c(new_n106), .o1(new_n108));
  oai012aa1n12x5               g013(.a(new_n101), .b(new_n108), .c(new_n104), .o1(new_n109));
  nand22aa1n12x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  orn002aa1n12x5               g015(.a(\a[6] ), .b(\b[5] ), .o(new_n111));
  nand42aa1n06x5               g016(.a(\b[3] ), .b(\a[4] ), .o1(new_n112));
  xnrc02aa1n12x5               g017(.a(\b[4] ), .b(\a[5] ), .out0(new_n113));
  nano32aa1n03x7               g018(.a(new_n113), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n114));
  nand42aa1d28x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nor022aa1n16x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nand42aa1n10x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  nano23aa1n09x5               g023(.a(new_n117), .b(new_n116), .c(new_n118), .d(new_n115), .out0(new_n119));
  nand03aa1n08x5               g024(.a(new_n109), .b(new_n114), .c(new_n119), .o1(new_n120));
  nona22aa1n09x5               g025(.a(new_n115), .b(new_n116), .c(new_n117), .out0(new_n121));
  nor002aa1d32x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  aob012aa1n06x5               g027(.a(new_n111), .b(new_n122), .c(new_n110), .out0(new_n123));
  aoi022aa1n12x5               g028(.a(new_n119), .b(new_n123), .c(new_n115), .d(new_n121), .o1(new_n124));
  oai112aa1n02x5               g029(.a(new_n120), .b(new_n124), .c(\b[8] ), .d(\a[9] ), .o1(new_n125));
  nor002aa1d32x5               g030(.a(\b[9] ), .b(\a[10] ), .o1(new_n126));
  nand02aa1n12x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n126), .b(new_n127), .out0(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n128), .b(new_n125), .c(new_n97), .out0(\s[10] ));
  nand02aa1d16x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor002aa1d32x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n127), .b(new_n126), .c(new_n125), .d(new_n97), .o1(new_n133));
  nano22aa1n02x4               g038(.a(new_n131), .b(new_n127), .c(new_n130), .out0(new_n134));
  aoai13aa1n02x5               g039(.a(new_n134), .b(new_n126), .c(new_n125), .d(new_n97), .o1(new_n135));
  aobi12aa1n02x5               g040(.a(new_n135), .b(new_n133), .c(new_n132), .out0(\s[11] ));
  inv000aa1d42x5               g041(.a(new_n131), .o1(new_n137));
  nor022aa1n16x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nand22aa1n06x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n135), .c(new_n137), .out0(\s[12] ));
  nona23aa1d18x5               g046(.a(new_n130), .b(new_n139), .c(new_n138), .d(new_n131), .out0(new_n142));
  norp02aa1n24x5               g047(.a(\b[8] ), .b(\a[9] ), .o1(new_n143));
  nona23aa1n09x5               g048(.a(new_n97), .b(new_n127), .c(new_n126), .d(new_n143), .out0(new_n144));
  nor042aa1d18x5               g049(.a(new_n144), .b(new_n142), .o1(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  oai112aa1n02x7               g051(.a(new_n127), .b(new_n130), .c(new_n126), .d(new_n143), .o1(new_n147));
  nona22aa1n03x5               g052(.a(new_n147), .b(new_n138), .c(new_n131), .out0(new_n148));
  and002aa1n18x5               g053(.a(new_n148), .b(new_n139), .o(new_n149));
  inv000aa1n06x5               g054(.a(new_n149), .o1(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n146), .c(new_n120), .d(new_n124), .o1(new_n151));
  nor002aa1d24x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  nand42aa1n08x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  norb02aa1n02x7               g058(.a(new_n153), .b(new_n152), .out0(new_n154));
  nanp02aa1n03x5               g059(.a(new_n120), .b(new_n124), .o1(new_n155));
  aoi112aa1n02x5               g060(.a(new_n154), .b(new_n149), .c(new_n155), .d(new_n145), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n156), .b(new_n151), .c(new_n154), .o1(\s[13] ));
  nor042aa1d18x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand22aa1n09x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  norb02aa1n03x5               g064(.a(new_n159), .b(new_n158), .out0(new_n160));
  aoi112aa1n02x5               g065(.a(new_n152), .b(new_n160), .c(new_n151), .d(new_n154), .o1(new_n161));
  aoai13aa1n02x5               g066(.a(new_n160), .b(new_n152), .c(new_n151), .d(new_n153), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(\s[14] ));
  nano23aa1n02x4               g068(.a(new_n152), .b(new_n158), .c(new_n159), .d(new_n153), .out0(new_n164));
  aoai13aa1n02x5               g069(.a(new_n164), .b(new_n149), .c(new_n155), .d(new_n145), .o1(new_n165));
  aoi012aa1d18x5               g070(.a(new_n158), .b(new_n152), .c(new_n159), .o1(new_n166));
  nor002aa1n20x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nand22aa1n03x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n165), .c(new_n166), .out0(\s[15] ));
  aob012aa1n02x5               g075(.a(new_n169), .b(new_n165), .c(new_n166), .out0(new_n171));
  nor002aa1d32x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nand02aa1d04x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  aoib12aa1n02x5               g079(.a(new_n167), .b(new_n173), .c(new_n172), .out0(new_n175));
  aobi12aa1n02x5               g080(.a(new_n166), .b(new_n151), .c(new_n164), .out0(new_n176));
  tech160nm_fioaoi03aa1n03p5x5 g081(.a(\a[15] ), .b(\b[14] ), .c(new_n176), .o1(new_n177));
  aoi022aa1n03x5               g082(.a(new_n177), .b(new_n174), .c(new_n171), .d(new_n175), .o1(\s[16] ));
  nona23aa1n09x5               g083(.a(new_n173), .b(new_n168), .c(new_n167), .d(new_n172), .out0(new_n179));
  nano22aa1n03x7               g084(.a(new_n179), .b(new_n154), .c(new_n160), .out0(new_n180));
  nand02aa1d04x5               g085(.a(new_n180), .b(new_n145), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n181), .b(new_n155), .out0(new_n182));
  aoi012aa1n02x7               g087(.a(new_n172), .b(\a[15] ), .c(\b[14] ), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n152), .b(\a[12] ), .c(\b[11] ), .o1(new_n184));
  nona23aa1n03x5               g089(.a(new_n159), .b(new_n153), .c(new_n167), .d(new_n158), .out0(new_n185));
  nano32aa1n03x7               g090(.a(new_n185), .b(new_n184), .c(new_n183), .d(new_n173), .out0(new_n186));
  tech160nm_fiaoi012aa1n03p5x5 g091(.a(new_n172), .b(new_n167), .c(new_n173), .o1(new_n187));
  oai012aa1n06x5               g092(.a(new_n187), .b(new_n179), .c(new_n166), .o1(new_n188));
  aoi012aa1n06x5               g093(.a(new_n188), .b(new_n186), .c(new_n148), .o1(new_n189));
  aoai13aa1n12x5               g094(.a(new_n189), .b(new_n181), .c(new_n120), .d(new_n124), .o1(new_n190));
  xorc02aa1n12x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  aoi112aa1n02x5               g096(.a(new_n188), .b(new_n191), .c(new_n186), .d(new_n148), .o1(new_n192));
  aoi022aa1n02x5               g097(.a(new_n192), .b(new_n182), .c(new_n190), .d(new_n191), .o1(\s[17] ));
  inv000aa1d42x5               g098(.a(\a[17] ), .o1(new_n194));
  nanb02aa1n02x5               g099(.a(\b[16] ), .b(new_n194), .out0(new_n195));
  nanp02aa1n02x5               g100(.a(new_n190), .b(new_n191), .o1(new_n196));
  xorc02aa1n12x5               g101(.a(\a[18] ), .b(\b[17] ), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n196), .c(new_n195), .out0(\s[18] ));
  and002aa1n06x5               g103(.a(new_n197), .b(new_n191), .o(new_n199));
  nor042aa1n02x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  aoi112aa1n09x5               g105(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n201));
  norp02aa1n02x5               g106(.a(new_n201), .b(new_n200), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  xorc02aa1n12x5               g108(.a(\a[19] ), .b(\b[18] ), .out0(new_n204));
  aoai13aa1n06x5               g109(.a(new_n204), .b(new_n203), .c(new_n190), .d(new_n199), .o1(new_n205));
  aoi112aa1n02x5               g110(.a(new_n204), .b(new_n203), .c(new_n190), .d(new_n199), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n205), .b(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n06x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand42aa1n16x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n12x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  orn002aa1n06x5               g116(.a(\a[19] ), .b(\b[18] ), .o(new_n212));
  norb02aa1n02x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  nanp02aa1n02x5               g118(.a(new_n205), .b(new_n212), .o1(new_n214));
  aoi022aa1n02x5               g119(.a(new_n214), .b(new_n211), .c(new_n205), .d(new_n213), .o1(\s[20] ));
  nand23aa1n03x5               g120(.a(new_n199), .b(new_n204), .c(new_n211), .o1(new_n216));
  nanb02aa1n06x5               g121(.a(new_n216), .b(new_n190), .out0(new_n217));
  oai112aa1n06x5               g122(.a(new_n204), .b(new_n211), .c(new_n201), .d(new_n200), .o1(new_n218));
  oaib12aa1n18x5               g123(.a(new_n210), .b(new_n209), .c(new_n212), .out0(new_n219));
  nanp02aa1n02x5               g124(.a(new_n218), .b(new_n219), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  xorc02aa1n12x5               g126(.a(\a[21] ), .b(\b[20] ), .out0(new_n222));
  xnbna2aa1n03x5               g127(.a(new_n222), .b(new_n217), .c(new_n221), .out0(\s[21] ));
  aob012aa1n03x5               g128(.a(new_n222), .b(new_n217), .c(new_n221), .out0(new_n224));
  tech160nm_fixorc02aa1n02p5x5 g129(.a(\a[22] ), .b(\b[21] ), .out0(new_n225));
  nor042aa1n06x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  norp02aa1n02x5               g131(.a(new_n225), .b(new_n226), .o1(new_n227));
  inv000aa1d42x5               g132(.a(new_n226), .o1(new_n228));
  and002aa1n02x5               g133(.a(\b[20] ), .b(\a[21] ), .o(new_n229));
  aoai13aa1n02x5               g134(.a(new_n228), .b(new_n229), .c(new_n217), .d(new_n221), .o1(new_n230));
  aoi022aa1n02x5               g135(.a(new_n230), .b(new_n225), .c(new_n224), .d(new_n227), .o1(\s[22] ));
  nand22aa1n03x5               g136(.a(new_n225), .b(new_n222), .o1(new_n232));
  nano32aa1n02x4               g137(.a(new_n232), .b(new_n199), .c(new_n204), .d(new_n211), .out0(new_n233));
  oao003aa1n03x5               g138(.a(\a[22] ), .b(\b[21] ), .c(new_n228), .carry(new_n234));
  aoai13aa1n12x5               g139(.a(new_n234), .b(new_n232), .c(new_n218), .d(new_n219), .o1(new_n235));
  xorc02aa1n12x5               g140(.a(\a[23] ), .b(\b[22] ), .out0(new_n236));
  aoai13aa1n06x5               g141(.a(new_n236), .b(new_n235), .c(new_n190), .d(new_n233), .o1(new_n237));
  aoi112aa1n02x5               g142(.a(new_n236), .b(new_n235), .c(new_n190), .d(new_n233), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n237), .b(new_n238), .out0(\s[23] ));
  tech160nm_fixorc02aa1n03p5x5 g144(.a(\a[24] ), .b(\b[23] ), .out0(new_n240));
  orn002aa1n02x5               g145(.a(\a[23] ), .b(\b[22] ), .o(new_n241));
  norb02aa1n02x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  nanp02aa1n02x5               g147(.a(new_n237), .b(new_n241), .o1(new_n243));
  aoi022aa1n02x5               g148(.a(new_n243), .b(new_n240), .c(new_n237), .d(new_n242), .o1(\s[24] ));
  and002aa1n06x5               g149(.a(new_n240), .b(new_n236), .o(new_n245));
  oaoi03aa1n02x5               g150(.a(\a[24] ), .b(\b[23] ), .c(new_n241), .o1(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(new_n235), .c(new_n245), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n245), .o1(new_n248));
  nona32aa1n06x5               g153(.a(new_n190), .b(new_n248), .c(new_n232), .d(new_n216), .out0(new_n249));
  xorc02aa1n12x5               g154(.a(\a[25] ), .b(\b[24] ), .out0(new_n250));
  xnbna2aa1n03x5               g155(.a(new_n250), .b(new_n249), .c(new_n247), .out0(\s[25] ));
  aob012aa1n03x5               g156(.a(new_n250), .b(new_n249), .c(new_n247), .out0(new_n252));
  xorc02aa1n02x5               g157(.a(\a[26] ), .b(\b[25] ), .out0(new_n253));
  orn002aa1n02x5               g158(.a(\a[25] ), .b(\b[24] ), .o(new_n254));
  norb02aa1n02x5               g159(.a(new_n254), .b(new_n253), .out0(new_n255));
  inv000aa1d42x5               g160(.a(new_n250), .o1(new_n256));
  aoai13aa1n03x5               g161(.a(new_n254), .b(new_n256), .c(new_n249), .d(new_n247), .o1(new_n257));
  aoi022aa1n03x5               g162(.a(new_n257), .b(new_n253), .c(new_n252), .d(new_n255), .o1(\s[26] ));
  and002aa1n06x5               g163(.a(new_n253), .b(new_n250), .o(new_n259));
  aoai13aa1n12x5               g164(.a(new_n259), .b(new_n246), .c(new_n235), .d(new_n245), .o1(new_n260));
  nano22aa1n02x4               g165(.a(new_n232), .b(new_n236), .c(new_n240), .out0(new_n261));
  nano22aa1n03x7               g166(.a(new_n216), .b(new_n261), .c(new_n259), .out0(new_n262));
  nanp02aa1n06x5               g167(.a(new_n190), .b(new_n262), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(\b[25] ), .b(\a[26] ), .o1(new_n264));
  oai022aa1n02x5               g169(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(new_n265), .b(new_n264), .o1(new_n266));
  nanp03aa1n09x5               g171(.a(new_n263), .b(new_n260), .c(new_n266), .o1(new_n267));
  xorc02aa1n12x5               g172(.a(\a[27] ), .b(\b[26] ), .out0(new_n268));
  aoi122aa1n02x5               g173(.a(new_n268), .b(new_n264), .c(new_n265), .d(new_n190), .e(new_n262), .o1(new_n269));
  aoi022aa1n02x5               g174(.a(new_n269), .b(new_n260), .c(new_n267), .d(new_n268), .o1(\s[27] ));
  nand02aa1n04x5               g175(.a(new_n267), .b(new_n268), .o1(new_n271));
  xorc02aa1n02x5               g176(.a(\a[28] ), .b(\b[27] ), .out0(new_n272));
  norp02aa1n02x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  norp02aa1n02x5               g178(.a(new_n272), .b(new_n273), .o1(new_n274));
  aoi022aa1n06x5               g179(.a(new_n190), .b(new_n262), .c(new_n264), .d(new_n265), .o1(new_n275));
  inv000aa1n06x5               g180(.a(new_n273), .o1(new_n276));
  inv000aa1d42x5               g181(.a(new_n268), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n276), .b(new_n277), .c(new_n275), .d(new_n260), .o1(new_n278));
  aoi022aa1n03x5               g183(.a(new_n278), .b(new_n272), .c(new_n271), .d(new_n274), .o1(\s[28] ));
  and002aa1n06x5               g184(.a(new_n272), .b(new_n268), .o(new_n280));
  nanp02aa1n03x5               g185(.a(new_n267), .b(new_n280), .o1(new_n281));
  tech160nm_fixorc02aa1n02p5x5 g186(.a(\a[29] ), .b(\b[28] ), .out0(new_n282));
  norp02aa1n02x5               g187(.a(\b[27] ), .b(\a[28] ), .o1(new_n283));
  aoi112aa1n02x5               g188(.a(\b[26] ), .b(\a[27] ), .c(\a[28] ), .d(\b[27] ), .o1(new_n284));
  norp03aa1n02x5               g189(.a(new_n282), .b(new_n284), .c(new_n283), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n280), .o1(new_n286));
  oaoi03aa1n12x5               g191(.a(\a[28] ), .b(\b[27] ), .c(new_n276), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n286), .c(new_n275), .d(new_n260), .o1(new_n289));
  aoi022aa1n03x5               g194(.a(new_n289), .b(new_n282), .c(new_n281), .d(new_n285), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g196(.a(new_n277), .b(new_n272), .c(new_n282), .out0(new_n292));
  nand42aa1n02x5               g197(.a(new_n267), .b(new_n292), .o1(new_n293));
  xorc02aa1n02x5               g198(.a(\a[30] ), .b(\b[29] ), .out0(new_n294));
  inv000aa1d42x5               g199(.a(\a[29] ), .o1(new_n295));
  inv000aa1d42x5               g200(.a(\b[28] ), .o1(new_n296));
  oa0022aa1n02x5               g201(.a(new_n284), .b(new_n283), .c(new_n296), .d(new_n295), .o(new_n297));
  aoi112aa1n02x5               g202(.a(new_n297), .b(new_n294), .c(new_n295), .d(new_n296), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n292), .o1(new_n299));
  oaoi03aa1n02x5               g204(.a(new_n295), .b(new_n296), .c(new_n287), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n299), .c(new_n275), .d(new_n260), .o1(new_n301));
  aoi022aa1n03x5               g206(.a(new_n301), .b(new_n294), .c(new_n293), .d(new_n298), .o1(\s[30] ));
  nanp03aa1n02x5               g207(.a(new_n280), .b(new_n282), .c(new_n294), .o1(new_n303));
  nanb02aa1n03x5               g208(.a(new_n303), .b(new_n267), .out0(new_n304));
  xorc02aa1n02x5               g209(.a(\a[31] ), .b(\b[30] ), .out0(new_n305));
  oao003aa1n02x5               g210(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n306));
  norb02aa1n02x5               g211(.a(new_n306), .b(new_n305), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n306), .b(new_n303), .c(new_n275), .d(new_n260), .o1(new_n308));
  aoi022aa1n03x5               g213(.a(new_n308), .b(new_n305), .c(new_n304), .d(new_n307), .o1(\s[31] ));
  xnbna2aa1n03x5               g214(.a(new_n108), .b(new_n102), .c(new_n103), .out0(\s[3] ));
  nanb02aa1n02x5               g215(.a(\b[3] ), .b(new_n99), .out0(new_n311));
  aob012aa1n02x5               g216(.a(new_n102), .b(new_n311), .c(new_n112), .out0(new_n312));
  oab012aa1n02x4               g217(.a(new_n312), .b(new_n104), .c(new_n108), .out0(new_n313));
  aoi013aa1n02x4               g218(.a(new_n313), .b(new_n109), .c(new_n112), .d(new_n311), .o1(\s[4] ));
  xnbna2aa1n03x5               g219(.a(new_n113), .b(new_n109), .c(new_n112), .out0(\s[5] ));
  xorc02aa1n02x5               g220(.a(\a[6] ), .b(\b[5] ), .out0(new_n316));
  inv000aa1d42x5               g221(.a(new_n122), .o1(new_n317));
  nanb03aa1n02x5               g222(.a(new_n113), .b(new_n109), .c(new_n112), .out0(new_n318));
  xnbna2aa1n03x5               g223(.a(new_n316), .b(new_n318), .c(new_n317), .out0(\s[6] ));
  tech160nm_fiao0012aa1n02p5x5 g224(.a(new_n123), .b(new_n109), .c(new_n114), .o(new_n320));
  xorb03aa1n02x5               g225(.a(new_n320), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  norb02aa1n02x5               g226(.a(new_n115), .b(new_n116), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n322), .b(new_n117), .c(new_n320), .d(new_n118), .o1(new_n323));
  aoi112aa1n02x5               g228(.a(new_n322), .b(new_n117), .c(new_n320), .d(new_n118), .o1(new_n324));
  norb02aa1n02x5               g229(.a(new_n323), .b(new_n324), .out0(\s[8] ));
  xorb03aa1n02x5               g230(.a(new_n155), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


