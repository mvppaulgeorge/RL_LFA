// Benchmark "adder" written by ABC on Wed Jul 17 19:38:42 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n319, new_n322, new_n323, new_n324, new_n326, new_n328;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  xnrc02aa1n12x5               g003(.a(\b[3] ), .b(\a[4] ), .out0(new_n99));
  tech160nm_fixnrc02aa1n05x5   g004(.a(\b[2] ), .b(\a[3] ), .out0(new_n100));
  nor042aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nand22aa1n09x5               g006(.a(\b[0] ), .b(\a[1] ), .o1(new_n102));
  tech160nm_finand02aa1n03p5x5 g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  oaih12aa1n06x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .o1(new_n104));
  nor002aa1d32x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  inv030aa1n02x5               g010(.a(new_n105), .o1(new_n106));
  oao003aa1n06x5               g011(.a(\a[4] ), .b(\b[3] ), .c(new_n106), .carry(new_n107));
  oai013aa1n09x5               g012(.a(new_n107), .b(new_n100), .c(new_n99), .d(new_n104), .o1(new_n108));
  xnrc02aa1n12x5               g013(.a(\b[7] ), .b(\a[8] ), .out0(new_n109));
  xnrc02aa1n12x5               g014(.a(\b[6] ), .b(\a[7] ), .out0(new_n110));
  nor042aa1n12x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand22aa1n04x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nor042aa1n06x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand42aa1n16x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nona23aa1n09x5               g019(.a(new_n114), .b(new_n112), .c(new_n111), .d(new_n113), .out0(new_n115));
  nor043aa1n03x5               g020(.a(new_n115), .b(new_n110), .c(new_n109), .o1(new_n116));
  aoi012aa1n12x5               g021(.a(new_n113), .b(new_n111), .c(new_n114), .o1(new_n117));
  nor042aa1n06x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  inv000aa1n02x5               g023(.a(new_n118), .o1(new_n119));
  oao003aa1n03x5               g024(.a(\a[8] ), .b(\b[7] ), .c(new_n119), .carry(new_n120));
  oai013aa1d12x5               g025(.a(new_n120), .b(new_n110), .c(new_n109), .d(new_n117), .o1(new_n121));
  tech160nm_fixorc02aa1n03p5x5 g026(.a(\a[9] ), .b(\b[8] ), .out0(new_n122));
  aoai13aa1n02x5               g027(.a(new_n122), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n123));
  xorc02aa1n12x5               g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  xnbna2aa1n03x5               g029(.a(new_n124), .b(new_n123), .c(new_n98), .out0(\s[10] ));
  inv030aa1n02x5               g030(.a(new_n99), .o1(new_n126));
  nona22aa1n09x5               g031(.a(new_n126), .b(new_n100), .c(new_n104), .out0(new_n127));
  inv030aa1n02x5               g032(.a(new_n109), .o1(new_n128));
  inv030aa1n02x5               g033(.a(new_n110), .o1(new_n129));
  nanb03aa1n06x5               g034(.a(new_n115), .b(new_n128), .c(new_n129), .out0(new_n130));
  nor003aa1n02x5               g035(.a(new_n109), .b(new_n110), .c(new_n117), .o1(new_n131));
  norb02aa1n03x5               g036(.a(new_n120), .b(new_n131), .out0(new_n132));
  aoai13aa1n06x5               g037(.a(new_n132), .b(new_n130), .c(new_n127), .d(new_n107), .o1(new_n133));
  and002aa1n02x5               g038(.a(new_n124), .b(new_n122), .o(new_n134));
  norp02aa1n02x5               g039(.a(\b[9] ), .b(\a[10] ), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(\b[9] ), .b(\a[10] ), .o1(new_n136));
  tech160nm_fioai012aa1n05x5   g041(.a(new_n136), .b(new_n135), .c(new_n97), .o1(new_n137));
  aob012aa1n03x5               g042(.a(new_n137), .b(new_n133), .c(new_n134), .out0(new_n138));
  xorb03aa1n02x5               g043(.a(new_n138), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nand02aa1n06x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  norp02aa1n12x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand42aa1n04x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nanb02aa1n02x5               g049(.a(new_n143), .b(new_n144), .out0(new_n145));
  aoai13aa1n03x5               g050(.a(new_n145), .b(new_n140), .c(new_n138), .d(new_n142), .o1(new_n146));
  nona22aa1n02x4               g051(.a(new_n144), .b(new_n143), .c(new_n140), .out0(new_n147));
  aoai13aa1n02x5               g052(.a(new_n146), .b(new_n147), .c(new_n142), .d(new_n138), .o1(\s[12] ));
  nona23aa1n03x5               g053(.a(new_n144), .b(new_n141), .c(new_n140), .d(new_n143), .out0(new_n149));
  nano22aa1n02x4               g054(.a(new_n149), .b(new_n122), .c(new_n124), .out0(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n151));
  oaih12aa1n02x5               g056(.a(new_n144), .b(new_n143), .c(new_n140), .o1(new_n152));
  tech160nm_fioai012aa1n05x5   g057(.a(new_n152), .b(new_n149), .c(new_n137), .o1(new_n153));
  inv000aa1n03x5               g058(.a(new_n153), .o1(new_n154));
  nanp02aa1n03x5               g059(.a(new_n151), .b(new_n154), .o1(new_n155));
  xorb03aa1n02x5               g060(.a(new_n155), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n09x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  nand42aa1d28x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nano22aa1n03x7               g063(.a(new_n157), .b(new_n155), .c(new_n158), .out0(new_n159));
  nor042aa1n06x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1d28x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nanb02aa1n02x5               g066(.a(new_n160), .b(new_n161), .out0(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n157), .c(new_n155), .d(new_n158), .o1(new_n163));
  nona22aa1n02x4               g068(.a(new_n161), .b(new_n160), .c(new_n157), .out0(new_n164));
  oai012aa1n03x5               g069(.a(new_n163), .b(new_n159), .c(new_n164), .o1(\s[14] ));
  nano23aa1d15x5               g070(.a(new_n157), .b(new_n160), .c(new_n161), .d(new_n158), .out0(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  aoi022aa1n02x5               g072(.a(new_n153), .b(new_n166), .c(new_n161), .d(new_n164), .o1(new_n168));
  tech160nm_fioai012aa1n03p5x5 g073(.a(new_n168), .b(new_n151), .c(new_n167), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1d18x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  tech160nm_finand02aa1n03p5x5 g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nanb02aa1n06x5               g077(.a(new_n171), .b(new_n172), .out0(new_n173));
  oaoi13aa1n02x7               g078(.a(new_n173), .b(new_n168), .c(new_n151), .d(new_n167), .o1(new_n174));
  norp02aa1n12x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand02aa1n06x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nanb02aa1n09x5               g081(.a(new_n175), .b(new_n176), .out0(new_n177));
  aoai13aa1n03x5               g082(.a(new_n177), .b(new_n171), .c(new_n169), .d(new_n172), .o1(new_n178));
  norb03aa1n02x5               g083(.a(new_n176), .b(new_n171), .c(new_n175), .out0(new_n179));
  oaib12aa1n03x5               g084(.a(new_n178), .b(new_n174), .c(new_n179), .out0(\s[16] ));
  nano23aa1n06x5               g085(.a(new_n140), .b(new_n143), .c(new_n144), .d(new_n141), .out0(new_n181));
  nona22aa1d24x5               g086(.a(new_n166), .b(new_n173), .c(new_n177), .out0(new_n182));
  nano32aa1d12x5               g087(.a(new_n182), .b(new_n181), .c(new_n124), .d(new_n122), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n121), .c(new_n108), .d(new_n116), .o1(new_n184));
  oai012aa1n02x5               g089(.a(new_n161), .b(new_n160), .c(new_n157), .o1(new_n185));
  aoi012aa1n02x5               g090(.a(new_n175), .b(new_n171), .c(new_n176), .o1(new_n186));
  oai013aa1n02x4               g091(.a(new_n186), .b(new_n185), .c(new_n173), .d(new_n177), .o1(new_n187));
  aoib12aa1n09x5               g092(.a(new_n187), .b(new_n153), .c(new_n182), .out0(new_n188));
  xorc02aa1n12x5               g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  xnbna2aa1n03x5               g094(.a(new_n189), .b(new_n184), .c(new_n188), .out0(\s[17] ));
  inv040aa1d30x5               g095(.a(\a[17] ), .o1(new_n191));
  nanb02aa1d24x5               g096(.a(\b[16] ), .b(new_n191), .out0(new_n192));
  oabi12aa1n06x5               g097(.a(new_n187), .b(new_n154), .c(new_n182), .out0(new_n193));
  aoai13aa1n03x5               g098(.a(new_n189), .b(new_n193), .c(new_n133), .d(new_n183), .o1(new_n194));
  xorc02aa1n12x5               g099(.a(\a[18] ), .b(\b[17] ), .out0(new_n195));
  xnbna2aa1n03x5               g100(.a(new_n195), .b(new_n194), .c(new_n192), .out0(\s[18] ));
  inv000aa1d42x5               g101(.a(\a[18] ), .o1(new_n197));
  xroi22aa1d06x4               g102(.a(new_n191), .b(\b[16] ), .c(new_n197), .d(\b[17] ), .out0(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n193), .c(new_n133), .d(new_n183), .o1(new_n199));
  nor042aa1n04x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nand42aa1n04x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nanb02aa1n02x5               g106(.a(new_n200), .b(new_n201), .out0(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  oaoi03aa1n12x5               g108(.a(\a[18] ), .b(\b[17] ), .c(new_n192), .o1(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n203), .b(new_n199), .c(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g112(.a(new_n198), .o1(new_n208));
  aoai13aa1n02x7               g113(.a(new_n205), .b(new_n208), .c(new_n184), .d(new_n188), .o1(new_n209));
  nor042aa1n04x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  nand02aa1d16x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nanb02aa1n02x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  aoai13aa1n03x5               g117(.a(new_n212), .b(new_n200), .c(new_n209), .d(new_n203), .o1(new_n213));
  norb03aa1n02x5               g118(.a(new_n211), .b(new_n200), .c(new_n210), .out0(new_n214));
  aoai13aa1n02x5               g119(.a(new_n214), .b(new_n202), .c(new_n199), .d(new_n205), .o1(new_n215));
  nanp02aa1n03x5               g120(.a(new_n213), .b(new_n215), .o1(\s[20] ));
  nano23aa1n09x5               g121(.a(new_n200), .b(new_n210), .c(new_n211), .d(new_n201), .out0(new_n217));
  nand23aa1n06x5               g122(.a(new_n217), .b(new_n189), .c(new_n195), .o1(new_n218));
  oaih12aa1n02x5               g123(.a(new_n211), .b(new_n210), .c(new_n200), .o1(new_n219));
  aobi12aa1n06x5               g124(.a(new_n219), .b(new_n217), .c(new_n204), .out0(new_n220));
  aoai13aa1n06x5               g125(.a(new_n220), .b(new_n218), .c(new_n184), .d(new_n188), .o1(new_n221));
  xorb03aa1n02x5               g126(.a(new_n221), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nand02aa1d24x5               g128(.a(\b[20] ), .b(\a[21] ), .o1(new_n224));
  nor042aa1n04x5               g129(.a(\b[21] ), .b(\a[22] ), .o1(new_n225));
  nand02aa1n16x5               g130(.a(\b[21] ), .b(\a[22] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  inv000aa1d42x5               g132(.a(new_n227), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n228), .b(new_n223), .c(new_n221), .d(new_n224), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n218), .o1(new_n230));
  aoai13aa1n02x5               g135(.a(new_n230), .b(new_n193), .c(new_n133), .d(new_n183), .o1(new_n231));
  nanb02aa1n02x5               g136(.a(new_n223), .b(new_n224), .out0(new_n232));
  norb03aa1n02x5               g137(.a(new_n226), .b(new_n223), .c(new_n225), .out0(new_n233));
  aoai13aa1n02x5               g138(.a(new_n233), .b(new_n232), .c(new_n231), .d(new_n220), .o1(new_n234));
  nanp02aa1n03x5               g139(.a(new_n229), .b(new_n234), .o1(\s[22] ));
  nano23aa1n06x5               g140(.a(new_n223), .b(new_n225), .c(new_n226), .d(new_n224), .out0(new_n236));
  nanp03aa1n02x5               g141(.a(new_n198), .b(new_n217), .c(new_n236), .o1(new_n237));
  inv000aa1n02x5               g142(.a(new_n220), .o1(new_n238));
  inv020aa1n02x5               g143(.a(new_n223), .o1(new_n239));
  tech160nm_fioaoi03aa1n04x5   g144(.a(\a[22] ), .b(\b[21] ), .c(new_n239), .o1(new_n240));
  aoi012aa1n02x5               g145(.a(new_n240), .b(new_n238), .c(new_n236), .o1(new_n241));
  aoai13aa1n04x5               g146(.a(new_n241), .b(new_n237), .c(new_n184), .d(new_n188), .o1(new_n242));
  xorb03aa1n02x5               g147(.a(new_n242), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1d32x5               g148(.a(\b[22] ), .b(\a[23] ), .o1(new_n244));
  nand02aa1d24x5               g149(.a(\b[22] ), .b(\a[23] ), .o1(new_n245));
  norb02aa1n02x5               g150(.a(new_n245), .b(new_n244), .out0(new_n246));
  nor002aa1d24x5               g151(.a(\b[23] ), .b(\a[24] ), .o1(new_n247));
  nand02aa1d28x5               g152(.a(\b[23] ), .b(\a[24] ), .o1(new_n248));
  nanb02aa1n02x5               g153(.a(new_n247), .b(new_n248), .out0(new_n249));
  aoai13aa1n03x5               g154(.a(new_n249), .b(new_n244), .c(new_n242), .d(new_n246), .o1(new_n250));
  nand02aa1n02x5               g155(.a(new_n242), .b(new_n246), .o1(new_n251));
  nona22aa1d24x5               g156(.a(new_n248), .b(new_n247), .c(new_n244), .out0(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  tech160nm_finand02aa1n03p5x5 g158(.a(new_n251), .b(new_n253), .o1(new_n254));
  nanp02aa1n03x5               g159(.a(new_n250), .b(new_n254), .o1(\s[24] ));
  nano23aa1n06x5               g160(.a(new_n244), .b(new_n247), .c(new_n248), .d(new_n245), .out0(new_n256));
  nand02aa1d06x5               g161(.a(new_n256), .b(new_n236), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n257), .o1(new_n258));
  nanb02aa1n02x5               g163(.a(new_n218), .b(new_n258), .out0(new_n259));
  nand22aa1n03x5               g164(.a(new_n217), .b(new_n204), .o1(new_n260));
  aoi022aa1n06x5               g165(.a(new_n256), .b(new_n240), .c(new_n248), .d(new_n252), .o1(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n257), .c(new_n260), .d(new_n219), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  aoai13aa1n04x5               g168(.a(new_n263), .b(new_n259), .c(new_n184), .d(new_n188), .o1(new_n264));
  xorb03aa1n02x5               g169(.a(new_n264), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g170(.a(\b[24] ), .b(\a[25] ), .o1(new_n266));
  tech160nm_fixorc02aa1n03p5x5 g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[25] ), .b(\a[26] ), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n266), .c(new_n264), .d(new_n267), .o1(new_n269));
  nand02aa1n02x5               g174(.a(new_n264), .b(new_n267), .o1(new_n270));
  norp02aa1n02x5               g175(.a(new_n268), .b(new_n266), .o1(new_n271));
  tech160nm_finand02aa1n03p5x5 g176(.a(new_n270), .b(new_n271), .o1(new_n272));
  nanp02aa1n03x5               g177(.a(new_n269), .b(new_n272), .o1(\s[26] ));
  norb02aa1n02x5               g178(.a(new_n267), .b(new_n268), .out0(new_n274));
  norb03aa1n03x5               g179(.a(new_n274), .b(new_n218), .c(new_n257), .out0(new_n275));
  inv000aa1n02x5               g180(.a(new_n275), .o1(new_n276));
  oaoi03aa1n02x5               g181(.a(\a[26] ), .b(\b[25] ), .c(new_n271), .o1(new_n277));
  aoi012aa1n06x5               g182(.a(new_n277), .b(new_n262), .c(new_n274), .o1(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n276), .c(new_n184), .d(new_n188), .o1(new_n279));
  xorb03aa1n03x5               g184(.a(new_n279), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g185(.a(\b[26] ), .b(\a[27] ), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnrc02aa1n12x5               g187(.a(\b[27] ), .b(\a[28] ), .out0(new_n283));
  aoai13aa1n03x5               g188(.a(new_n283), .b(new_n281), .c(new_n279), .d(new_n282), .o1(new_n284));
  aoai13aa1n03x5               g189(.a(new_n275), .b(new_n193), .c(new_n133), .d(new_n183), .o1(new_n285));
  inv000aa1d42x5               g190(.a(new_n282), .o1(new_n286));
  nor042aa1n03x5               g191(.a(new_n283), .b(new_n281), .o1(new_n287));
  aoai13aa1n02x5               g192(.a(new_n287), .b(new_n286), .c(new_n285), .d(new_n278), .o1(new_n288));
  nanp02aa1n03x5               g193(.a(new_n284), .b(new_n288), .o1(\s[28] ));
  norb02aa1n03x5               g194(.a(new_n282), .b(new_n283), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  xorc02aa1n12x5               g196(.a(\a[29] ), .b(\b[28] ), .out0(new_n292));
  inv000aa1d42x5               g197(.a(new_n292), .o1(new_n293));
  tech160nm_fiaoi012aa1n05x5   g198(.a(new_n287), .b(\a[28] ), .c(\b[27] ), .o1(new_n294));
  norp02aa1n02x5               g199(.a(new_n294), .b(new_n293), .o1(new_n295));
  aoai13aa1n02x5               g200(.a(new_n295), .b(new_n291), .c(new_n285), .d(new_n278), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n293), .b(new_n294), .c(new_n279), .d(new_n290), .o1(new_n297));
  nanp02aa1n03x5               g202(.a(new_n297), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n102), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g204(.a(new_n283), .b(new_n282), .c(new_n292), .out0(new_n300));
  nand02aa1n02x5               g205(.a(new_n279), .b(new_n300), .o1(new_n301));
  norp02aa1n02x5               g206(.a(\b[28] ), .b(\a[29] ), .o1(new_n302));
  aoi012aa1n02x5               g207(.a(new_n302), .b(new_n294), .c(new_n292), .o1(new_n303));
  xorc02aa1n02x5               g208(.a(\a[30] ), .b(\b[29] ), .out0(new_n304));
  inv000aa1n02x5               g209(.a(new_n300), .o1(new_n305));
  oai012aa1n02x5               g210(.a(new_n304), .b(\b[28] ), .c(\a[29] ), .o1(new_n306));
  tech160nm_fiaoi012aa1n05x5   g211(.a(new_n306), .b(new_n294), .c(new_n292), .o1(new_n307));
  aoai13aa1n02x7               g212(.a(new_n307), .b(new_n305), .c(new_n285), .d(new_n278), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n304), .c(new_n301), .d(new_n303), .o1(\s[30] ));
  nano23aa1n09x5               g214(.a(new_n293), .b(new_n283), .c(new_n304), .d(new_n282), .out0(new_n310));
  inv000aa1d42x5               g215(.a(new_n310), .o1(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[30] ), .b(\a[31] ), .out0(new_n312));
  aoi012aa1n02x5               g217(.a(new_n307), .b(\a[30] ), .c(\b[29] ), .o1(new_n313));
  norp02aa1n02x5               g218(.a(new_n313), .b(new_n312), .o1(new_n314));
  aoai13aa1n02x7               g219(.a(new_n314), .b(new_n311), .c(new_n285), .d(new_n278), .o1(new_n315));
  aoai13aa1n03x5               g220(.a(new_n312), .b(new_n313), .c(new_n279), .d(new_n310), .o1(new_n316));
  nanp02aa1n03x5               g221(.a(new_n316), .b(new_n315), .o1(\s[31] ));
  xnrb03aa1n02x5               g222(.a(new_n104), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  orn002aa1n02x5               g223(.a(new_n100), .b(new_n104), .o(new_n319));
  xnbna2aa1n03x5               g224(.a(new_n126), .b(new_n319), .c(new_n106), .out0(\s[4] ));
  xorb03aa1n02x5               g225(.a(new_n108), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g226(.a(new_n113), .b(new_n114), .out0(new_n322));
  aoai13aa1n02x5               g227(.a(new_n322), .b(new_n111), .c(new_n108), .d(new_n112), .o1(new_n323));
  aoi112aa1n02x5               g228(.a(new_n111), .b(new_n322), .c(new_n108), .d(new_n112), .o1(new_n324));
  nanb02aa1n02x5               g229(.a(new_n324), .b(new_n323), .out0(\s[6] ));
  aoai13aa1n02x5               g230(.a(new_n117), .b(new_n115), .c(new_n127), .d(new_n107), .o1(new_n326));
  xorb03aa1n02x5               g231(.a(new_n326), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanp02aa1n02x5               g232(.a(new_n326), .b(new_n129), .o1(new_n328));
  xnbna2aa1n03x5               g233(.a(new_n128), .b(new_n328), .c(new_n119), .out0(\s[8] ));
  xorb03aa1n02x5               g234(.a(new_n133), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


