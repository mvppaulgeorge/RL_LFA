// Benchmark "adder" written by ABC on Wed Jul 17 19:43:37 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n285, new_n286, new_n287, new_n288,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n338,
    new_n339, new_n341, new_n342, new_n343, new_n345, new_n346, new_n348,
    new_n349, new_n351;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1d32x5               g002(.a(\b[2] ), .b(\a[3] ), .o1(new_n98));
  and002aa1n12x5               g003(.a(\b[3] ), .b(\a[4] ), .o(new_n99));
  nor002aa1n03x5               g004(.a(\b[3] ), .b(\a[4] ), .o1(new_n100));
  nor043aa1n06x5               g005(.a(new_n99), .b(new_n100), .c(new_n98), .o1(new_n101));
  nand42aa1n03x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanb02aa1n06x5               g007(.a(new_n98), .b(new_n102), .out0(new_n103));
  nor002aa1n08x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand22aa1n09x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nand42aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  oai012aa1n12x5               g011(.a(new_n106), .b(new_n104), .c(new_n105), .o1(new_n107));
  oaih12aa1n12x5               g012(.a(new_n101), .b(new_n107), .c(new_n103), .o1(new_n108));
  nor042aa1n09x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  aoi022aa1n06x5               g014(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n110));
  nor042aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nona22aa1n02x4               g016(.a(new_n110), .b(new_n111), .c(new_n109), .out0(new_n112));
  nor042aa1n06x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  aoi022aa1d24x5               g018(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n114));
  nand22aa1n04x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nor022aa1n08x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n114), .b(new_n115), .c(new_n116), .d(new_n113), .out0(new_n117));
  nona22aa1n03x5               g022(.a(new_n108), .b(new_n117), .c(new_n112), .out0(new_n118));
  nand42aa1n02x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nand42aa1n06x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nano22aa1n03x7               g025(.a(new_n113), .b(new_n119), .c(new_n120), .out0(new_n121));
  norb02aa1n03x5               g026(.a(new_n115), .b(new_n116), .out0(new_n122));
  inv040aa1n02x5               g027(.a(new_n109), .o1(new_n123));
  oai112aa1n02x5               g028(.a(new_n123), .b(new_n120), .c(\b[4] ), .d(\a[5] ), .o1(new_n124));
  tech160nm_fiaoi012aa1n04x5   g029(.a(new_n116), .b(new_n113), .c(new_n115), .o1(new_n125));
  inv000aa1n02x5               g030(.a(new_n125), .o1(new_n126));
  aoi013aa1n06x4               g031(.a(new_n126), .b(new_n124), .c(new_n121), .d(new_n122), .o1(new_n127));
  nand02aa1d06x5               g032(.a(new_n118), .b(new_n127), .o1(new_n128));
  nanp02aa1n02x5               g033(.a(\b[8] ), .b(\a[9] ), .o1(new_n129));
  aoi012aa1n02x5               g034(.a(new_n97), .b(new_n128), .c(new_n129), .o1(new_n130));
  xorc02aa1n02x5               g035(.a(\a[10] ), .b(\b[9] ), .out0(new_n131));
  nor042aa1n03x5               g036(.a(new_n117), .b(new_n112), .o1(new_n132));
  norb03aa1n09x5               g037(.a(new_n120), .b(new_n109), .c(new_n111), .out0(new_n133));
  tech160nm_fioai012aa1n05x5   g038(.a(new_n125), .b(new_n117), .c(new_n133), .o1(new_n134));
  aoi012aa1n12x5               g039(.a(new_n134), .b(new_n132), .c(new_n108), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n129), .b(new_n97), .out0(new_n136));
  nand42aa1d28x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  oaih22aa1n06x5               g043(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n139));
  norp02aa1n02x5               g044(.a(new_n139), .b(new_n138), .o1(new_n140));
  oaib12aa1n02x5               g045(.a(new_n140), .b(new_n135), .c(new_n136), .out0(new_n141));
  oai012aa1n02x5               g046(.a(new_n141), .b(new_n130), .c(new_n131), .o1(\s[10] ));
  nand42aa1n08x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nor002aa1d32x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nano22aa1n03x7               g049(.a(new_n144), .b(new_n137), .c(new_n143), .out0(new_n145));
  aoai13aa1n06x5               g050(.a(new_n145), .b(new_n139), .c(new_n128), .d(new_n136), .o1(new_n146));
  nanb02aa1n02x5               g051(.a(new_n144), .b(new_n143), .out0(new_n147));
  aoai13aa1n02x5               g052(.a(new_n137), .b(new_n139), .c(new_n128), .d(new_n136), .o1(new_n148));
  aobi12aa1n02x5               g053(.a(new_n146), .b(new_n148), .c(new_n147), .out0(\s[11] ));
  orn002aa1n02x5               g054(.a(\a[11] ), .b(\b[10] ), .o(new_n150));
  xorc02aa1n02x5               g055(.a(\a[12] ), .b(\b[11] ), .out0(new_n151));
  xnbna2aa1n03x5               g056(.a(new_n151), .b(new_n146), .c(new_n150), .out0(\s[12] ));
  inv040aa1d32x5               g057(.a(\a[12] ), .o1(new_n153));
  inv030aa1d32x5               g058(.a(\b[11] ), .o1(new_n154));
  nand22aa1n03x5               g059(.a(new_n154), .b(new_n153), .o1(new_n155));
  nand02aa1n02x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  nand02aa1d04x5               g061(.a(new_n155), .b(new_n156), .o1(new_n157));
  nona23aa1n02x4               g062(.a(new_n145), .b(new_n129), .c(new_n157), .d(new_n139), .out0(new_n158));
  nanb03aa1n12x5               g063(.a(new_n144), .b(new_n137), .c(new_n143), .out0(new_n159));
  oaoi03aa1n06x5               g064(.a(new_n153), .b(new_n154), .c(new_n144), .o1(new_n160));
  oai013aa1n02x4               g065(.a(new_n160), .b(new_n140), .c(new_n159), .d(new_n157), .o1(new_n161));
  oabi12aa1n06x5               g066(.a(new_n161), .b(new_n135), .c(new_n158), .out0(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1d18x5               g068(.a(\b[12] ), .b(\a[13] ), .o1(new_n164));
  nanp02aa1n04x5               g069(.a(\b[12] ), .b(\a[13] ), .o1(new_n165));
  nor002aa1d32x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nand02aa1d28x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  aoi112aa1n02x5               g073(.a(new_n164), .b(new_n168), .c(new_n162), .d(new_n165), .o1(new_n169));
  aoai13aa1n02x5               g074(.a(new_n168), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(\s[14] ));
  oab012aa1n06x5               g076(.a(new_n97), .b(\a[10] ), .c(\b[9] ), .out0(new_n172));
  nano23aa1n03x7               g077(.a(new_n159), .b(new_n157), .c(new_n172), .d(new_n129), .out0(new_n173));
  nano23aa1n09x5               g078(.a(new_n164), .b(new_n166), .c(new_n167), .d(new_n165), .out0(new_n174));
  aoai13aa1n06x5               g079(.a(new_n174), .b(new_n161), .c(new_n128), .d(new_n173), .o1(new_n175));
  aoi012aa1d24x5               g080(.a(new_n166), .b(new_n164), .c(new_n167), .o1(new_n176));
  nor002aa1d32x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  nanp02aa1n06x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nanb02aa1n02x5               g083(.a(new_n177), .b(new_n178), .out0(new_n179));
  xobna2aa1n03x5               g084(.a(new_n179), .b(new_n175), .c(new_n176), .out0(\s[15] ));
  tech160nm_fiao0012aa1n02p5x5 g085(.a(new_n179), .b(new_n175), .c(new_n176), .o(new_n181));
  nor042aa1n06x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nand02aa1n04x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  norb02aa1n02x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  aoib12aa1n02x5               g089(.a(new_n177), .b(new_n183), .c(new_n182), .out0(new_n185));
  inv000aa1d42x5               g090(.a(new_n177), .o1(new_n186));
  aoai13aa1n02x7               g091(.a(new_n186), .b(new_n179), .c(new_n175), .d(new_n176), .o1(new_n187));
  aoi022aa1n03x5               g092(.a(new_n181), .b(new_n185), .c(new_n187), .d(new_n184), .o1(\s[16] ));
  nona23aa1n03x5               g093(.a(new_n167), .b(new_n165), .c(new_n164), .d(new_n166), .out0(new_n189));
  nona23aa1d18x5               g094(.a(new_n183), .b(new_n178), .c(new_n177), .d(new_n182), .out0(new_n190));
  nor042aa1n03x5               g095(.a(new_n190), .b(new_n189), .o1(new_n191));
  nand22aa1n03x5               g096(.a(new_n173), .b(new_n191), .o1(new_n192));
  aoi112aa1n03x5               g097(.a(new_n159), .b(new_n157), .c(new_n172), .d(new_n137), .o1(new_n193));
  inv000aa1n02x5               g098(.a(new_n160), .o1(new_n194));
  tech160nm_fioai012aa1n03p5x5 g099(.a(new_n183), .b(new_n182), .c(new_n177), .o1(new_n195));
  tech160nm_fioai012aa1n04x5   g100(.a(new_n195), .b(new_n190), .c(new_n176), .o1(new_n196));
  oaoi13aa1n12x5               g101(.a(new_n196), .b(new_n191), .c(new_n193), .d(new_n194), .o1(new_n197));
  oai012aa1d24x5               g102(.a(new_n197), .b(new_n135), .c(new_n192), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nor042aa1n04x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  tech160nm_fixorc02aa1n03p5x5 g105(.a(\a[17] ), .b(\b[16] ), .out0(new_n201));
  nor022aa1n08x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nand42aa1n16x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  norb02aa1n03x5               g108(.a(new_n203), .b(new_n202), .out0(new_n204));
  aoi112aa1n02x5               g109(.a(new_n200), .b(new_n204), .c(new_n198), .d(new_n201), .o1(new_n205));
  aoai13aa1n02x5               g110(.a(new_n204), .b(new_n200), .c(new_n198), .d(new_n201), .o1(new_n206));
  norb02aa1n02x5               g111(.a(new_n206), .b(new_n205), .out0(\s[18] ));
  and002aa1n06x5               g112(.a(new_n201), .b(new_n204), .o(new_n208));
  aoi012aa1d18x5               g113(.a(new_n202), .b(new_n200), .c(new_n203), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor042aa1n04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  tech160nm_finand02aa1n05x5   g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  nanb02aa1d24x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  inv000aa1d42x5               g118(.a(new_n213), .o1(new_n214));
  aoai13aa1n12x5               g119(.a(new_n214), .b(new_n210), .c(new_n198), .d(new_n208), .o1(new_n215));
  aoi112aa1n02x5               g120(.a(new_n214), .b(new_n210), .c(new_n198), .d(new_n208), .o1(new_n216));
  norb02aa1n03x4               g121(.a(new_n215), .b(new_n216), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g123(.a(\a[20] ), .o1(new_n219));
  inv030aa1d32x5               g124(.a(\b[19] ), .o1(new_n220));
  nand02aa1d04x5               g125(.a(new_n220), .b(new_n219), .o1(new_n221));
  nand22aa1n04x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand22aa1n09x5               g127(.a(new_n221), .b(new_n222), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoi012aa1n02x5               g129(.a(new_n211), .b(new_n221), .c(new_n222), .o1(new_n225));
  tech160nm_fioai012aa1n03p5x5 g130(.a(new_n215), .b(\b[18] ), .c(\a[19] ), .o1(new_n226));
  aoi022aa1n02x7               g131(.a(new_n226), .b(new_n224), .c(new_n215), .d(new_n225), .o1(\s[20] ));
  nano23aa1n02x4               g132(.a(new_n223), .b(new_n213), .c(new_n201), .d(new_n204), .out0(new_n228));
  oaoi03aa1n03x5               g133(.a(new_n219), .b(new_n220), .c(new_n211), .o1(new_n229));
  oai013aa1d12x5               g134(.a(new_n229), .b(new_n209), .c(new_n213), .d(new_n223), .o1(new_n230));
  nor042aa1n04x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  nand42aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  aoai13aa1n12x5               g138(.a(new_n233), .b(new_n230), .c(new_n198), .d(new_n228), .o1(new_n234));
  aoi112aa1n02x5               g139(.a(new_n233), .b(new_n230), .c(new_n198), .d(new_n228), .o1(new_n235));
  norb02aa1n03x4               g140(.a(new_n234), .b(new_n235), .out0(\s[21] ));
  nor022aa1n16x5               g141(.a(\b[21] ), .b(\a[22] ), .o1(new_n237));
  nand02aa1n04x5               g142(.a(\b[21] ), .b(\a[22] ), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n238), .b(new_n237), .out0(new_n239));
  aoib12aa1n02x5               g144(.a(new_n231), .b(new_n238), .c(new_n237), .out0(new_n240));
  tech160nm_fioai012aa1n03p5x5 g145(.a(new_n234), .b(\b[20] ), .c(\a[21] ), .o1(new_n241));
  aoi022aa1n02x7               g146(.a(new_n241), .b(new_n239), .c(new_n234), .d(new_n240), .o1(\s[22] ));
  nano23aa1n03x5               g147(.a(new_n177), .b(new_n182), .c(new_n183), .d(new_n178), .out0(new_n243));
  nanp02aa1n02x5               g148(.a(new_n243), .b(new_n174), .o1(new_n244));
  nor042aa1n03x5               g149(.a(new_n158), .b(new_n244), .o1(new_n245));
  oai112aa1n02x5               g150(.a(new_n145), .b(new_n151), .c(new_n139), .d(new_n138), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n176), .o1(new_n247));
  aobi12aa1n02x5               g152(.a(new_n195), .b(new_n243), .c(new_n247), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n244), .c(new_n246), .d(new_n160), .o1(new_n249));
  nor042aa1n04x5               g154(.a(new_n213), .b(new_n223), .o1(new_n250));
  nona23aa1n09x5               g155(.a(new_n238), .b(new_n232), .c(new_n231), .d(new_n237), .out0(new_n251));
  nano32aa1n02x4               g156(.a(new_n251), .b(new_n250), .c(new_n204), .d(new_n201), .out0(new_n252));
  aoai13aa1n06x5               g157(.a(new_n252), .b(new_n249), .c(new_n128), .d(new_n245), .o1(new_n253));
  nano23aa1n06x5               g158(.a(new_n231), .b(new_n237), .c(new_n238), .d(new_n232), .out0(new_n254));
  ao0012aa1n12x5               g159(.a(new_n237), .b(new_n231), .c(new_n238), .o(new_n255));
  aoi012aa1n02x5               g160(.a(new_n255), .b(new_n230), .c(new_n254), .o1(new_n256));
  nor002aa1n16x5               g161(.a(\b[22] ), .b(\a[23] ), .o1(new_n257));
  nand42aa1n06x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  norb02aa1d21x5               g163(.a(new_n258), .b(new_n257), .out0(new_n259));
  aob012aa1n03x5               g164(.a(new_n259), .b(new_n253), .c(new_n256), .out0(new_n260));
  aoi112aa1n02x5               g165(.a(new_n259), .b(new_n255), .c(new_n230), .d(new_n254), .o1(new_n261));
  aobi12aa1n02x7               g166(.a(new_n260), .b(new_n261), .c(new_n253), .out0(\s[23] ));
  nor002aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .o1(new_n263));
  nand42aa1n06x5               g168(.a(\b[23] ), .b(\a[24] ), .o1(new_n264));
  norb02aa1n02x7               g169(.a(new_n264), .b(new_n263), .out0(new_n265));
  aoib12aa1n02x5               g170(.a(new_n257), .b(new_n264), .c(new_n263), .out0(new_n266));
  inv000aa1d42x5               g171(.a(new_n257), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n259), .o1(new_n268));
  aoai13aa1n02x5               g173(.a(new_n267), .b(new_n268), .c(new_n253), .d(new_n256), .o1(new_n269));
  aoi022aa1n02x7               g174(.a(new_n269), .b(new_n265), .c(new_n260), .d(new_n266), .o1(\s[24] ));
  nano23aa1n03x5               g175(.a(new_n257), .b(new_n263), .c(new_n264), .d(new_n258), .out0(new_n271));
  nanp02aa1n03x5               g176(.a(new_n271), .b(new_n254), .o1(new_n272));
  nano32aa1n03x7               g177(.a(new_n272), .b(new_n250), .c(new_n204), .d(new_n201), .out0(new_n273));
  and002aa1n02x5               g178(.a(new_n198), .b(new_n273), .o(new_n274));
  nona22aa1n03x5               g179(.a(new_n210), .b(new_n213), .c(new_n223), .out0(new_n275));
  oaoi03aa1n02x5               g180(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .o1(new_n276));
  aoi012aa1n06x5               g181(.a(new_n276), .b(new_n271), .c(new_n255), .o1(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n272), .c(new_n275), .d(new_n229), .o1(new_n278));
  xorc02aa1n12x5               g183(.a(\a[25] ), .b(\b[24] ), .out0(new_n279));
  aoai13aa1n06x5               g184(.a(new_n279), .b(new_n278), .c(new_n198), .d(new_n273), .o1(new_n280));
  nano22aa1n03x7               g185(.a(new_n251), .b(new_n259), .c(new_n265), .out0(new_n281));
  nand22aa1n04x5               g186(.a(new_n230), .b(new_n281), .o1(new_n282));
  nanb03aa1n02x5               g187(.a(new_n279), .b(new_n282), .c(new_n277), .out0(new_n283));
  oa0012aa1n03x5               g188(.a(new_n280), .b(new_n274), .c(new_n283), .o(\s[25] ));
  tech160nm_fixorc02aa1n05x5   g189(.a(\a[26] ), .b(\b[25] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(\a[25] ), .o1(new_n286));
  aoib12aa1n02x5               g191(.a(new_n285), .b(new_n286), .c(\b[24] ), .out0(new_n287));
  oaib12aa1n03x5               g192(.a(new_n280), .b(\b[24] ), .c(new_n286), .out0(new_n288));
  aoi022aa1n02x7               g193(.a(new_n288), .b(new_n285), .c(new_n280), .d(new_n287), .o1(\s[26] ));
  and002aa1n02x5               g194(.a(new_n285), .b(new_n279), .o(new_n290));
  inv030aa1n02x5               g195(.a(new_n290), .o1(new_n291));
  nano32aa1d12x5               g196(.a(new_n291), .b(new_n208), .c(new_n281), .d(new_n250), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n249), .c(new_n128), .d(new_n245), .o1(new_n293));
  nanp02aa1n02x5               g198(.a(\b[25] ), .b(\a[26] ), .o1(new_n294));
  oai022aa1n02x5               g199(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n295));
  aoi022aa1n06x5               g200(.a(new_n278), .b(new_n290), .c(new_n294), .d(new_n295), .o1(new_n296));
  xorc02aa1n02x5               g201(.a(\a[27] ), .b(\b[26] ), .out0(new_n297));
  xnbna2aa1n03x5               g202(.a(new_n297), .b(new_n293), .c(new_n296), .out0(\s[27] ));
  nanp02aa1n02x5               g203(.a(new_n295), .b(new_n294), .o1(new_n299));
  aoai13aa1n12x5               g204(.a(new_n299), .b(new_n291), .c(new_n282), .d(new_n277), .o1(new_n300));
  aoai13aa1n06x5               g205(.a(new_n297), .b(new_n300), .c(new_n198), .d(new_n292), .o1(new_n301));
  xorc02aa1n02x5               g206(.a(\a[28] ), .b(\b[27] ), .out0(new_n302));
  norp02aa1n02x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  norp02aa1n02x5               g208(.a(new_n302), .b(new_n303), .o1(new_n304));
  inv000aa1d42x5               g209(.a(\a[27] ), .o1(new_n305));
  oaib12aa1n06x5               g210(.a(new_n301), .b(\b[26] ), .c(new_n305), .out0(new_n306));
  aoi022aa1n02x7               g211(.a(new_n306), .b(new_n302), .c(new_n301), .d(new_n304), .o1(\s[28] ));
  inv000aa1d42x5               g212(.a(\a[28] ), .o1(new_n308));
  xroi22aa1d04x5               g213(.a(new_n305), .b(\b[26] ), .c(new_n308), .d(\b[27] ), .out0(new_n309));
  aoai13aa1n06x5               g214(.a(new_n309), .b(new_n300), .c(new_n198), .d(new_n292), .o1(new_n310));
  inv000aa1d42x5               g215(.a(\b[27] ), .o1(new_n311));
  oao003aa1n09x5               g216(.a(new_n308), .b(new_n311), .c(new_n303), .carry(new_n312));
  inv000aa1d42x5               g217(.a(new_n312), .o1(new_n313));
  nand42aa1n02x5               g218(.a(new_n310), .b(new_n313), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[29] ), .b(\b[28] ), .out0(new_n315));
  norp02aa1n02x5               g220(.a(new_n312), .b(new_n315), .o1(new_n316));
  aoi022aa1n02x7               g221(.a(new_n314), .b(new_n315), .c(new_n310), .d(new_n316), .o1(\s[29] ));
  xorb03aa1n02x5               g222(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g223(.a(new_n297), .b(new_n315), .c(new_n302), .o(new_n319));
  aoai13aa1n06x5               g224(.a(new_n319), .b(new_n300), .c(new_n198), .d(new_n292), .o1(new_n320));
  inv000aa1d42x5               g225(.a(\a[29] ), .o1(new_n321));
  inv000aa1d42x5               g226(.a(\b[28] ), .o1(new_n322));
  oaoi03aa1n02x5               g227(.a(new_n321), .b(new_n322), .c(new_n312), .o1(new_n323));
  nand42aa1n02x5               g228(.a(new_n320), .b(new_n323), .o1(new_n324));
  xorc02aa1n02x5               g229(.a(\a[30] ), .b(\b[29] ), .out0(new_n325));
  oabi12aa1n02x5               g230(.a(new_n325), .b(\a[29] ), .c(\b[28] ), .out0(new_n326));
  oaoi13aa1n02x5               g231(.a(new_n326), .b(new_n312), .c(new_n321), .d(new_n322), .o1(new_n327));
  aoi022aa1n02x7               g232(.a(new_n324), .b(new_n325), .c(new_n320), .d(new_n327), .o1(\s[30] ));
  xnrc02aa1n02x5               g233(.a(\b[30] ), .b(\a[31] ), .out0(new_n329));
  and003aa1n02x5               g234(.a(new_n309), .b(new_n325), .c(new_n315), .o(new_n330));
  aoai13aa1n03x5               g235(.a(new_n330), .b(new_n300), .c(new_n198), .d(new_n292), .o1(new_n331));
  oao003aa1n02x5               g236(.a(\a[30] ), .b(\b[29] ), .c(new_n323), .carry(new_n332));
  aoi012aa1n03x5               g237(.a(new_n329), .b(new_n331), .c(new_n332), .o1(new_n333));
  aobi12aa1n03x5               g238(.a(new_n330), .b(new_n293), .c(new_n296), .out0(new_n334));
  nano22aa1n02x4               g239(.a(new_n334), .b(new_n329), .c(new_n332), .out0(new_n335));
  nor002aa1n02x5               g240(.a(new_n333), .b(new_n335), .o1(\s[31] ));
  xnrb03aa1n02x5               g241(.a(new_n107), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  norp02aa1n02x5               g242(.a(new_n99), .b(new_n100), .o1(new_n338));
  oab012aa1n02x4               g243(.a(new_n98), .b(new_n107), .c(new_n103), .out0(new_n339));
  oai012aa1n02x5               g244(.a(new_n108), .b(new_n339), .c(new_n338), .o1(\s[4] ));
  norb02aa1n02x5               g245(.a(new_n110), .b(new_n111), .out0(new_n341));
  nanb02aa1n02x5               g246(.a(new_n99), .b(new_n108), .out0(new_n342));
  xnrc02aa1n02x5               g247(.a(\b[4] ), .b(\a[5] ), .out0(new_n343));
  aoi022aa1n02x5               g248(.a(new_n342), .b(new_n343), .c(new_n341), .d(new_n108), .o1(\s[5] ));
  aoi012aa1n02x5               g249(.a(new_n111), .b(new_n108), .c(new_n110), .o1(new_n345));
  aob012aa1n02x5               g250(.a(new_n133), .b(new_n108), .c(new_n341), .out0(new_n346));
  aoai13aa1n02x5               g251(.a(new_n346), .b(new_n345), .c(new_n123), .d(new_n120), .o1(\s[6] ));
  nanb02aa1n02x5               g252(.a(new_n113), .b(new_n119), .out0(new_n348));
  aoai13aa1n02x5               g253(.a(new_n120), .b(new_n124), .c(new_n108), .d(new_n341), .o1(new_n349));
  aoi022aa1n02x5               g254(.a(new_n349), .b(new_n348), .c(new_n346), .d(new_n121), .o1(\s[7] ));
  aoi012aa1n02x5               g255(.a(new_n113), .b(new_n346), .c(new_n114), .o1(new_n351));
  xnrc02aa1n02x5               g256(.a(new_n351), .b(new_n122), .out0(\s[8] ));
  xnbna2aa1n03x5               g257(.a(new_n136), .b(new_n118), .c(new_n127), .out0(\s[9] ));
endmodule


