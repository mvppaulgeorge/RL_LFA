// Benchmark "adder" written by ABC on Thu Jul 18 03:42:02 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n314, new_n315, new_n316, new_n318,
    new_n319, new_n321, new_n323, new_n324, new_n325, new_n327;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  inv000aa1d42x5               g003(.a(\a[3] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\a[4] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(\b[2] ), .o1(new_n101));
  aboi22aa1n03x5               g006(.a(\b[3] ), .b(new_n100), .c(new_n99), .d(new_n101), .out0(new_n102));
  xnrc02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .out0(new_n103));
  nanp02aa1n02x5               g008(.a(\b[1] ), .b(\a[2] ), .o1(new_n104));
  nand22aa1n04x5               g009(.a(\b[0] ), .b(\a[1] ), .o1(new_n105));
  nor042aa1n02x5               g010(.a(\b[1] ), .b(\a[2] ), .o1(new_n106));
  tech160nm_fioai012aa1n04x5   g011(.a(new_n104), .b(new_n106), .c(new_n105), .o1(new_n107));
  oai012aa1n06x5               g012(.a(new_n102), .b(new_n103), .c(new_n107), .o1(new_n108));
  nor022aa1n16x5               g013(.a(\b[5] ), .b(\a[6] ), .o1(new_n109));
  inv000aa1d42x5               g014(.a(new_n109), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  oai112aa1n02x5               g016(.a(new_n110), .b(new_n111), .c(\b[7] ), .d(\a[8] ), .o1(new_n112));
  inv000aa1d42x5               g017(.a(\a[5] ), .o1(new_n113));
  aoi022aa1n02x7               g018(.a(\b[4] ), .b(\a[5] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n114));
  oaib12aa1n02x5               g019(.a(new_n114), .b(\b[4] ), .c(new_n113), .out0(new_n115));
  inv000aa1d42x5               g020(.a(\a[8] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[7] ), .o1(new_n117));
  nor042aa1n02x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  inv000aa1n02x5               g023(.a(new_n118), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  oai112aa1n02x5               g025(.a(new_n119), .b(new_n120), .c(new_n117), .d(new_n116), .o1(new_n121));
  nor043aa1n03x5               g026(.a(new_n121), .b(new_n112), .c(new_n115), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(new_n116), .b(new_n117), .c(new_n118), .o1(new_n123));
  oai112aa1n02x5               g028(.a(new_n111), .b(new_n120), .c(\b[7] ), .d(\a[8] ), .o1(new_n124));
  oai022aa1n02x5               g029(.a(new_n116), .b(new_n117), .c(\a[7] ), .d(\b[6] ), .o1(new_n125));
  oab012aa1n02x4               g030(.a(new_n109), .b(\a[5] ), .c(\b[4] ), .out0(new_n126));
  oai013aa1n03x5               g031(.a(new_n123), .b(new_n124), .c(new_n126), .d(new_n125), .o1(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n122), .d(new_n108), .o1(new_n129));
  tech160nm_fixnrc02aa1n04x5   g034(.a(\b[9] ), .b(\a[10] ), .out0(new_n130));
  xobna2aa1n03x5               g035(.a(new_n130), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  oai022aa1n02x5               g036(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n132));
  aob012aa1n02x5               g037(.a(new_n132), .b(\b[9] ), .c(\a[10] ), .out0(new_n133));
  aoai13aa1n04x5               g038(.a(new_n133), .b(new_n130), .c(new_n129), .d(new_n98), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nand02aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  aoi012aa1n02x5               g042(.a(new_n136), .b(new_n134), .c(new_n137), .o1(new_n138));
  norp02aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand02aa1d04x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  inv000aa1d42x5               g046(.a(new_n141), .o1(new_n142));
  aoi112aa1n02x5               g047(.a(new_n136), .b(new_n142), .c(new_n134), .d(new_n137), .o1(new_n143));
  oab012aa1n02x5               g048(.a(new_n143), .b(new_n138), .c(new_n141), .out0(\s[12] ));
  aoi012aa1n12x5               g049(.a(new_n127), .b(new_n122), .c(new_n108), .o1(new_n145));
  inv000aa1n06x5               g050(.a(new_n145), .o1(new_n146));
  nona23aa1d18x5               g051(.a(new_n140), .b(new_n137), .c(new_n136), .d(new_n139), .out0(new_n147));
  norb03aa1d15x5               g052(.a(new_n128), .b(new_n147), .c(new_n130), .out0(new_n148));
  ao0012aa1n03x7               g053(.a(new_n139), .b(new_n136), .c(new_n140), .o(new_n149));
  oabi12aa1n06x5               g054(.a(new_n149), .b(new_n147), .c(new_n133), .out0(new_n150));
  nor042aa1n06x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(\b[12] ), .b(\a[13] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  aoai13aa1n02x5               g058(.a(new_n153), .b(new_n150), .c(new_n146), .d(new_n148), .o1(new_n154));
  aoi112aa1n02x5               g059(.a(new_n153), .b(new_n150), .c(new_n146), .d(new_n148), .o1(new_n155));
  norb02aa1n02x5               g060(.a(new_n154), .b(new_n155), .out0(\s[13] ));
  inv000aa1n06x5               g061(.a(new_n151), .o1(new_n157));
  xorc02aa1n02x5               g062(.a(\a[14] ), .b(\b[13] ), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n154), .c(new_n157), .out0(\s[14] ));
  xnrc02aa1n02x5               g064(.a(\b[13] ), .b(\a[14] ), .out0(new_n160));
  nano22aa1n03x7               g065(.a(new_n160), .b(new_n157), .c(new_n152), .out0(new_n161));
  aoai13aa1n06x5               g066(.a(new_n161), .b(new_n150), .c(new_n146), .d(new_n148), .o1(new_n162));
  oaoi03aa1n09x5               g067(.a(\a[14] ), .b(\b[13] ), .c(new_n157), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  xorc02aa1n12x5               g069(.a(\a[15] ), .b(\b[14] ), .out0(new_n165));
  xnbna2aa1n03x5               g070(.a(new_n165), .b(new_n162), .c(new_n164), .out0(\s[15] ));
  aob012aa1n02x5               g071(.a(new_n165), .b(new_n162), .c(new_n164), .out0(new_n167));
  nor042aa1n03x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n165), .o1(new_n170));
  aoai13aa1n02x5               g075(.a(new_n169), .b(new_n170), .c(new_n162), .d(new_n164), .o1(new_n171));
  xorc02aa1n02x5               g076(.a(\a[16] ), .b(\b[15] ), .out0(new_n172));
  norp02aa1n02x5               g077(.a(new_n172), .b(new_n168), .o1(new_n173));
  aoi022aa1n02x5               g078(.a(new_n171), .b(new_n172), .c(new_n167), .d(new_n173), .o1(\s[16] ));
  nand22aa1n04x5               g079(.a(new_n172), .b(new_n165), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(new_n158), .b(new_n153), .o1(new_n176));
  nona22aa1n09x5               g081(.a(new_n148), .b(new_n176), .c(new_n175), .out0(new_n177));
  aoi012aa1n06x5               g082(.a(new_n163), .b(new_n150), .c(new_n161), .o1(new_n178));
  oao003aa1n02x5               g083(.a(\a[16] ), .b(\b[15] ), .c(new_n169), .carry(new_n179));
  oai122aa1n12x5               g084(.a(new_n179), .b(new_n178), .c(new_n175), .d(new_n177), .e(new_n145), .o1(new_n180));
  xorb03aa1n02x5               g085(.a(new_n180), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g086(.a(\a[17] ), .o1(new_n182));
  nanb02aa1n03x5               g087(.a(\b[16] ), .b(new_n182), .out0(new_n183));
  nor042aa1n06x5               g088(.a(new_n145), .b(new_n177), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n185));
  nano23aa1n06x5               g090(.a(new_n136), .b(new_n139), .c(new_n140), .d(new_n137), .out0(new_n186));
  aoai13aa1n04x5               g091(.a(new_n161), .b(new_n149), .c(new_n186), .d(new_n185), .o1(new_n187));
  aoai13aa1n04x5               g092(.a(new_n179), .b(new_n175), .c(new_n187), .d(new_n164), .o1(new_n188));
  xorc02aa1n02x5               g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  oai012aa1n02x5               g094(.a(new_n189), .b(new_n188), .c(new_n184), .o1(new_n190));
  xorc02aa1n02x5               g095(.a(\a[18] ), .b(\b[17] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n190), .c(new_n183), .out0(\s[18] ));
  inv000aa1d42x5               g097(.a(\a[18] ), .o1(new_n193));
  xroi22aa1d04x5               g098(.a(new_n182), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n194));
  oaih12aa1n02x5               g099(.a(new_n194), .b(new_n188), .c(new_n184), .o1(new_n195));
  oai022aa1n03x5               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oaib12aa1n09x5               g101(.a(new_n196), .b(new_n193), .c(\b[17] ), .out0(new_n197));
  nor002aa1n20x5               g102(.a(\b[18] ), .b(\a[19] ), .o1(new_n198));
  nand02aa1d08x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n199), .b(new_n198), .out0(new_n200));
  xnbna2aa1n03x5               g105(.a(new_n200), .b(new_n195), .c(new_n197), .out0(\s[19] ));
  xnrc02aa1n02x5               g106(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n12x5               g107(.a(\a[18] ), .b(\b[17] ), .c(new_n183), .o1(new_n203));
  aoai13aa1n03x5               g108(.a(new_n200), .b(new_n203), .c(new_n180), .d(new_n194), .o1(new_n204));
  inv000aa1d42x5               g109(.a(new_n198), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n200), .o1(new_n206));
  aoai13aa1n02x5               g111(.a(new_n205), .b(new_n206), .c(new_n195), .d(new_n197), .o1(new_n207));
  nor042aa1n04x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand22aa1n12x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoib12aa1n02x5               g115(.a(new_n198), .b(new_n209), .c(new_n208), .out0(new_n211));
  aoi022aa1n03x5               g116(.a(new_n207), .b(new_n210), .c(new_n204), .d(new_n211), .o1(\s[20] ));
  nona23aa1d18x5               g117(.a(new_n209), .b(new_n199), .c(new_n198), .d(new_n208), .out0(new_n213));
  nano22aa1n03x7               g118(.a(new_n213), .b(new_n189), .c(new_n191), .out0(new_n214));
  oaih12aa1n02x5               g119(.a(new_n214), .b(new_n188), .c(new_n184), .o1(new_n215));
  aoi012aa1n12x5               g120(.a(new_n208), .b(new_n198), .c(new_n209), .o1(new_n216));
  oai012aa1d24x5               g121(.a(new_n216), .b(new_n213), .c(new_n197), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  xorc02aa1n02x5               g123(.a(\a[21] ), .b(\b[20] ), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n215), .c(new_n218), .out0(\s[21] ));
  aoai13aa1n03x5               g125(.a(new_n219), .b(new_n217), .c(new_n180), .d(new_n214), .o1(new_n221));
  nor002aa1d32x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n219), .o1(new_n224));
  aoai13aa1n02x5               g129(.a(new_n223), .b(new_n224), .c(new_n215), .d(new_n218), .o1(new_n225));
  xorc02aa1n02x5               g130(.a(\a[22] ), .b(\b[21] ), .out0(new_n226));
  norp02aa1n02x5               g131(.a(new_n226), .b(new_n222), .o1(new_n227));
  aoi022aa1n03x5               g132(.a(new_n225), .b(new_n226), .c(new_n221), .d(new_n227), .o1(\s[22] ));
  nano23aa1n06x5               g133(.a(new_n198), .b(new_n208), .c(new_n209), .d(new_n199), .out0(new_n229));
  nanp02aa1n02x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  tech160nm_fixnrc02aa1n05x5   g135(.a(\b[21] ), .b(\a[22] ), .out0(new_n231));
  nano22aa1n12x5               g136(.a(new_n231), .b(new_n223), .c(new_n230), .out0(new_n232));
  and003aa1n02x5               g137(.a(new_n194), .b(new_n232), .c(new_n229), .o(new_n233));
  oaih12aa1n02x5               g138(.a(new_n233), .b(new_n188), .c(new_n184), .o1(new_n234));
  oao003aa1n12x5               g139(.a(\a[22] ), .b(\b[21] ), .c(new_n223), .carry(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi012aa1d24x5               g141(.a(new_n236), .b(new_n217), .c(new_n232), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  xnbna2aa1n03x5               g143(.a(new_n238), .b(new_n234), .c(new_n237), .out0(\s[23] ));
  inv000aa1d42x5               g144(.a(new_n237), .o1(new_n240));
  aoai13aa1n02x7               g145(.a(new_n238), .b(new_n240), .c(new_n180), .d(new_n233), .o1(new_n241));
  nor042aa1n06x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  inv000aa1d42x5               g148(.a(new_n238), .o1(new_n244));
  aoai13aa1n02x5               g149(.a(new_n243), .b(new_n244), .c(new_n234), .d(new_n237), .o1(new_n245));
  tech160nm_fixorc02aa1n02p5x5 g150(.a(\a[24] ), .b(\b[23] ), .out0(new_n246));
  norp02aa1n02x5               g151(.a(new_n246), .b(new_n242), .o1(new_n247));
  aoi022aa1n03x5               g152(.a(new_n245), .b(new_n246), .c(new_n241), .d(new_n247), .o1(\s[24] ));
  and002aa1n12x5               g153(.a(new_n246), .b(new_n238), .o(new_n249));
  inv020aa1n04x5               g154(.a(new_n249), .o1(new_n250));
  nano32aa1n02x4               g155(.a(new_n250), .b(new_n194), .c(new_n229), .d(new_n232), .out0(new_n251));
  oaih12aa1n02x5               g156(.a(new_n251), .b(new_n188), .c(new_n184), .o1(new_n252));
  inv040aa1n02x5               g157(.a(new_n216), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n232), .b(new_n253), .c(new_n229), .d(new_n203), .o1(new_n254));
  oao003aa1n02x5               g159(.a(\a[24] ), .b(\b[23] ), .c(new_n243), .carry(new_n255));
  aoai13aa1n12x5               g160(.a(new_n255), .b(new_n250), .c(new_n254), .d(new_n235), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n256), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  xnbna2aa1n03x5               g163(.a(new_n258), .b(new_n252), .c(new_n257), .out0(\s[25] ));
  aoai13aa1n03x5               g164(.a(new_n258), .b(new_n256), .c(new_n180), .d(new_n251), .o1(new_n260));
  nor042aa1n03x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n258), .o1(new_n263));
  aoai13aa1n02x5               g168(.a(new_n262), .b(new_n263), .c(new_n252), .d(new_n257), .o1(new_n264));
  xorc02aa1n02x5               g169(.a(\a[26] ), .b(\b[25] ), .out0(new_n265));
  norp02aa1n02x5               g170(.a(new_n265), .b(new_n261), .o1(new_n266));
  aoi022aa1n03x5               g171(.a(new_n264), .b(new_n265), .c(new_n260), .d(new_n266), .o1(\s[26] ));
  and002aa1n02x5               g172(.a(new_n265), .b(new_n258), .o(new_n268));
  inv000aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  nano32aa1n03x7               g174(.a(new_n269), .b(new_n214), .c(new_n232), .d(new_n249), .out0(new_n270));
  oai012aa1n09x5               g175(.a(new_n270), .b(new_n188), .c(new_n184), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[26] ), .b(\b[25] ), .c(new_n262), .carry(new_n272));
  aobi12aa1n12x5               g177(.a(new_n272), .b(new_n256), .c(new_n268), .out0(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n271), .out0(\s[27] ));
  aoai13aa1n03x5               g180(.a(new_n249), .b(new_n236), .c(new_n217), .d(new_n232), .o1(new_n276));
  aoai13aa1n04x5               g181(.a(new_n272), .b(new_n269), .c(new_n276), .d(new_n255), .o1(new_n277));
  aoai13aa1n02x7               g182(.a(new_n274), .b(new_n277), .c(new_n180), .d(new_n270), .o1(new_n278));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  inv000aa1n03x5               g184(.a(new_n279), .o1(new_n280));
  inv000aa1n02x5               g185(.a(new_n274), .o1(new_n281));
  aoai13aa1n02x5               g186(.a(new_n280), .b(new_n281), .c(new_n273), .d(new_n271), .o1(new_n282));
  tech160nm_fixorc02aa1n03p5x5 g187(.a(\a[28] ), .b(\b[27] ), .out0(new_n283));
  norp02aa1n02x5               g188(.a(new_n283), .b(new_n279), .o1(new_n284));
  aoi022aa1n03x5               g189(.a(new_n282), .b(new_n283), .c(new_n278), .d(new_n284), .o1(\s[28] ));
  and002aa1n02x5               g190(.a(new_n283), .b(new_n274), .o(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n277), .c(new_n180), .d(new_n270), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n286), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n280), .carry(new_n289));
  aoai13aa1n02x7               g194(.a(new_n289), .b(new_n288), .c(new_n273), .d(new_n271), .o1(new_n290));
  tech160nm_fixorc02aa1n03p5x5 g195(.a(\a[29] ), .b(\b[28] ), .out0(new_n291));
  norb02aa1n02x5               g196(.a(new_n289), .b(new_n291), .out0(new_n292));
  aoi022aa1n03x5               g197(.a(new_n290), .b(new_n291), .c(new_n287), .d(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n105), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g199(.a(new_n281), .b(new_n283), .c(new_n291), .out0(new_n295));
  aoai13aa1n02x7               g200(.a(new_n295), .b(new_n277), .c(new_n180), .d(new_n270), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n295), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n297), .c(new_n273), .d(new_n271), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[30] ), .b(\b[29] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n298), .b(new_n300), .out0(new_n301));
  aoi022aa1n03x5               g206(.a(new_n299), .b(new_n300), .c(new_n296), .d(new_n301), .o1(\s[30] ));
  xorc02aa1n02x5               g207(.a(\a[31] ), .b(\b[30] ), .out0(new_n303));
  nano32aa1n03x7               g208(.a(new_n281), .b(new_n300), .c(new_n283), .d(new_n291), .out0(new_n304));
  aoai13aa1n02x5               g209(.a(new_n304), .b(new_n277), .c(new_n180), .d(new_n270), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n304), .o1(new_n306));
  oao003aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n306), .c(new_n273), .d(new_n271), .o1(new_n308));
  and002aa1n02x5               g213(.a(\b[29] ), .b(\a[30] ), .o(new_n309));
  oabi12aa1n02x5               g214(.a(new_n303), .b(\a[30] ), .c(\b[29] ), .out0(new_n310));
  oab012aa1n02x4               g215(.a(new_n310), .b(new_n298), .c(new_n309), .out0(new_n311));
  aoi022aa1n03x5               g216(.a(new_n308), .b(new_n303), .c(new_n305), .d(new_n311), .o1(\s[31] ));
  xorb03aa1n02x5               g217(.a(new_n107), .b(\b[2] ), .c(new_n99), .out0(\s[3] ));
  norp02aa1n02x5               g218(.a(new_n103), .b(new_n107), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[4] ), .b(\b[3] ), .out0(new_n315));
  aoi012aa1n02x5               g220(.a(new_n315), .b(new_n99), .c(new_n101), .o1(new_n316));
  aboi22aa1n03x5               g221(.a(new_n314), .b(new_n316), .c(new_n108), .d(new_n315), .out0(\s[4] ));
  xnrc02aa1n02x5               g222(.a(\b[4] ), .b(\a[5] ), .out0(new_n318));
  oaib12aa1n02x5               g223(.a(new_n108), .b(new_n100), .c(\b[3] ), .out0(new_n319));
  aboi22aa1n03x5               g224(.a(new_n115), .b(new_n108), .c(new_n319), .d(new_n318), .out0(\s[5] ));
  obai22aa1n02x7               g225(.a(new_n108), .b(new_n115), .c(\a[5] ), .d(\b[4] ), .out0(new_n321));
  xorb03aa1n02x5               g226(.a(new_n321), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norb02aa1n02x5               g227(.a(new_n120), .b(new_n118), .out0(new_n323));
  aoai13aa1n02x5               g228(.a(new_n323), .b(new_n109), .c(new_n321), .d(new_n111), .o1(new_n324));
  aoi112aa1n02x5               g229(.a(new_n323), .b(new_n109), .c(new_n321), .d(new_n111), .o1(new_n325));
  norb02aa1n02x5               g230(.a(new_n324), .b(new_n325), .out0(\s[7] ));
  xorc02aa1n02x5               g231(.a(\a[8] ), .b(\b[7] ), .out0(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n327), .b(new_n324), .c(new_n119), .out0(\s[8] ));
  xorb03aa1n02x5               g233(.a(new_n145), .b(\b[8] ), .c(new_n97), .out0(\s[9] ));
endmodule


