// Benchmark "adder" written by ABC on Thu Jul 18 02:35:06 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n185, new_n186, new_n187, new_n188,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n317,
    new_n320, new_n321, new_n322, new_n324, new_n325, new_n327, new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n20x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand02aa1d16x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[7] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[6] ), .o1(new_n103));
  nand42aa1n06x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  nor002aa1d32x5               g009(.a(\b[7] ), .b(\a[8] ), .o1(new_n105));
  aoai13aa1n02x5               g010(.a(new_n104), .b(new_n105), .c(new_n103), .d(new_n102), .o1(new_n106));
  xnrc02aa1n12x5               g011(.a(\b[6] ), .b(\a[7] ), .out0(new_n107));
  nand42aa1n16x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  inv000aa1n02x5               g013(.a(new_n108), .o1(new_n109));
  inv040aa1n02x5               g014(.a(new_n105), .o1(new_n110));
  nor042aa1n12x5               g015(.a(\b[5] ), .b(\a[6] ), .o1(new_n111));
  nor042aa1d18x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  oai112aa1n04x5               g017(.a(new_n110), .b(new_n104), .c(new_n111), .d(new_n112), .o1(new_n113));
  oai013aa1n03x5               g018(.a(new_n106), .b(new_n113), .c(new_n107), .d(new_n109), .o1(new_n114));
  nand42aa1n02x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  nand02aa1d06x5               g020(.a(\b[0] ), .b(\a[1] ), .o1(new_n116));
  nor042aa1n03x5               g021(.a(\b[1] ), .b(\a[2] ), .o1(new_n117));
  oai012aa1d24x5               g022(.a(new_n115), .b(new_n117), .c(new_n116), .o1(new_n118));
  nor022aa1n08x5               g023(.a(\b[2] ), .b(\a[3] ), .o1(new_n119));
  nand42aa1n02x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  nor002aa1n20x5               g025(.a(\b[3] ), .b(\a[4] ), .o1(new_n121));
  nand22aa1n12x5               g026(.a(\b[3] ), .b(\a[4] ), .o1(new_n122));
  nona23aa1n09x5               g027(.a(new_n122), .b(new_n120), .c(new_n119), .d(new_n121), .out0(new_n123));
  ao0012aa1n03x7               g028(.a(new_n121), .b(new_n119), .c(new_n122), .o(new_n124));
  oabi12aa1n18x5               g029(.a(new_n124), .b(new_n123), .c(new_n118), .out0(new_n125));
  nanb02aa1n18x5               g030(.a(new_n111), .b(new_n108), .out0(new_n126));
  nand02aa1n03x5               g031(.a(\b[4] ), .b(\a[5] ), .o1(new_n127));
  nona23aa1n02x4               g032(.a(new_n104), .b(new_n127), .c(new_n112), .d(new_n105), .out0(new_n128));
  nor043aa1n03x5               g033(.a(new_n128), .b(new_n126), .c(new_n107), .o1(new_n129));
  nanp02aa1n09x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n100), .out0(new_n131));
  aoai13aa1n03x5               g036(.a(new_n131), .b(new_n114), .c(new_n125), .d(new_n129), .o1(new_n132));
  xobna2aa1n03x5               g037(.a(new_n99), .b(new_n132), .c(new_n101), .out0(\s[10] ));
  nor002aa1d32x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand02aa1n10x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  oai022aa1n02x5               g041(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  nanp02aa1n03x5               g043(.a(new_n132), .b(new_n138), .o1(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n136), .b(new_n139), .c(new_n98), .out0(\s[11] ));
  nanb03aa1n09x5               g045(.a(new_n134), .b(new_n135), .c(new_n98), .out0(new_n141));
  aoib12aa1n06x5               g046(.a(new_n134), .b(new_n139), .c(new_n141), .out0(new_n142));
  xnrb03aa1n03x5               g047(.a(new_n142), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n12x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand02aa1n16x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nano23aa1n09x5               g050(.a(new_n97), .b(new_n144), .c(new_n145), .d(new_n98), .out0(new_n146));
  nano23aa1n09x5               g051(.a(new_n100), .b(new_n134), .c(new_n135), .d(new_n130), .out0(new_n147));
  nand22aa1n09x5               g052(.a(new_n147), .b(new_n146), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n03x5               g054(.a(new_n149), .b(new_n114), .c(new_n125), .d(new_n129), .o1(new_n150));
  inv030aa1n03x5               g055(.a(new_n144), .o1(new_n151));
  oai112aa1n06x5               g056(.a(new_n151), .b(new_n145), .c(new_n100), .d(new_n97), .o1(new_n152));
  tech160nm_fiaoi012aa1n03p5x5 g057(.a(new_n144), .b(new_n134), .c(new_n145), .o1(new_n153));
  oai012aa1n12x5               g058(.a(new_n153), .b(new_n152), .c(new_n141), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(new_n150), .b(new_n155), .o1(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1n03x5               g062(.a(\b[12] ), .b(\a[13] ), .o1(new_n158));
  nand42aa1n08x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  aoi012aa1n02x5               g064(.a(new_n158), .b(new_n156), .c(new_n159), .o1(new_n160));
  xnrb03aa1n02x5               g065(.a(new_n160), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nand42aa1n06x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  tech160nm_fiao0012aa1n04x5   g068(.a(new_n162), .b(new_n158), .c(new_n163), .o(new_n164));
  inv000aa1d42x5               g069(.a(new_n164), .o1(new_n165));
  nona23aa1n09x5               g070(.a(new_n163), .b(new_n159), .c(new_n158), .d(new_n162), .out0(new_n166));
  aoai13aa1n04x5               g071(.a(new_n165), .b(new_n166), .c(new_n150), .d(new_n155), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n03x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nand22aa1n06x5               g074(.a(\b[14] ), .b(\a[15] ), .o1(new_n170));
  nor042aa1n02x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nand02aa1n06x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  aoai13aa1n02x5               g078(.a(new_n173), .b(new_n169), .c(new_n167), .d(new_n170), .o1(new_n174));
  aoi112aa1n02x5               g079(.a(new_n173), .b(new_n169), .c(new_n167), .d(new_n170), .o1(new_n175));
  norb02aa1n03x4               g080(.a(new_n174), .b(new_n175), .out0(\s[16] ));
  nano23aa1n03x7               g081(.a(new_n158), .b(new_n162), .c(new_n163), .d(new_n159), .out0(new_n177));
  nano23aa1n06x5               g082(.a(new_n169), .b(new_n171), .c(new_n172), .d(new_n170), .out0(new_n178));
  nano22aa1n06x5               g083(.a(new_n148), .b(new_n177), .c(new_n178), .out0(new_n179));
  aoai13aa1n12x5               g084(.a(new_n179), .b(new_n114), .c(new_n125), .d(new_n129), .o1(new_n180));
  aoai13aa1n04x5               g085(.a(new_n178), .b(new_n164), .c(new_n154), .d(new_n177), .o1(new_n181));
  tech160nm_fiaoi012aa1n04x5   g086(.a(new_n171), .b(new_n169), .c(new_n172), .o1(new_n182));
  nand23aa1n06x5               g087(.a(new_n180), .b(new_n181), .c(new_n182), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g089(.a(\a[18] ), .o1(new_n185));
  inv030aa1d32x5               g090(.a(\a[17] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[16] ), .o1(new_n187));
  oaoi03aa1n03x5               g092(.a(new_n186), .b(new_n187), .c(new_n183), .o1(new_n188));
  xorb03aa1n02x5               g093(.a(new_n188), .b(\b[17] ), .c(new_n185), .out0(\s[18] ));
  oaoi13aa1n03x5               g094(.a(new_n166), .b(new_n153), .c(new_n152), .d(new_n141), .o1(new_n190));
  inv000aa1n02x5               g095(.a(new_n182), .o1(new_n191));
  oaoi13aa1n09x5               g096(.a(new_n191), .b(new_n178), .c(new_n190), .d(new_n164), .o1(new_n192));
  xroi22aa1d06x4               g097(.a(new_n186), .b(\b[16] ), .c(new_n185), .d(\b[17] ), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[17] ), .o1(new_n195));
  oai022aa1d18x5               g100(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n196));
  oa0012aa1n02x5               g101(.a(new_n196), .b(new_n195), .c(new_n185), .o(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  aoai13aa1n06x5               g103(.a(new_n198), .b(new_n194), .c(new_n192), .d(new_n180), .o1(new_n199));
  xorb03aa1n02x5               g104(.a(new_n199), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n16x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  nand02aa1d06x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  nanb02aa1n12x5               g109(.a(new_n202), .b(new_n204), .out0(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n206), .b(new_n197), .c(new_n183), .d(new_n193), .o1(new_n207));
  nor002aa1n12x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  nand02aa1d08x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanb02aa1d30x5               g114(.a(new_n208), .b(new_n209), .out0(new_n210));
  tech160nm_fiaoi012aa1n02p5x5 g115(.a(new_n210), .b(new_n207), .c(new_n203), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n210), .o1(new_n212));
  aoi112aa1n03x4               g117(.a(new_n202), .b(new_n212), .c(new_n199), .d(new_n204), .o1(new_n213));
  nor002aa1n02x5               g118(.a(new_n211), .b(new_n213), .o1(\s[20] ));
  nona22aa1n12x5               g119(.a(new_n193), .b(new_n205), .c(new_n210), .out0(new_n215));
  oai112aa1n06x5               g120(.a(new_n196), .b(new_n204), .c(new_n195), .d(new_n185), .o1(new_n216));
  nona22aa1n09x5               g121(.a(new_n216), .b(new_n208), .c(new_n202), .out0(new_n217));
  nand02aa1d12x5               g122(.a(new_n217), .b(new_n209), .o1(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n215), .c(new_n192), .d(new_n180), .o1(new_n219));
  xorb03aa1n02x5               g124(.a(new_n219), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n09x5               g125(.a(\b[20] ), .b(\a[21] ), .o1(new_n221));
  inv000aa1n06x5               g126(.a(new_n221), .o1(new_n222));
  inv000aa1n02x5               g127(.a(new_n215), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n218), .o1(new_n224));
  nand02aa1d08x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  norb02aa1n06x5               g130(.a(new_n225), .b(new_n221), .out0(new_n226));
  aoai13aa1n06x5               g131(.a(new_n226), .b(new_n224), .c(new_n183), .d(new_n223), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  tech160nm_fiaoi012aa1n03p5x5 g133(.a(new_n228), .b(new_n227), .c(new_n222), .o1(new_n229));
  xorc02aa1n02x5               g134(.a(\a[22] ), .b(\b[21] ), .out0(new_n230));
  aoi112aa1n03x4               g135(.a(new_n221), .b(new_n230), .c(new_n219), .d(new_n226), .o1(new_n231));
  nor042aa1n03x5               g136(.a(new_n229), .b(new_n231), .o1(\s[22] ));
  xorc02aa1n02x5               g137(.a(\a[23] ), .b(\b[22] ), .out0(new_n233));
  nand42aa1n02x5               g138(.a(new_n230), .b(new_n226), .o1(new_n234));
  nona22aa1n03x5               g139(.a(new_n183), .b(new_n215), .c(new_n234), .out0(new_n235));
  nano22aa1n02x4               g140(.a(new_n228), .b(new_n222), .c(new_n225), .out0(new_n236));
  xnrc02aa1n03x5               g141(.a(\b[22] ), .b(\a[23] ), .out0(new_n237));
  oaoi03aa1n03x5               g142(.a(\a[22] ), .b(\b[21] ), .c(new_n222), .o1(new_n238));
  aoi113aa1n02x5               g143(.a(new_n238), .b(new_n237), .c(new_n217), .d(new_n236), .e(new_n209), .o1(new_n239));
  nand42aa1n03x5               g144(.a(new_n235), .b(new_n239), .o1(new_n240));
  oabi12aa1n02x5               g145(.a(new_n238), .b(new_n218), .c(new_n234), .out0(new_n241));
  aoi013aa1n02x4               g146(.a(new_n241), .b(new_n183), .c(new_n223), .d(new_n236), .o1(new_n242));
  oaih12aa1n02x5               g147(.a(new_n240), .b(new_n242), .c(new_n233), .o1(\s[23] ));
  and002aa1n02x5               g148(.a(\b[22] ), .b(\a[23] ), .o(new_n244));
  xorc02aa1n12x5               g149(.a(\a[24] ), .b(\b[23] ), .out0(new_n245));
  aoai13aa1n02x7               g150(.a(new_n245), .b(new_n244), .c(new_n235), .d(new_n239), .o1(new_n246));
  nona22aa1n03x5               g151(.a(new_n240), .b(new_n245), .c(new_n244), .out0(new_n247));
  nanp02aa1n03x5               g152(.a(new_n247), .b(new_n246), .o1(\s[24] ));
  nona23aa1d18x5               g153(.a(new_n226), .b(new_n245), .c(new_n237), .d(new_n228), .out0(new_n249));
  nor042aa1n06x5               g154(.a(new_n215), .b(new_n249), .o1(new_n250));
  inv020aa1n03x5               g155(.a(new_n250), .o1(new_n251));
  orn002aa1n02x5               g156(.a(\a[23] ), .b(\b[22] ), .o(new_n252));
  oaoi03aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .c(new_n252), .o1(new_n253));
  aoi013aa1n06x4               g158(.a(new_n253), .b(new_n238), .c(new_n245), .d(new_n233), .o1(new_n254));
  oai012aa1n12x5               g159(.a(new_n254), .b(new_n218), .c(new_n249), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  aoai13aa1n04x5               g161(.a(new_n256), .b(new_n251), .c(new_n192), .d(new_n180), .o1(new_n257));
  xorb03aa1n02x5               g162(.a(new_n257), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g163(.a(\b[24] ), .b(\a[25] ), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n259), .o1(new_n260));
  tech160nm_fixorc02aa1n03p5x5 g165(.a(\a[25] ), .b(\b[24] ), .out0(new_n261));
  aoai13aa1n06x5               g166(.a(new_n261), .b(new_n255), .c(new_n183), .d(new_n250), .o1(new_n262));
  xorc02aa1n12x5               g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  tech160nm_fiaoi012aa1n03p5x5 g169(.a(new_n264), .b(new_n262), .c(new_n260), .o1(new_n265));
  aoi112aa1n03x4               g170(.a(new_n259), .b(new_n263), .c(new_n257), .d(new_n261), .o1(new_n266));
  nor042aa1n03x5               g171(.a(new_n265), .b(new_n266), .o1(\s[26] ));
  and002aa1n03x5               g172(.a(new_n263), .b(new_n261), .o(new_n268));
  inv040aa1n02x5               g173(.a(new_n268), .o1(new_n269));
  nor043aa1d12x5               g174(.a(new_n269), .b(new_n215), .c(new_n249), .o1(new_n270));
  inv020aa1n03x5               g175(.a(new_n270), .o1(new_n271));
  oao003aa1n02x5               g176(.a(\a[26] ), .b(\b[25] ), .c(new_n260), .carry(new_n272));
  aobi12aa1n06x5               g177(.a(new_n272), .b(new_n255), .c(new_n268), .out0(new_n273));
  aoai13aa1n12x5               g178(.a(new_n273), .b(new_n271), .c(new_n192), .d(new_n180), .o1(new_n274));
  xorb03aa1n03x5               g179(.a(new_n274), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  inv000aa1n06x5               g181(.a(new_n276), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[28] ), .b(\b[27] ), .out0(new_n278));
  inv000aa1d42x5               g183(.a(new_n278), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  nano22aa1n02x4               g185(.a(new_n234), .b(new_n233), .c(new_n245), .out0(new_n281));
  nanp03aa1n02x5               g186(.a(new_n281), .b(new_n209), .c(new_n217), .o1(new_n282));
  aoai13aa1n06x5               g187(.a(new_n272), .b(new_n269), .c(new_n282), .d(new_n254), .o1(new_n283));
  aoai13aa1n03x5               g188(.a(new_n280), .b(new_n283), .c(new_n183), .d(new_n270), .o1(new_n284));
  tech160nm_fiaoi012aa1n03p5x5 g189(.a(new_n279), .b(new_n284), .c(new_n277), .o1(new_n285));
  aoi112aa1n03x4               g190(.a(new_n278), .b(new_n276), .c(new_n274), .d(new_n280), .o1(new_n286));
  nor002aa1n02x5               g191(.a(new_n285), .b(new_n286), .o1(\s[28] ));
  nano22aa1n02x4               g192(.a(new_n279), .b(new_n277), .c(new_n280), .out0(new_n288));
  aoai13aa1n03x5               g193(.a(new_n288), .b(new_n283), .c(new_n183), .d(new_n270), .o1(new_n289));
  oao003aa1n12x5               g194(.a(\a[28] ), .b(\b[27] ), .c(new_n277), .carry(new_n290));
  xorc02aa1n12x5               g195(.a(\a[29] ), .b(\b[28] ), .out0(new_n291));
  inv000aa1d42x5               g196(.a(new_n291), .o1(new_n292));
  tech160nm_fiaoi012aa1n03p5x5 g197(.a(new_n292), .b(new_n289), .c(new_n290), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n290), .o1(new_n294));
  aoi112aa1n03x4               g199(.a(new_n291), .b(new_n294), .c(new_n274), .d(new_n288), .o1(new_n295));
  nor002aa1n02x5               g200(.a(new_n293), .b(new_n295), .o1(\s[29] ));
  xorb03aa1n02x5               g201(.a(new_n116), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g202(.a(new_n292), .b(new_n278), .c(new_n280), .d(new_n277), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n298), .b(new_n283), .c(new_n183), .d(new_n270), .o1(new_n299));
  oao003aa1n12x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n290), .carry(new_n300));
  xorc02aa1n12x5               g205(.a(\a[30] ), .b(\b[29] ), .out0(new_n301));
  inv000aa1d42x5               g206(.a(new_n301), .o1(new_n302));
  tech160nm_fiaoi012aa1n03p5x5 g207(.a(new_n302), .b(new_n299), .c(new_n300), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n300), .o1(new_n304));
  aoi112aa1n03x4               g209(.a(new_n301), .b(new_n304), .c(new_n274), .d(new_n298), .o1(new_n305));
  nor002aa1n02x5               g210(.a(new_n303), .b(new_n305), .o1(\s[30] ));
  xnrc02aa1n02x5               g211(.a(\b[30] ), .b(\a[31] ), .out0(new_n307));
  and003aa1n02x5               g212(.a(new_n288), .b(new_n301), .c(new_n291), .o(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n283), .c(new_n183), .d(new_n270), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n300), .carry(new_n310));
  tech160nm_fiaoi012aa1n03p5x5 g215(.a(new_n307), .b(new_n309), .c(new_n310), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n307), .o1(new_n312));
  inv000aa1n02x5               g217(.a(new_n310), .o1(new_n313));
  aoi112aa1n03x4               g218(.a(new_n312), .b(new_n313), .c(new_n274), .d(new_n308), .o1(new_n314));
  norp02aa1n03x5               g219(.a(new_n311), .b(new_n314), .o1(\s[31] ));
  xnrb03aa1n02x5               g220(.a(new_n118), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g221(.a(\a[3] ), .b(\b[2] ), .c(new_n118), .o1(new_n317));
  xorb03aa1n02x5               g222(.a(new_n317), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g223(.a(new_n125), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g224(.a(new_n126), .o1(new_n320));
  oaoi13aa1n02x5               g225(.a(new_n320), .b(new_n127), .c(new_n125), .d(new_n112), .o1(new_n321));
  oai112aa1n04x5               g226(.a(new_n320), .b(new_n127), .c(new_n125), .d(new_n112), .o1(new_n322));
  norb02aa1n02x5               g227(.a(new_n322), .b(new_n321), .out0(\s[6] ));
  oaoi13aa1n02x5               g228(.a(new_n107), .b(new_n322), .c(\a[6] ), .d(\b[5] ), .o1(new_n324));
  oai112aa1n02x5               g229(.a(new_n322), .b(new_n107), .c(\b[5] ), .d(\a[6] ), .o1(new_n325));
  norb02aa1n02x5               g230(.a(new_n325), .b(new_n324), .out0(\s[7] ));
  tech160nm_fiaoi012aa1n05x5   g231(.a(new_n324), .b(new_n102), .c(new_n103), .o1(new_n327));
  xnbna2aa1n03x5               g232(.a(new_n327), .b(new_n104), .c(new_n110), .out0(\s[8] ));
  aoi112aa1n02x5               g233(.a(new_n131), .b(new_n114), .c(new_n125), .d(new_n129), .o1(new_n329));
  norb02aa1n02x5               g234(.a(new_n132), .b(new_n329), .out0(\s[9] ));
endmodule


