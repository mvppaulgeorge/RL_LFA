// Benchmark "adder" written by ABC on Thu Jul 18 03:13:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n313, new_n315, new_n316, new_n319,
    new_n320, new_n322, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n02x5               g001(.a(\a[9] ), .b(\b[8] ), .o(new_n97));
  inv000aa1d42x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oaoi03aa1n02x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n101));
  xnrc02aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .out0(new_n102));
  xnrc02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .out0(new_n103));
  orn002aa1n02x5               g008(.a(\a[4] ), .b(\b[3] ), .o(new_n104));
  aoi112aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .c(\a[4] ), .d(\b[3] ), .o1(new_n105));
  norb02aa1n03x5               g010(.a(new_n104), .b(new_n105), .out0(new_n106));
  oai013aa1n02x4               g011(.a(new_n106), .b(new_n101), .c(new_n102), .d(new_n103), .o1(new_n107));
  xorc02aa1n02x5               g012(.a(\a[6] ), .b(\b[5] ), .out0(new_n108));
  tech160nm_fixorc02aa1n02p5x5 g013(.a(\a[5] ), .b(\b[4] ), .out0(new_n109));
  xorc02aa1n12x5               g014(.a(\a[8] ), .b(\b[7] ), .out0(new_n110));
  nanp02aa1n02x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nor042aa1n12x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nanb02aa1n02x5               g017(.a(new_n112), .b(new_n111), .out0(new_n113));
  nano32aa1n02x4               g018(.a(new_n113), .b(new_n110), .c(new_n109), .d(new_n108), .out0(new_n114));
  nanp02aa1n02x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nano22aa1n09x5               g020(.a(new_n112), .b(new_n115), .c(new_n111), .out0(new_n116));
  oai022aa1n06x5               g021(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n117));
  inv000aa1d42x5               g022(.a(new_n112), .o1(new_n118));
  oaoi03aa1n02x5               g023(.a(\a[8] ), .b(\b[7] ), .c(new_n118), .o1(new_n119));
  aoi013aa1n09x5               g024(.a(new_n119), .b(new_n116), .c(new_n110), .d(new_n117), .o1(new_n120));
  inv000aa1d42x5               g025(.a(new_n120), .o1(new_n121));
  xnrc02aa1n12x5               g026(.a(\b[8] ), .b(\a[9] ), .out0(new_n122));
  inv000aa1d42x5               g027(.a(new_n122), .o1(new_n123));
  aoai13aa1n02x5               g028(.a(new_n123), .b(new_n121), .c(new_n114), .d(new_n107), .o1(new_n124));
  xorc02aa1n06x5               g029(.a(\a[10] ), .b(\b[9] ), .out0(new_n125));
  xnbna2aa1n03x5               g030(.a(new_n125), .b(new_n124), .c(new_n97), .out0(\s[10] ));
  oai022aa1n09x5               g031(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n127));
  nanb02aa1n03x5               g032(.a(new_n127), .b(new_n124), .out0(new_n128));
  nanp02aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanp02aa1n02x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  nor002aa1n03x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nanb03aa1n02x5               g036(.a(new_n131), .b(new_n129), .c(new_n130), .out0(new_n132));
  nanb02aa1n06x5               g037(.a(new_n131), .b(new_n130), .out0(new_n133));
  oao003aa1n02x5               g038(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n134));
  xorc02aa1n02x5               g039(.a(\a[4] ), .b(\b[3] ), .out0(new_n135));
  xorc02aa1n02x5               g040(.a(\a[3] ), .b(\b[2] ), .out0(new_n136));
  nanp03aa1n02x5               g041(.a(new_n134), .b(new_n135), .c(new_n136), .o1(new_n137));
  xnrc02aa1n02x5               g042(.a(\b[5] ), .b(\a[6] ), .out0(new_n138));
  nona23aa1n09x5               g043(.a(new_n109), .b(new_n110), .c(new_n138), .d(new_n113), .out0(new_n139));
  aoai13aa1n12x5               g044(.a(new_n120), .b(new_n139), .c(new_n137), .d(new_n106), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n129), .b(new_n127), .c(new_n140), .d(new_n123), .o1(new_n141));
  aboi22aa1n03x5               g046(.a(new_n132), .b(new_n128), .c(new_n141), .d(new_n133), .out0(\s[11] ));
  xorc02aa1n06x5               g047(.a(\a[12] ), .b(\b[11] ), .out0(new_n143));
  aoi113aa1n02x5               g048(.a(new_n143), .b(new_n131), .c(new_n128), .d(new_n130), .e(new_n129), .o1(new_n144));
  obai22aa1n02x7               g049(.a(new_n128), .b(new_n132), .c(\a[11] ), .d(\b[10] ), .out0(new_n145));
  aoi012aa1n02x5               g050(.a(new_n144), .b(new_n145), .c(new_n143), .o1(\s[12] ));
  nona23aa1d18x5               g051(.a(new_n143), .b(new_n125), .c(new_n122), .d(new_n133), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  aoi022aa1n02x5               g053(.a(\b[11] ), .b(\a[12] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n149));
  aoai13aa1n02x5               g054(.a(new_n149), .b(new_n131), .c(new_n127), .d(new_n129), .o1(new_n150));
  oai012aa1n02x5               g055(.a(new_n150), .b(\b[11] ), .c(\a[12] ), .o1(new_n151));
  xorc02aa1n02x5               g056(.a(\a[13] ), .b(\b[12] ), .out0(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n151), .c(new_n140), .d(new_n148), .o1(new_n153));
  aoi112aa1n02x5               g058(.a(new_n152), .b(new_n151), .c(new_n140), .d(new_n148), .o1(new_n154));
  norb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(\s[13] ));
  inv000aa1d42x5               g060(.a(\a[13] ), .o1(new_n156));
  inv000aa1d42x5               g061(.a(\b[12] ), .o1(new_n157));
  nand42aa1n03x5               g062(.a(new_n157), .b(new_n156), .o1(new_n158));
  norp02aa1n02x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nand42aa1n03x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  xnbna2aa1n03x5               g066(.a(new_n161), .b(new_n153), .c(new_n158), .out0(\s[14] ));
  nanp02aa1n02x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  nano32aa1n02x4               g068(.a(new_n159), .b(new_n158), .c(new_n160), .d(new_n163), .out0(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n151), .c(new_n140), .d(new_n148), .o1(new_n165));
  aoai13aa1n06x5               g070(.a(new_n160), .b(new_n159), .c(new_n156), .d(new_n157), .o1(new_n166));
  xorc02aa1n02x5               g071(.a(\a[15] ), .b(\b[14] ), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n165), .c(new_n166), .out0(\s[15] ));
  aob012aa1n02x5               g073(.a(new_n167), .b(new_n165), .c(new_n166), .out0(new_n169));
  norp02aa1n02x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(new_n172));
  orn002aa1n02x5               g077(.a(\a[15] ), .b(\b[14] ), .o(new_n173));
  norb02aa1n02x5               g078(.a(new_n173), .b(new_n172), .out0(new_n174));
  nand02aa1d06x5               g079(.a(\b[14] ), .b(\a[15] ), .o1(new_n175));
  inv000aa1d42x5               g080(.a(new_n175), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n173), .b(new_n176), .c(new_n165), .d(new_n166), .o1(new_n177));
  aoi022aa1n02x5               g082(.a(new_n177), .b(new_n172), .c(new_n169), .d(new_n174), .o1(\s[16] ));
  nano32aa1n02x4               g083(.a(new_n170), .b(new_n173), .c(new_n171), .d(new_n175), .out0(new_n179));
  nanp02aa1n02x5               g084(.a(new_n179), .b(new_n164), .o1(new_n180));
  nor042aa1n03x5               g085(.a(new_n147), .b(new_n180), .o1(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n121), .c(new_n114), .d(new_n107), .o1(new_n182));
  oai122aa1n02x7               g087(.a(new_n173), .b(new_n166), .c(new_n176), .d(\b[15] ), .e(\a[16] ), .o1(new_n183));
  nanp02aa1n02x5               g088(.a(new_n183), .b(new_n171), .o1(new_n184));
  oaib12aa1n06x5               g089(.a(new_n184), .b(new_n180), .c(new_n151), .out0(new_n185));
  nanb02aa1n06x5               g090(.a(new_n185), .b(new_n182), .out0(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g092(.a(\a[17] ), .o1(new_n188));
  nanb02aa1n02x5               g093(.a(\b[16] ), .b(new_n188), .out0(new_n189));
  xorc02aa1n02x5               g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  aoai13aa1n02x5               g095(.a(new_n190), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n191));
  xorc02aa1n02x5               g096(.a(\a[18] ), .b(\b[17] ), .out0(new_n192));
  xnbna2aa1n03x5               g097(.a(new_n192), .b(new_n191), .c(new_n189), .out0(\s[18] ));
  inv000aa1d42x5               g098(.a(\a[18] ), .o1(new_n194));
  xroi22aa1d04x5               g099(.a(new_n188), .b(\b[16] ), .c(new_n194), .d(\b[17] ), .out0(new_n195));
  aoai13aa1n02x5               g100(.a(new_n195), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n196));
  oai022aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oaib12aa1n02x5               g102(.a(new_n197), .b(new_n194), .c(\b[17] ), .out0(new_n198));
  nor042aa1n06x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nanp02aa1n02x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  inv000aa1d42x5               g106(.a(new_n201), .o1(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n196), .c(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n02x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n205));
  aoai13aa1n02x5               g110(.a(new_n202), .b(new_n205), .c(new_n186), .d(new_n195), .o1(new_n206));
  nor042aa1n02x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  nanp02aa1n02x5               g112(.a(\b[19] ), .b(\a[20] ), .o1(new_n208));
  norb02aa1n02x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  aoib12aa1n02x5               g114(.a(new_n199), .b(new_n208), .c(new_n207), .out0(new_n210));
  inv000aa1n02x5               g115(.a(new_n199), .o1(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n201), .c(new_n196), .d(new_n198), .o1(new_n212));
  aoi022aa1n02x5               g117(.a(new_n212), .b(new_n209), .c(new_n206), .d(new_n210), .o1(\s[20] ));
  nano23aa1n06x5               g118(.a(new_n199), .b(new_n207), .c(new_n208), .d(new_n200), .out0(new_n214));
  nand23aa1n04x5               g119(.a(new_n214), .b(new_n190), .c(new_n192), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n217));
  nona23aa1n09x5               g122(.a(new_n208), .b(new_n200), .c(new_n199), .d(new_n207), .out0(new_n218));
  oaoi03aa1n06x5               g123(.a(\a[20] ), .b(\b[19] ), .c(new_n211), .o1(new_n219));
  oabi12aa1n12x5               g124(.a(new_n219), .b(new_n218), .c(new_n198), .out0(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[20] ), .b(\a[21] ), .out0(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  xnbna2aa1n03x5               g128(.a(new_n223), .b(new_n217), .c(new_n221), .out0(\s[21] ));
  aoai13aa1n02x5               g129(.a(new_n223), .b(new_n220), .c(new_n186), .d(new_n216), .o1(new_n225));
  xnrc02aa1n02x5               g130(.a(\b[21] ), .b(\a[22] ), .out0(new_n226));
  nor042aa1n06x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  norb02aa1n02x5               g132(.a(new_n226), .b(new_n227), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n227), .o1(new_n229));
  aoai13aa1n02x5               g134(.a(new_n229), .b(new_n222), .c(new_n217), .d(new_n221), .o1(new_n230));
  aboi22aa1n03x5               g135(.a(new_n226), .b(new_n230), .c(new_n225), .d(new_n228), .out0(\s[22] ));
  nor042aa1n04x5               g136(.a(new_n226), .b(new_n222), .o1(new_n232));
  norb02aa1n02x5               g137(.a(new_n232), .b(new_n215), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n234));
  oao003aa1n02x5               g139(.a(\a[22] ), .b(\b[21] ), .c(new_n229), .carry(new_n235));
  inv000aa1n02x5               g140(.a(new_n235), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n220), .c(new_n232), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  aob012aa1n03x5               g143(.a(new_n238), .b(new_n234), .c(new_n237), .out0(new_n239));
  aoi112aa1n02x5               g144(.a(new_n238), .b(new_n236), .c(new_n220), .d(new_n232), .o1(new_n240));
  aobi12aa1n02x5               g145(.a(new_n239), .b(new_n240), .c(new_n234), .out0(\s[23] ));
  xorc02aa1n02x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  nor042aa1n03x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  norp02aa1n02x5               g148(.a(new_n242), .b(new_n243), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n243), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n238), .o1(new_n246));
  aoai13aa1n02x5               g151(.a(new_n245), .b(new_n246), .c(new_n234), .d(new_n237), .o1(new_n247));
  aoi022aa1n02x5               g152(.a(new_n247), .b(new_n242), .c(new_n239), .d(new_n244), .o1(\s[24] ));
  nano32aa1n02x4               g153(.a(new_n215), .b(new_n242), .c(new_n232), .d(new_n238), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n232), .b(new_n219), .c(new_n214), .d(new_n205), .o1(new_n251));
  and002aa1n06x5               g156(.a(new_n242), .b(new_n238), .o(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  oao003aa1n02x5               g158(.a(\a[24] ), .b(\b[23] ), .c(new_n245), .carry(new_n254));
  aoai13aa1n12x5               g159(.a(new_n254), .b(new_n253), .c(new_n251), .d(new_n235), .o1(new_n255));
  inv000aa1d42x5               g160(.a(new_n255), .o1(new_n256));
  xorc02aa1n12x5               g161(.a(\a[25] ), .b(\b[24] ), .out0(new_n257));
  xnbna2aa1n03x5               g162(.a(new_n257), .b(new_n250), .c(new_n256), .out0(\s[25] ));
  aoai13aa1n02x5               g163(.a(new_n257), .b(new_n255), .c(new_n186), .d(new_n249), .o1(new_n259));
  xorc02aa1n02x5               g164(.a(\a[26] ), .b(\b[25] ), .out0(new_n260));
  nor042aa1n03x5               g165(.a(\b[24] ), .b(\a[25] ), .o1(new_n261));
  norp02aa1n02x5               g166(.a(new_n260), .b(new_n261), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n261), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n257), .o1(new_n264));
  aoai13aa1n02x5               g169(.a(new_n263), .b(new_n264), .c(new_n250), .d(new_n256), .o1(new_n265));
  aoi022aa1n02x5               g170(.a(new_n265), .b(new_n260), .c(new_n259), .d(new_n262), .o1(\s[26] ));
  and002aa1n02x5               g171(.a(new_n260), .b(new_n257), .o(new_n267));
  inv000aa1n02x5               g172(.a(new_n267), .o1(new_n268));
  nano23aa1n06x5               g173(.a(new_n268), .b(new_n215), .c(new_n252), .d(new_n232), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n185), .c(new_n140), .d(new_n181), .o1(new_n270));
  oao003aa1n02x5               g175(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n271));
  inv000aa1d42x5               g176(.a(new_n271), .o1(new_n272));
  aoi012aa1n12x5               g177(.a(new_n272), .b(new_n255), .c(new_n267), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[27] ), .b(\b[26] ), .out0(new_n274));
  xnbna2aa1n03x5               g179(.a(new_n274), .b(new_n273), .c(new_n270), .out0(\s[27] ));
  aoai13aa1n06x5               g180(.a(new_n252), .b(new_n236), .c(new_n220), .d(new_n232), .o1(new_n276));
  aoai13aa1n04x5               g181(.a(new_n271), .b(new_n268), .c(new_n276), .d(new_n254), .o1(new_n277));
  aoai13aa1n02x5               g182(.a(new_n274), .b(new_n277), .c(new_n186), .d(new_n269), .o1(new_n278));
  tech160nm_fixorc02aa1n04x5   g183(.a(\a[28] ), .b(\b[27] ), .out0(new_n279));
  norp02aa1n02x5               g184(.a(\b[26] ), .b(\a[27] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(new_n281));
  inv000aa1n03x5               g186(.a(new_n280), .o1(new_n282));
  inv000aa1d42x5               g187(.a(new_n274), .o1(new_n283));
  aoai13aa1n02x5               g188(.a(new_n282), .b(new_n283), .c(new_n273), .d(new_n270), .o1(new_n284));
  aoi022aa1n02x5               g189(.a(new_n284), .b(new_n279), .c(new_n278), .d(new_n281), .o1(\s[28] ));
  and002aa1n02x5               g190(.a(new_n279), .b(new_n274), .o(new_n286));
  aoai13aa1n02x5               g191(.a(new_n286), .b(new_n277), .c(new_n186), .d(new_n269), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n286), .o1(new_n288));
  oao003aa1n02x5               g193(.a(\a[28] ), .b(\b[27] ), .c(new_n282), .carry(new_n289));
  aoai13aa1n02x5               g194(.a(new_n289), .b(new_n288), .c(new_n273), .d(new_n270), .o1(new_n290));
  xorc02aa1n02x5               g195(.a(\a[29] ), .b(\b[28] ), .out0(new_n291));
  norb02aa1n02x5               g196(.a(new_n289), .b(new_n291), .out0(new_n292));
  aoi022aa1n02x5               g197(.a(new_n290), .b(new_n291), .c(new_n287), .d(new_n292), .o1(\s[29] ));
  xorb03aa1n02x5               g198(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g199(.a(new_n283), .b(new_n279), .c(new_n291), .out0(new_n295));
  aoai13aa1n03x5               g200(.a(new_n295), .b(new_n277), .c(new_n186), .d(new_n269), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n295), .o1(new_n297));
  oao003aa1n02x5               g202(.a(\a[29] ), .b(\b[28] ), .c(new_n289), .carry(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n297), .c(new_n273), .d(new_n270), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[30] ), .b(\b[29] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n298), .b(new_n300), .out0(new_n301));
  aoi022aa1n02x5               g206(.a(new_n299), .b(new_n300), .c(new_n296), .d(new_n301), .o1(\s[30] ));
  nano32aa1n02x4               g207(.a(new_n283), .b(new_n300), .c(new_n279), .d(new_n291), .out0(new_n303));
  aoai13aa1n06x5               g208(.a(new_n303), .b(new_n277), .c(new_n186), .d(new_n269), .o1(new_n304));
  xorc02aa1n02x5               g209(.a(\a[31] ), .b(\b[30] ), .out0(new_n305));
  and002aa1n02x5               g210(.a(\b[29] ), .b(\a[30] ), .o(new_n306));
  oabi12aa1n02x5               g211(.a(new_n305), .b(\a[30] ), .c(\b[29] ), .out0(new_n307));
  oab012aa1n02x4               g212(.a(new_n307), .b(new_n298), .c(new_n306), .out0(new_n308));
  inv000aa1n02x5               g213(.a(new_n303), .o1(new_n309));
  oao003aa1n02x5               g214(.a(\a[30] ), .b(\b[29] ), .c(new_n298), .carry(new_n310));
  aoai13aa1n02x5               g215(.a(new_n310), .b(new_n309), .c(new_n273), .d(new_n270), .o1(new_n311));
  aoi022aa1n02x5               g216(.a(new_n311), .b(new_n305), .c(new_n304), .d(new_n308), .o1(\s[31] ));
  inv000aa1d42x5               g217(.a(\a[3] ), .o1(new_n313));
  xorb03aa1n02x5               g218(.a(new_n101), .b(\b[2] ), .c(new_n313), .out0(\s[3] ));
  nanp02aa1n02x5               g219(.a(new_n134), .b(new_n136), .o1(new_n315));
  aoib12aa1n02x5               g220(.a(new_n135), .b(new_n313), .c(\b[2] ), .out0(new_n316));
  aoi022aa1n02x5               g221(.a(new_n107), .b(new_n104), .c(new_n316), .d(new_n315), .o1(\s[4] ));
  xnbna2aa1n03x5               g222(.a(new_n109), .b(new_n137), .c(new_n106), .out0(\s[5] ));
  norp02aa1n02x5               g223(.a(\b[4] ), .b(\a[5] ), .o1(new_n319));
  aoi012aa1n02x5               g224(.a(new_n319), .b(new_n107), .c(new_n109), .o1(new_n320));
  xnrc02aa1n02x5               g225(.a(new_n320), .b(new_n108), .out0(\s[6] ));
  nanp02aa1n02x5               g226(.a(new_n320), .b(new_n108), .o1(new_n322));
  xnbna2aa1n03x5               g227(.a(new_n113), .b(new_n322), .c(new_n115), .out0(\s[7] ));
  nanp02aa1n02x5               g228(.a(new_n322), .b(new_n116), .o1(new_n324));
  xnbna2aa1n03x5               g229(.a(new_n110), .b(new_n324), .c(new_n118), .out0(\s[8] ));
  xorb03aa1n02x5               g230(.a(new_n140), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


