// Benchmark "adder" written by ABC on Wed Jul 17 22:09:20 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n326, new_n328, new_n330, new_n332, new_n333,
    new_n335, new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n03x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n03x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n09x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  nor002aa1n02x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nanp02aa1n04x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  oai012aa1n02x5               g006(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  norp02aa1n02x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nano23aa1n03x7               g010(.a(new_n102), .b(new_n105), .c(new_n103), .d(new_n104), .out0(new_n106));
  nanp02aa1n02x5               g011(.a(\b[0] ), .b(\a[1] ), .o1(new_n107));
  norp02aa1n02x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  norb03aa1n02x5               g013(.a(new_n101), .b(new_n108), .c(new_n107), .out0(new_n109));
  nanb02aa1n06x5               g014(.a(new_n109), .b(new_n106), .out0(new_n110));
  norp02aa1n02x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  aoi012aa1n02x5               g016(.a(new_n105), .b(new_n111), .c(new_n103), .o1(new_n112));
  xorc02aa1n02x5               g017(.a(\a[7] ), .b(\b[6] ), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  nanp02aa1n04x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nanb02aa1n02x5               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  tech160nm_fixorc02aa1n02p5x5 g022(.a(\a[8] ), .b(\b[7] ), .out0(new_n118));
  nona23aa1n06x5               g023(.a(new_n118), .b(new_n113), .c(new_n114), .d(new_n117), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\a[8] ), .o1(new_n120));
  orn002aa1n02x5               g025(.a(\a[7] ), .b(\b[6] ), .o(new_n121));
  norp02aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  oaih12aa1n02x5               g027(.a(new_n115), .b(new_n116), .c(new_n122), .o1(new_n123));
  nanp02aa1n02x5               g028(.a(new_n123), .b(new_n121), .o1(new_n124));
  aoi022aa1n02x5               g029(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n125));
  aboi22aa1n03x5               g030(.a(\b[7] ), .b(new_n120), .c(new_n124), .d(new_n125), .out0(new_n126));
  aoai13aa1n12x5               g031(.a(new_n126), .b(new_n119), .c(new_n110), .d(new_n112), .o1(new_n127));
  xorc02aa1n12x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n99), .b(new_n100), .c(new_n127), .d(new_n128), .o1(new_n129));
  nand22aa1n03x5               g034(.a(new_n127), .b(new_n128), .o1(new_n130));
  nona22aa1n02x4               g035(.a(new_n130), .b(new_n100), .c(new_n99), .out0(new_n131));
  nanp02aa1n02x5               g036(.a(new_n131), .b(new_n129), .o1(\s[10] ));
  inv000aa1d42x5               g037(.a(\a[11] ), .o1(new_n133));
  inv000aa1d42x5               g038(.a(\b[10] ), .o1(new_n134));
  nand42aa1n03x5               g039(.a(new_n134), .b(new_n133), .o1(new_n135));
  nanp02aa1n02x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  aoi022aa1n02x5               g041(.a(new_n131), .b(new_n98), .c(new_n135), .d(new_n136), .o1(new_n137));
  aoi022aa1n02x5               g042(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n138));
  aoi013aa1n02x4               g043(.a(new_n137), .b(new_n135), .c(new_n131), .d(new_n138), .o1(\s[11] ));
  aob012aa1n02x5               g044(.a(new_n135), .b(new_n131), .c(new_n138), .out0(new_n140));
  tech160nm_fixorc02aa1n03p5x5 g045(.a(\a[12] ), .b(\b[11] ), .out0(new_n141));
  aoi122aa1n06x5               g046(.a(new_n141), .b(new_n134), .c(new_n133), .d(new_n131), .e(new_n138), .o1(new_n142));
  tech160nm_fiaoi012aa1n02p5x5 g047(.a(new_n142), .b(new_n140), .c(new_n141), .o1(\s[12] ));
  nanp02aa1n02x5               g048(.a(new_n135), .b(new_n136), .o1(new_n144));
  nona23aa1n08x5               g049(.a(new_n141), .b(new_n128), .c(new_n99), .d(new_n144), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  oa0022aa1n02x5               g051(.a(\a[12] ), .b(\b[11] ), .c(\a[11] ), .d(\b[10] ), .o(new_n147));
  oai112aa1n02x5               g052(.a(new_n136), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n148));
  aoi022aa1n02x5               g053(.a(new_n148), .b(new_n147), .c(\a[12] ), .d(\b[11] ), .o1(new_n149));
  xorc02aa1n02x5               g054(.a(\a[13] ), .b(\b[12] ), .out0(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n149), .c(new_n127), .d(new_n146), .o1(new_n151));
  aoi112aa1n02x5               g056(.a(new_n150), .b(new_n149), .c(new_n127), .d(new_n146), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n151), .b(new_n152), .out0(\s[13] ));
  nor042aa1n06x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  xorc02aa1n02x5               g060(.a(\a[14] ), .b(\b[13] ), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n151), .c(new_n155), .out0(\s[14] ));
  inv000aa1d42x5               g062(.a(\a[13] ), .o1(new_n158));
  inv000aa1d42x5               g063(.a(\a[14] ), .o1(new_n159));
  xroi22aa1d04x5               g064(.a(new_n158), .b(\b[12] ), .c(new_n159), .d(\b[13] ), .out0(new_n160));
  aoai13aa1n06x5               g065(.a(new_n160), .b(new_n149), .c(new_n127), .d(new_n146), .o1(new_n161));
  oao003aa1n02x5               g066(.a(\a[14] ), .b(\b[13] ), .c(new_n155), .carry(new_n162));
  xorc02aa1n02x5               g067(.a(\a[15] ), .b(\b[14] ), .out0(new_n163));
  xnbna2aa1n03x5               g068(.a(new_n163), .b(new_n161), .c(new_n162), .out0(\s[15] ));
  aob012aa1n03x5               g069(.a(new_n163), .b(new_n161), .c(new_n162), .out0(new_n165));
  nor042aa1n03x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  inv000aa1d42x5               g071(.a(new_n166), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n163), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n167), .b(new_n168), .c(new_n161), .d(new_n162), .o1(new_n169));
  xorc02aa1n02x5               g074(.a(\a[16] ), .b(\b[15] ), .out0(new_n170));
  norp02aa1n02x5               g075(.a(new_n170), .b(new_n166), .o1(new_n171));
  aoi022aa1n03x5               g076(.a(new_n169), .b(new_n170), .c(new_n165), .d(new_n171), .o1(\s[16] ));
  nanp02aa1n02x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  xnrc02aa1n02x5               g078(.a(\b[15] ), .b(\a[16] ), .out0(new_n174));
  nano22aa1n12x5               g079(.a(new_n174), .b(new_n167), .c(new_n173), .out0(new_n175));
  nano22aa1d15x5               g080(.a(new_n145), .b(new_n160), .c(new_n175), .out0(new_n176));
  nanp02aa1n09x5               g081(.a(new_n127), .b(new_n176), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  aoi012aa1n02x5               g083(.a(new_n154), .b(\a[12] ), .c(\b[11] ), .o1(new_n179));
  obai22aa1n02x7               g084(.a(\b[12] ), .b(new_n158), .c(\b[13] ), .d(\a[14] ), .out0(new_n180));
  nanb03aa1n02x5               g085(.a(new_n180), .b(new_n178), .c(new_n179), .out0(new_n181));
  aoai13aa1n02x5               g086(.a(new_n162), .b(new_n181), .c(new_n148), .d(new_n147), .o1(new_n182));
  oao003aa1n02x5               g087(.a(\a[16] ), .b(\b[15] ), .c(new_n167), .carry(new_n183));
  aobi12aa1n02x5               g088(.a(new_n183), .b(new_n182), .c(new_n175), .out0(new_n184));
  xorc02aa1n12x5               g089(.a(\a[17] ), .b(\b[16] ), .out0(new_n185));
  xnbna2aa1n03x5               g090(.a(new_n185), .b(new_n177), .c(new_n184), .out0(\s[17] ));
  inv000aa1d42x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  nanp02aa1n02x5               g093(.a(new_n188), .b(new_n187), .o1(new_n189));
  inv000aa1d42x5               g094(.a(new_n175), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(\b[11] ), .b(\a[12] ), .o1(new_n191));
  nano32aa1n02x4               g096(.a(new_n180), .b(new_n155), .c(new_n178), .d(new_n191), .out0(new_n192));
  aob012aa1n02x5               g097(.a(new_n192), .b(new_n148), .c(new_n147), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n183), .b(new_n190), .c(new_n193), .d(new_n162), .o1(new_n194));
  aoai13aa1n02x5               g099(.a(new_n185), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n195));
  nor002aa1n02x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nand42aa1n02x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  norb02aa1n06x4               g102(.a(new_n197), .b(new_n196), .out0(new_n198));
  xnbna2aa1n03x5               g103(.a(new_n198), .b(new_n195), .c(new_n189), .out0(\s[18] ));
  and002aa1n02x5               g104(.a(new_n185), .b(new_n198), .o(new_n200));
  aoai13aa1n02x5               g105(.a(new_n200), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n201));
  aoi013aa1n06x5               g106(.a(new_n196), .b(new_n197), .c(new_n187), .d(new_n188), .o1(new_n202));
  nor042aa1n06x5               g107(.a(\b[18] ), .b(\a[19] ), .o1(new_n203));
  nand42aa1n02x5               g108(.a(\b[18] ), .b(\a[19] ), .o1(new_n204));
  norb02aa1n02x5               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n201), .c(new_n202), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nand02aa1d08x5               g112(.a(new_n177), .b(new_n184), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n189), .o1(new_n209));
  aoai13aa1n03x5               g114(.a(new_n205), .b(new_n209), .c(new_n208), .d(new_n200), .o1(new_n210));
  inv000aa1n03x5               g115(.a(new_n203), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n205), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n211), .b(new_n212), .c(new_n201), .d(new_n202), .o1(new_n213));
  nor002aa1n03x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand42aa1n02x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  inv000aa1d42x5               g121(.a(\a[19] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[18] ), .o1(new_n218));
  aboi22aa1n03x5               g123(.a(new_n214), .b(new_n215), .c(new_n217), .d(new_n218), .out0(new_n219));
  aoi022aa1n03x5               g124(.a(new_n213), .b(new_n216), .c(new_n210), .d(new_n219), .o1(\s[20] ));
  nano23aa1n06x5               g125(.a(new_n203), .b(new_n214), .c(new_n215), .d(new_n204), .out0(new_n221));
  nand23aa1n06x5               g126(.a(new_n221), .b(new_n185), .c(new_n198), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  aoai13aa1n02x5               g128(.a(new_n223), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n224));
  nona23aa1n09x5               g129(.a(new_n215), .b(new_n204), .c(new_n203), .d(new_n214), .out0(new_n225));
  oaoi03aa1n09x5               g130(.a(\a[20] ), .b(\b[19] ), .c(new_n211), .o1(new_n226));
  inv040aa1n03x5               g131(.a(new_n226), .o1(new_n227));
  oai012aa1d24x5               g132(.a(new_n227), .b(new_n225), .c(new_n202), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  xnbna2aa1n03x5               g136(.a(new_n231), .b(new_n224), .c(new_n229), .out0(\s[21] ));
  aoai13aa1n06x5               g137(.a(new_n231), .b(new_n228), .c(new_n208), .d(new_n223), .o1(new_n233));
  nor042aa1n03x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  inv000aa1n03x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n02x5               g140(.a(new_n235), .b(new_n230), .c(new_n224), .d(new_n229), .o1(new_n236));
  xnrc02aa1n12x5               g141(.a(\b[21] ), .b(\a[22] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n237), .b(new_n234), .out0(new_n239));
  aoi022aa1n02x5               g144(.a(new_n236), .b(new_n238), .c(new_n233), .d(new_n239), .o1(\s[22] ));
  nor042aa1n06x5               g145(.a(new_n237), .b(new_n230), .o1(new_n241));
  norb02aa1n03x5               g146(.a(new_n241), .b(new_n222), .out0(new_n242));
  aoai13aa1n02x5               g147(.a(new_n242), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n243));
  oao003aa1n12x5               g148(.a(\a[22] ), .b(\b[21] ), .c(new_n235), .carry(new_n244));
  inv000aa1d42x5               g149(.a(new_n244), .o1(new_n245));
  aoi012aa1d18x5               g150(.a(new_n245), .b(new_n228), .c(new_n241), .o1(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xorc02aa1n12x5               g152(.a(\a[23] ), .b(\b[22] ), .out0(new_n248));
  aoai13aa1n06x5               g153(.a(new_n248), .b(new_n247), .c(new_n208), .d(new_n242), .o1(new_n249));
  aoi112aa1n02x5               g154(.a(new_n248), .b(new_n245), .c(new_n228), .d(new_n241), .o1(new_n250));
  aobi12aa1n02x7               g155(.a(new_n249), .b(new_n250), .c(new_n243), .out0(\s[23] ));
  nor042aa1n03x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n248), .o1(new_n254));
  aoai13aa1n02x5               g159(.a(new_n253), .b(new_n254), .c(new_n243), .d(new_n246), .o1(new_n255));
  xorc02aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  norp02aa1n02x5               g161(.a(new_n256), .b(new_n252), .o1(new_n257));
  aoi022aa1n02x5               g162(.a(new_n255), .b(new_n256), .c(new_n249), .d(new_n257), .o1(\s[24] ));
  nano32aa1n03x7               g163(.a(new_n222), .b(new_n256), .c(new_n241), .d(new_n248), .out0(new_n259));
  aoai13aa1n02x5               g164(.a(new_n259), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n260));
  aoai13aa1n04x5               g165(.a(new_n241), .b(new_n226), .c(new_n221), .d(new_n209), .o1(new_n261));
  and002aa1n02x5               g166(.a(new_n256), .b(new_n248), .o(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  oao003aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .c(new_n253), .carry(new_n264));
  aoai13aa1n12x5               g169(.a(new_n264), .b(new_n263), .c(new_n261), .d(new_n244), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n265), .o1(new_n266));
  xorc02aa1n12x5               g171(.a(\a[25] ), .b(\b[24] ), .out0(new_n267));
  xnbna2aa1n03x5               g172(.a(new_n267), .b(new_n260), .c(new_n266), .out0(\s[25] ));
  aoai13aa1n03x5               g173(.a(new_n267), .b(new_n265), .c(new_n208), .d(new_n259), .o1(new_n269));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n267), .o1(new_n272));
  aoai13aa1n02x5               g177(.a(new_n271), .b(new_n272), .c(new_n260), .d(new_n266), .o1(new_n273));
  xorc02aa1n02x5               g178(.a(\a[26] ), .b(\b[25] ), .out0(new_n274));
  norp02aa1n02x5               g179(.a(new_n274), .b(new_n270), .o1(new_n275));
  aoi022aa1n03x5               g180(.a(new_n273), .b(new_n274), .c(new_n269), .d(new_n275), .o1(\s[26] ));
  and002aa1n02x5               g181(.a(new_n274), .b(new_n267), .o(new_n277));
  inv000aa1n02x5               g182(.a(new_n277), .o1(new_n278));
  nano23aa1d12x5               g183(.a(new_n278), .b(new_n222), .c(new_n262), .d(new_n241), .out0(new_n279));
  aoai13aa1n06x5               g184(.a(new_n279), .b(new_n194), .c(new_n127), .d(new_n176), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n262), .b(new_n245), .c(new_n228), .d(new_n241), .o1(new_n281));
  nanp02aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .o1(new_n282));
  oai022aa1n02x5               g187(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n283));
  nanp02aa1n02x5               g188(.a(new_n283), .b(new_n282), .o1(new_n284));
  aoai13aa1n06x5               g189(.a(new_n284), .b(new_n278), .c(new_n281), .d(new_n264), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n285), .c(new_n208), .d(new_n279), .o1(new_n287));
  aoi122aa1n02x5               g192(.a(new_n286), .b(new_n282), .c(new_n283), .d(new_n265), .e(new_n277), .o1(new_n288));
  aobi12aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n280), .out0(\s[27] ));
  aoi022aa1n09x5               g194(.a(new_n265), .b(new_n277), .c(new_n282), .d(new_n283), .o1(new_n290));
  norp02aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o1(new_n291));
  inv000aa1n03x5               g196(.a(new_n291), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n286), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n292), .b(new_n293), .c(new_n290), .d(new_n280), .o1(new_n294));
  tech160nm_fixorc02aa1n03p5x5 g199(.a(\a[28] ), .b(\b[27] ), .out0(new_n295));
  norp02aa1n02x5               g200(.a(new_n295), .b(new_n291), .o1(new_n296));
  aoi022aa1n03x5               g201(.a(new_n294), .b(new_n295), .c(new_n287), .d(new_n296), .o1(\s[28] ));
  and002aa1n02x5               g202(.a(new_n295), .b(new_n286), .o(new_n298));
  aoai13aa1n02x5               g203(.a(new_n298), .b(new_n285), .c(new_n208), .d(new_n279), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n298), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .carry(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n300), .c(new_n290), .d(new_n280), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[29] ), .b(\b[28] ), .out0(new_n303));
  norb02aa1n02x5               g208(.a(new_n301), .b(new_n303), .out0(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n299), .d(new_n304), .o1(\s[29] ));
  xorb03aa1n02x5               g210(.a(new_n107), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1d33x5               g211(.a(new_n293), .b(new_n295), .c(new_n303), .out0(new_n307));
  aoai13aa1n02x5               g212(.a(new_n307), .b(new_n285), .c(new_n208), .d(new_n279), .o1(new_n308));
  inv000aa1d42x5               g213(.a(new_n307), .o1(new_n309));
  oaoi03aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .o1(new_n310));
  inv000aa1n03x5               g215(.a(new_n310), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n309), .c(new_n290), .d(new_n280), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .out0(new_n313));
  and002aa1n02x5               g218(.a(\b[28] ), .b(\a[29] ), .o(new_n314));
  oabi12aa1n02x5               g219(.a(new_n313), .b(\a[29] ), .c(\b[28] ), .out0(new_n315));
  oab012aa1n02x4               g220(.a(new_n315), .b(new_n301), .c(new_n314), .out0(new_n316));
  aoi022aa1n03x5               g221(.a(new_n312), .b(new_n313), .c(new_n308), .d(new_n316), .o1(\s[30] ));
  nano32aa1n03x7               g222(.a(new_n293), .b(new_n313), .c(new_n295), .d(new_n303), .out0(new_n318));
  aoai13aa1n02x5               g223(.a(new_n318), .b(new_n285), .c(new_n208), .d(new_n279), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n318), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n320), .c(new_n290), .d(new_n280), .o1(new_n322));
  xorc02aa1n02x5               g227(.a(\a[31] ), .b(\b[30] ), .out0(new_n323));
  norb02aa1n02x5               g228(.a(new_n321), .b(new_n323), .out0(new_n324));
  aoi022aa1n03x5               g229(.a(new_n322), .b(new_n323), .c(new_n319), .d(new_n324), .o1(\s[31] ));
  oai012aa1n02x5               g230(.a(new_n101), .b(new_n108), .c(new_n107), .o1(new_n326));
  xnrb03aa1n02x5               g231(.a(new_n326), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g232(.a(\a[3] ), .b(\b[2] ), .c(new_n326), .o1(new_n328));
  xorb03aa1n02x5               g233(.a(new_n328), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorc02aa1n02x5               g234(.a(\a[5] ), .b(\b[4] ), .out0(new_n330));
  xnbna2aa1n03x5               g235(.a(new_n330), .b(new_n110), .c(new_n112), .out0(\s[5] ));
  orn002aa1n02x5               g236(.a(\a[5] ), .b(\b[4] ), .o(new_n332));
  aoai13aa1n02x5               g237(.a(new_n332), .b(new_n114), .c(new_n110), .d(new_n112), .o1(new_n333));
  xorb03aa1n02x5               g238(.a(new_n333), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  aoai13aa1n02x5               g239(.a(new_n113), .b(new_n116), .c(new_n333), .d(new_n115), .o1(new_n335));
  aoi112aa1n02x5               g240(.a(new_n116), .b(new_n113), .c(new_n333), .d(new_n115), .o1(new_n336));
  norb02aa1n02x5               g241(.a(new_n335), .b(new_n336), .out0(\s[7] ));
  xnbna2aa1n03x5               g242(.a(new_n118), .b(new_n335), .c(new_n121), .out0(\s[8] ));
  xorb03aa1n02x5               g243(.a(new_n127), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


