// Benchmark "adder" written by ABC on Thu Jul 18 12:21:13 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n356, new_n357, new_n359, new_n361,
    new_n362, new_n363, new_n364, new_n367, new_n369, new_n370;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n06x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n20x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nor002aa1d32x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  inv000aa1d42x5               g005(.a(new_n100), .o1(new_n101));
  inv040aa1d32x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand02aa1d08x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oaoi03aa1n12x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  nor002aa1d32x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nand22aa1n12x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nor002aa1d32x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  nand02aa1n10x5               g013(.a(\b[2] ), .b(\a[3] ), .o1(new_n109));
  nona23aa1d18x5               g014(.a(new_n109), .b(new_n107), .c(new_n106), .d(new_n108), .out0(new_n110));
  oaih12aa1n06x5               g015(.a(new_n107), .b(new_n108), .c(new_n106), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n111), .b(new_n110), .c(new_n105), .o1(new_n112));
  nor022aa1n12x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nand42aa1n04x5               g018(.a(\b[4] ), .b(\a[5] ), .o1(new_n114));
  nor002aa1d32x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nand42aa1n04x5               g020(.a(\b[5] ), .b(\a[6] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  xnrc02aa1n12x5               g022(.a(\b[6] ), .b(\a[7] ), .out0(new_n118));
  xnrc02aa1n12x5               g023(.a(\b[7] ), .b(\a[8] ), .out0(new_n119));
  nor043aa1n03x5               g024(.a(new_n117), .b(new_n118), .c(new_n119), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\a[8] ), .o1(new_n121));
  nor002aa1n04x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  nanp02aa1n02x5               g027(.a(\b[7] ), .b(\a[8] ), .o1(new_n123));
  oai022aa1n04x7               g028(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  aoi022aa1d24x5               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  aoai13aa1n04x5               g030(.a(new_n123), .b(new_n122), .c(new_n124), .d(new_n125), .o1(new_n126));
  oaib12aa1n06x5               g031(.a(new_n126), .b(\b[7] ), .c(new_n121), .out0(new_n127));
  nand42aa1n06x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n100), .out0(new_n129));
  aoai13aa1n02x5               g034(.a(new_n129), .b(new_n127), .c(new_n112), .d(new_n120), .o1(new_n130));
  xnbna2aa1n03x5               g035(.a(new_n99), .b(new_n130), .c(new_n101), .out0(\s[10] ));
  nand42aa1n02x5               g036(.a(new_n103), .b(new_n102), .o1(new_n132));
  nanp02aa1n04x5               g037(.a(\b[1] ), .b(\a[2] ), .o1(new_n133));
  aob012aa1n06x5               g038(.a(new_n132), .b(new_n104), .c(new_n133), .out0(new_n134));
  norb02aa1n06x5               g039(.a(new_n107), .b(new_n106), .out0(new_n135));
  norb02aa1n06x5               g040(.a(new_n109), .b(new_n108), .out0(new_n136));
  nand23aa1n04x5               g041(.a(new_n134), .b(new_n135), .c(new_n136), .o1(new_n137));
  nano23aa1n03x7               g042(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n138));
  nona22aa1n03x5               g043(.a(new_n138), .b(new_n118), .c(new_n119), .out0(new_n139));
  inv000aa1d42x5               g044(.a(\b[7] ), .o1(new_n140));
  inv020aa1n02x5               g045(.a(new_n122), .o1(new_n141));
  tech160nm_fioai012aa1n03p5x5 g046(.a(new_n125), .b(new_n115), .c(new_n113), .o1(new_n142));
  nanp02aa1n04x5               g047(.a(new_n142), .b(new_n141), .o1(new_n143));
  oaoi03aa1n09x5               g048(.a(new_n121), .b(new_n140), .c(new_n143), .o1(new_n144));
  aoai13aa1n06x5               g049(.a(new_n144), .b(new_n139), .c(new_n137), .d(new_n111), .o1(new_n145));
  oai022aa1n02x5               g050(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n146));
  nand42aa1n16x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  nor002aa1n20x5               g052(.a(\b[10] ), .b(\a[11] ), .o1(new_n148));
  nano22aa1n02x4               g053(.a(new_n148), .b(new_n98), .c(new_n147), .out0(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n146), .c(new_n145), .d(new_n129), .o1(new_n150));
  nanb02aa1n02x5               g055(.a(new_n148), .b(new_n147), .out0(new_n151));
  aoai13aa1n02x5               g056(.a(new_n98), .b(new_n146), .c(new_n145), .d(new_n129), .o1(new_n152));
  aobi12aa1n02x5               g057(.a(new_n150), .b(new_n152), .c(new_n151), .out0(\s[11] ));
  inv000aa1n04x5               g058(.a(new_n148), .o1(new_n154));
  nor042aa1d18x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand42aa1n16x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  norb02aa1n02x5               g061(.a(new_n156), .b(new_n155), .out0(new_n157));
  nona23aa1n02x4               g062(.a(new_n150), .b(new_n156), .c(new_n155), .d(new_n148), .out0(new_n158));
  aoai13aa1n02x5               g063(.a(new_n158), .b(new_n157), .c(new_n150), .d(new_n154), .o1(\s[12] ));
  nano23aa1n09x5               g064(.a(new_n155), .b(new_n148), .c(new_n156), .d(new_n147), .out0(new_n160));
  nano23aa1n09x5               g065(.a(new_n97), .b(new_n100), .c(new_n128), .d(new_n98), .out0(new_n161));
  nand22aa1n06x5               g066(.a(new_n161), .b(new_n160), .o1(new_n162));
  nanb02aa1n02x5               g067(.a(new_n162), .b(new_n145), .out0(new_n163));
  nanp02aa1n03x5               g068(.a(new_n112), .b(new_n120), .o1(new_n164));
  nanb03aa1n06x5               g069(.a(new_n155), .b(new_n156), .c(new_n147), .out0(new_n165));
  oai112aa1n04x5               g070(.a(new_n154), .b(new_n98), .c(new_n100), .d(new_n97), .o1(new_n166));
  tech160nm_fioai012aa1n03p5x5 g071(.a(new_n156), .b(new_n155), .c(new_n148), .o1(new_n167));
  oai012aa1n09x5               g072(.a(new_n167), .b(new_n166), .c(new_n165), .o1(new_n168));
  inv000aa1n06x5               g073(.a(new_n168), .o1(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n162), .c(new_n164), .d(new_n144), .o1(new_n170));
  nor002aa1n20x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nand42aa1d28x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n172), .b(new_n171), .out0(new_n173));
  nano32aa1n02x4               g078(.a(new_n165), .b(new_n146), .c(new_n154), .d(new_n98), .out0(new_n174));
  norb03aa1n02x5               g079(.a(new_n167), .b(new_n174), .c(new_n173), .out0(new_n175));
  aoi022aa1n02x5               g080(.a(new_n170), .b(new_n173), .c(new_n163), .d(new_n175), .o1(\s[13] ));
  inv000aa1d42x5               g081(.a(new_n171), .o1(new_n177));
  nanp02aa1n02x5               g082(.a(new_n170), .b(new_n173), .o1(new_n178));
  nor042aa1n04x5               g083(.a(\b[13] ), .b(\a[14] ), .o1(new_n179));
  nand42aa1d28x5               g084(.a(\b[13] ), .b(\a[14] ), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  oai022aa1d18x5               g086(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n182));
  nanb03aa1n02x5               g087(.a(new_n182), .b(new_n178), .c(new_n180), .out0(new_n183));
  aoai13aa1n03x5               g088(.a(new_n183), .b(new_n181), .c(new_n177), .d(new_n178), .o1(\s[14] ));
  nano23aa1d15x5               g089(.a(new_n171), .b(new_n179), .c(new_n180), .d(new_n172), .out0(new_n185));
  oaoi03aa1n02x5               g090(.a(\a[14] ), .b(\b[13] ), .c(new_n177), .o1(new_n186));
  xorc02aa1n12x5               g091(.a(\a[15] ), .b(\b[14] ), .out0(new_n187));
  aoai13aa1n06x5               g092(.a(new_n187), .b(new_n186), .c(new_n170), .d(new_n185), .o1(new_n188));
  aoi112aa1n02x5               g093(.a(new_n187), .b(new_n186), .c(new_n170), .d(new_n185), .o1(new_n189));
  norb02aa1n02x5               g094(.a(new_n188), .b(new_n189), .out0(\s[15] ));
  inv000aa1d42x5               g095(.a(\a[15] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\b[14] ), .o1(new_n192));
  nanp02aa1n02x5               g097(.a(new_n192), .b(new_n191), .o1(new_n193));
  nor042aa1d18x5               g098(.a(\b[15] ), .b(\a[16] ), .o1(new_n194));
  and002aa1n12x5               g099(.a(\b[15] ), .b(\a[16] ), .o(new_n195));
  nor042aa1n04x5               g100(.a(new_n195), .b(new_n194), .o1(new_n196));
  oai022aa1n02x5               g101(.a(\a[15] ), .b(\b[14] ), .c(\b[15] ), .d(\a[16] ), .o1(new_n197));
  nona22aa1n03x5               g102(.a(new_n188), .b(new_n195), .c(new_n197), .out0(new_n198));
  aoai13aa1n02x5               g103(.a(new_n198), .b(new_n196), .c(new_n193), .d(new_n188), .o1(\s[16] ));
  nand23aa1d12x5               g104(.a(new_n185), .b(new_n187), .c(new_n196), .o1(new_n200));
  nor042aa1n06x5               g105(.a(new_n200), .b(new_n162), .o1(new_n201));
  aoai13aa1n12x5               g106(.a(new_n201), .b(new_n127), .c(new_n112), .d(new_n120), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n194), .o1(new_n203));
  oai112aa1n04x5               g108(.a(new_n182), .b(new_n180), .c(new_n192), .d(new_n191), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n203), .b(new_n195), .c(new_n204), .d(new_n193), .o1(new_n205));
  aoib12aa1n09x5               g110(.a(new_n205), .b(new_n168), .c(new_n200), .out0(new_n206));
  nanp02aa1n12x5               g111(.a(new_n202), .b(new_n206), .o1(new_n207));
  nor042aa1d18x5               g112(.a(\b[16] ), .b(\a[17] ), .o1(new_n208));
  nand42aa1n02x5               g113(.a(\b[16] ), .b(\a[17] ), .o1(new_n209));
  norb02aa1n02x5               g114(.a(new_n209), .b(new_n208), .out0(new_n210));
  aoi022aa1n02x5               g115(.a(new_n204), .b(new_n193), .c(\a[16] ), .d(\b[15] ), .o1(new_n211));
  nona22aa1n02x4               g116(.a(new_n203), .b(new_n211), .c(new_n210), .out0(new_n212));
  aoib12aa1n02x5               g117(.a(new_n212), .b(new_n168), .c(new_n200), .out0(new_n213));
  aoi022aa1n02x5               g118(.a(new_n207), .b(new_n210), .c(new_n213), .d(new_n202), .o1(\s[17] ));
  inv000aa1d42x5               g119(.a(new_n208), .o1(new_n215));
  oabi12aa1n06x5               g120(.a(new_n205), .b(new_n169), .c(new_n200), .out0(new_n216));
  aoai13aa1n02x5               g121(.a(new_n210), .b(new_n216), .c(new_n145), .d(new_n201), .o1(new_n217));
  nor042aa1n06x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  nand02aa1n06x5               g123(.a(\b[17] ), .b(\a[18] ), .o1(new_n219));
  norb02aa1n02x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  nona23aa1n02x4               g125(.a(new_n217), .b(new_n219), .c(new_n218), .d(new_n208), .out0(new_n221));
  aoai13aa1n02x5               g126(.a(new_n221), .b(new_n220), .c(new_n215), .d(new_n217), .o1(\s[18] ));
  nano23aa1n06x5               g127(.a(new_n208), .b(new_n218), .c(new_n219), .d(new_n209), .out0(new_n223));
  oaoi03aa1n02x5               g128(.a(\a[18] ), .b(\b[17] ), .c(new_n215), .o1(new_n224));
  nor002aa1n16x5               g129(.a(\b[18] ), .b(\a[19] ), .o1(new_n225));
  nand02aa1n03x5               g130(.a(\b[18] ), .b(\a[19] ), .o1(new_n226));
  norb02aa1n06x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n207), .d(new_n223), .o1(new_n228));
  aoi112aa1n02x5               g133(.a(new_n227), .b(new_n224), .c(new_n207), .d(new_n223), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n228), .b(new_n229), .out0(\s[19] ));
  xnrc02aa1n02x5               g135(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1n02x5               g136(.a(new_n225), .o1(new_n232));
  nor042aa1n04x5               g137(.a(\b[19] ), .b(\a[20] ), .o1(new_n233));
  nand22aa1n04x5               g138(.a(\b[19] ), .b(\a[20] ), .o1(new_n234));
  norb02aa1n06x4               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  norb03aa1n02x5               g140(.a(new_n234), .b(new_n225), .c(new_n233), .out0(new_n236));
  tech160nm_finand02aa1n03p5x5 g141(.a(new_n228), .b(new_n236), .o1(new_n237));
  aoai13aa1n03x5               g142(.a(new_n237), .b(new_n235), .c(new_n232), .d(new_n228), .o1(\s[20] ));
  nand23aa1n03x5               g143(.a(new_n223), .b(new_n227), .c(new_n235), .o1(new_n239));
  inv040aa1n03x5               g144(.a(new_n239), .o1(new_n240));
  nanb03aa1n06x5               g145(.a(new_n233), .b(new_n234), .c(new_n226), .out0(new_n241));
  oai112aa1n03x5               g146(.a(new_n232), .b(new_n219), .c(new_n218), .d(new_n208), .o1(new_n242));
  aoi012aa1n06x5               g147(.a(new_n233), .b(new_n225), .c(new_n234), .o1(new_n243));
  tech160nm_fioai012aa1n05x5   g148(.a(new_n243), .b(new_n242), .c(new_n241), .o1(new_n244));
  nor002aa1d32x5               g149(.a(\b[20] ), .b(\a[21] ), .o1(new_n245));
  nanp02aa1n04x5               g150(.a(\b[20] ), .b(\a[21] ), .o1(new_n246));
  norb02aa1n02x5               g151(.a(new_n246), .b(new_n245), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n244), .c(new_n207), .d(new_n240), .o1(new_n248));
  nano22aa1n03x7               g153(.a(new_n233), .b(new_n226), .c(new_n234), .out0(new_n249));
  tech160nm_fioai012aa1n03p5x5 g154(.a(new_n219), .b(\b[18] ), .c(\a[19] ), .o1(new_n250));
  oab012aa1n06x5               g155(.a(new_n250), .b(new_n208), .c(new_n218), .out0(new_n251));
  inv020aa1n02x5               g156(.a(new_n243), .o1(new_n252));
  aoi112aa1n02x5               g157(.a(new_n252), .b(new_n247), .c(new_n251), .d(new_n249), .o1(new_n253));
  aobi12aa1n02x5               g158(.a(new_n253), .b(new_n207), .c(new_n240), .out0(new_n254));
  norb02aa1n03x4               g159(.a(new_n248), .b(new_n254), .out0(\s[21] ));
  inv000aa1d42x5               g160(.a(new_n245), .o1(new_n256));
  nor042aa1n03x5               g161(.a(\b[21] ), .b(\a[22] ), .o1(new_n257));
  nand42aa1n04x5               g162(.a(\b[21] ), .b(\a[22] ), .o1(new_n258));
  norb02aa1n02x5               g163(.a(new_n258), .b(new_n257), .out0(new_n259));
  norb03aa1n02x5               g164(.a(new_n258), .b(new_n245), .c(new_n257), .out0(new_n260));
  nand42aa1n03x5               g165(.a(new_n248), .b(new_n260), .o1(new_n261));
  aoai13aa1n03x5               g166(.a(new_n261), .b(new_n259), .c(new_n256), .d(new_n248), .o1(\s[22] ));
  nano23aa1d15x5               g167(.a(new_n245), .b(new_n257), .c(new_n258), .d(new_n246), .out0(new_n263));
  inv000aa1n02x5               g168(.a(new_n263), .o1(new_n264));
  nano32aa1n02x4               g169(.a(new_n264), .b(new_n223), .c(new_n227), .d(new_n235), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n263), .b(new_n252), .c(new_n251), .d(new_n249), .o1(new_n266));
  oaoi03aa1n12x5               g171(.a(\a[22] ), .b(\b[21] ), .c(new_n256), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n267), .o1(new_n268));
  nanp02aa1n02x5               g173(.a(new_n266), .b(new_n268), .o1(new_n269));
  xorc02aa1n12x5               g174(.a(\a[23] ), .b(\b[22] ), .out0(new_n270));
  aoai13aa1n06x5               g175(.a(new_n270), .b(new_n269), .c(new_n207), .d(new_n265), .o1(new_n271));
  nona22aa1n02x4               g176(.a(new_n266), .b(new_n267), .c(new_n270), .out0(new_n272));
  aoi012aa1n02x5               g177(.a(new_n272), .b(new_n207), .c(new_n265), .o1(new_n273));
  norb02aa1n03x4               g178(.a(new_n271), .b(new_n273), .out0(\s[23] ));
  norp02aa1n02x5               g179(.a(\b[22] ), .b(\a[23] ), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[24] ), .b(\b[23] ), .out0(new_n277));
  oai022aa1n02x5               g182(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n278));
  aoi012aa1n02x5               g183(.a(new_n278), .b(\a[24] ), .c(\b[23] ), .o1(new_n279));
  nand42aa1n03x5               g184(.a(new_n271), .b(new_n279), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n277), .c(new_n276), .d(new_n271), .o1(\s[24] ));
  nano32aa1n03x7               g186(.a(new_n239), .b(new_n277), .c(new_n263), .d(new_n270), .out0(new_n282));
  nand22aa1n03x5               g187(.a(new_n277), .b(new_n270), .o1(new_n283));
  aob012aa1n02x5               g188(.a(new_n278), .b(\b[23] ), .c(\a[24] ), .out0(new_n284));
  aoai13aa1n04x5               g189(.a(new_n284), .b(new_n283), .c(new_n266), .d(new_n268), .o1(new_n285));
  xorc02aa1n12x5               g190(.a(\a[25] ), .b(\b[24] ), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n285), .c(new_n207), .d(new_n282), .o1(new_n287));
  inv000aa1n02x5               g192(.a(new_n283), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n267), .c(new_n244), .d(new_n263), .o1(new_n289));
  nanb03aa1n02x5               g194(.a(new_n286), .b(new_n289), .c(new_n284), .out0(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(new_n207), .c(new_n282), .o1(new_n291));
  norb02aa1n02x5               g196(.a(new_n287), .b(new_n291), .out0(\s[25] ));
  norp02aa1n02x5               g197(.a(\b[24] ), .b(\a[25] ), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  tech160nm_fixorc02aa1n05x5   g199(.a(\a[26] ), .b(\b[25] ), .out0(new_n295));
  nanp02aa1n02x5               g200(.a(\b[25] ), .b(\a[26] ), .o1(new_n296));
  oai022aa1n02x5               g201(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n297));
  norb02aa1n02x5               g202(.a(new_n296), .b(new_n297), .out0(new_n298));
  tech160nm_finand02aa1n03p5x5 g203(.a(new_n287), .b(new_n298), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n295), .c(new_n294), .d(new_n287), .o1(\s[26] ));
  nand02aa1n04x5               g205(.a(new_n295), .b(new_n286), .o1(new_n301));
  nano23aa1n03x7               g206(.a(new_n239), .b(new_n301), .c(new_n288), .d(new_n263), .out0(new_n302));
  aoai13aa1n06x5               g207(.a(new_n302), .b(new_n216), .c(new_n145), .d(new_n201), .o1(new_n303));
  nona32aa1n09x5               g208(.a(new_n240), .b(new_n301), .c(new_n283), .d(new_n264), .out0(new_n304));
  aoi012aa1n06x5               g209(.a(new_n304), .b(new_n202), .c(new_n206), .o1(new_n305));
  nanp02aa1n02x5               g210(.a(new_n297), .b(new_n296), .o1(new_n306));
  aoai13aa1n06x5               g211(.a(new_n306), .b(new_n301), .c(new_n289), .d(new_n284), .o1(new_n307));
  xorc02aa1n12x5               g212(.a(\a[27] ), .b(\b[26] ), .out0(new_n308));
  oaih12aa1n02x5               g213(.a(new_n308), .b(new_n307), .c(new_n305), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n301), .o1(new_n310));
  aoi122aa1n02x5               g215(.a(new_n308), .b(new_n296), .c(new_n297), .d(new_n285), .e(new_n310), .o1(new_n311));
  aobi12aa1n02x7               g216(.a(new_n309), .b(new_n311), .c(new_n303), .out0(\s[27] ));
  nor002aa1n03x5               g217(.a(\b[26] ), .b(\a[27] ), .o1(new_n313));
  inv020aa1n02x5               g218(.a(new_n313), .o1(new_n314));
  nor002aa1n03x5               g219(.a(\b[27] ), .b(\a[28] ), .o1(new_n315));
  and002aa1n12x5               g220(.a(\b[27] ), .b(\a[28] ), .o(new_n316));
  nor002aa1n02x5               g221(.a(new_n316), .b(new_n315), .o1(new_n317));
  aoi022aa1n06x5               g222(.a(new_n285), .b(new_n310), .c(new_n296), .d(new_n297), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n308), .o1(new_n319));
  norp03aa1n02x5               g224(.a(new_n316), .b(new_n315), .c(new_n313), .o1(new_n320));
  aoai13aa1n06x5               g225(.a(new_n320), .b(new_n319), .c(new_n318), .d(new_n303), .o1(new_n321));
  aoai13aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n309), .d(new_n314), .o1(\s[28] ));
  and002aa1n02x5               g227(.a(new_n308), .b(new_n317), .o(new_n323));
  oaih12aa1n02x5               g228(.a(new_n323), .b(new_n307), .c(new_n305), .o1(new_n324));
  inv000aa1d42x5               g229(.a(new_n323), .o1(new_n325));
  oab012aa1n06x5               g230(.a(new_n315), .b(new_n314), .c(new_n316), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n326), .b(new_n325), .c(new_n318), .d(new_n303), .o1(new_n327));
  xorc02aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .out0(new_n328));
  norb02aa1n02x5               g233(.a(new_n326), .b(new_n328), .out0(new_n329));
  aoi022aa1n03x5               g234(.a(new_n327), .b(new_n328), .c(new_n324), .d(new_n329), .o1(\s[29] ));
  xorb03aa1n02x5               g235(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g236(.a(new_n319), .b(new_n328), .c(new_n317), .out0(new_n332));
  oaih12aa1n02x5               g237(.a(new_n332), .b(new_n307), .c(new_n305), .o1(new_n333));
  inv000aa1n02x5               g238(.a(new_n332), .o1(new_n334));
  tech160nm_fioaoi03aa1n03p5x5 g239(.a(\a[29] ), .b(\b[28] ), .c(new_n326), .o1(new_n335));
  inv000aa1d42x5               g240(.a(new_n335), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n334), .c(new_n318), .d(new_n303), .o1(new_n337));
  xorc02aa1n02x5               g242(.a(\a[30] ), .b(\b[29] ), .out0(new_n338));
  and002aa1n02x5               g243(.a(\b[28] ), .b(\a[29] ), .o(new_n339));
  oabi12aa1n02x5               g244(.a(new_n338), .b(\a[29] ), .c(\b[28] ), .out0(new_n340));
  oab012aa1n02x4               g245(.a(new_n340), .b(new_n326), .c(new_n339), .out0(new_n341));
  aoi022aa1n03x5               g246(.a(new_n337), .b(new_n338), .c(new_n333), .d(new_n341), .o1(\s[30] ));
  nano32aa1n02x4               g247(.a(new_n319), .b(new_n338), .c(new_n317), .d(new_n328), .out0(new_n343));
  oai012aa1n02x5               g248(.a(new_n343), .b(new_n307), .c(new_n305), .o1(new_n344));
  xorc02aa1n02x5               g249(.a(\a[31] ), .b(\b[30] ), .out0(new_n345));
  inv000aa1d42x5               g250(.a(\a[30] ), .o1(new_n346));
  inv000aa1d42x5               g251(.a(\b[29] ), .o1(new_n347));
  oabi12aa1n02x5               g252(.a(new_n345), .b(\a[30] ), .c(\b[29] ), .out0(new_n348));
  oaoi13aa1n02x5               g253(.a(new_n348), .b(new_n335), .c(new_n346), .d(new_n347), .o1(new_n349));
  inv000aa1n02x5               g254(.a(new_n343), .o1(new_n350));
  tech160nm_fioaoi03aa1n03p5x5 g255(.a(new_n346), .b(new_n347), .c(new_n335), .o1(new_n351));
  aoai13aa1n03x5               g256(.a(new_n351), .b(new_n350), .c(new_n318), .d(new_n303), .o1(new_n352));
  aoi022aa1n03x5               g257(.a(new_n352), .b(new_n345), .c(new_n344), .d(new_n349), .o1(\s[31] ));
  nanp03aa1n02x5               g258(.a(new_n132), .b(new_n104), .c(new_n133), .o1(new_n354));
  xnbna2aa1n03x5               g259(.a(new_n136), .b(new_n354), .c(new_n132), .out0(\s[3] ));
  inv000aa1d42x5               g260(.a(new_n108), .o1(new_n356));
  nanp02aa1n02x5               g261(.a(new_n134), .b(new_n136), .o1(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n135), .b(new_n357), .c(new_n356), .out0(\s[4] ));
  norb02aa1n02x5               g263(.a(new_n114), .b(new_n113), .out0(new_n359));
  xnbna2aa1n03x5               g264(.a(new_n359), .b(new_n137), .c(new_n111), .out0(\s[5] ));
  nanb02aa1n02x5               g265(.a(new_n115), .b(new_n116), .out0(new_n361));
  aoai13aa1n02x5               g266(.a(new_n361), .b(new_n113), .c(new_n112), .d(new_n114), .o1(new_n362));
  norb03aa1n02x5               g267(.a(new_n116), .b(new_n113), .c(new_n115), .out0(new_n363));
  aob012aa1n02x5               g268(.a(new_n363), .b(new_n112), .c(new_n359), .out0(new_n364));
  nanp02aa1n02x5               g269(.a(new_n362), .b(new_n364), .o1(\s[6] ));
  xnbna2aa1n03x5               g270(.a(new_n118), .b(new_n364), .c(new_n116), .out0(\s[7] ));
  nanb03aa1n02x5               g271(.a(new_n118), .b(new_n364), .c(new_n116), .out0(new_n367));
  xobna2aa1n03x5               g272(.a(new_n119), .b(new_n367), .c(new_n141), .out0(\s[8] ));
  obai22aa1n02x7               g273(.a(new_n128), .b(new_n100), .c(\a[8] ), .d(\b[7] ), .out0(new_n369));
  aoi012aa1n02x5               g274(.a(new_n369), .b(new_n143), .c(new_n123), .o1(new_n370));
  aoi022aa1n02x5               g275(.a(new_n145), .b(new_n129), .c(new_n164), .d(new_n370), .o1(\s[9] ));
endmodule


