// Benchmark "adder" written by ABC on Wed Jul 17 17:47:59 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n175, new_n176, new_n177,
    new_n178, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n345,
    new_n346, new_n347, new_n350, new_n352, new_n353, new_n354, new_n355,
    new_n357, new_n358;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1n06x5               g002(.a(new_n97), .o1(new_n98));
  orn002aa1n02x7               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  tech160nm_finand02aa1n05x5   g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aob012aa1n12x5               g005(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(new_n101));
  nor042aa1n09x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nand22aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanb02aa1n03x5               g008(.a(new_n102), .b(new_n103), .out0(new_n104));
  nor042aa1n04x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor042aa1n12x5               g010(.a(new_n105), .b(new_n102), .o1(new_n106));
  aoai13aa1n04x5               g011(.a(new_n106), .b(new_n104), .c(new_n101), .d(new_n99), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[4] ), .b(\a[5] ), .o1(new_n108));
  norp02aa1n02x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  aoi012aa1n02x5               g014(.a(new_n109), .b(\a[6] ), .c(\b[5] ), .o1(new_n110));
  inv000aa1d42x5               g015(.a(\a[8] ), .o1(new_n111));
  inv000aa1d42x5               g016(.a(\b[7] ), .o1(new_n112));
  aoi022aa1n02x7               g017(.a(new_n112), .b(new_n111), .c(\a[4] ), .d(\b[3] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nor042aa1n04x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n04x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nor002aa1n16x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nona23aa1n03x5               g022(.a(new_n116), .b(new_n114), .c(new_n117), .d(new_n115), .out0(new_n118));
  nano32aa1n03x7               g023(.a(new_n118), .b(new_n113), .c(new_n110), .d(new_n108), .out0(new_n119));
  nanp02aa1n04x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nano22aa1n03x7               g025(.a(new_n115), .b(new_n120), .c(new_n116), .out0(new_n121));
  oai022aa1n04x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  xorc02aa1n12x5               g027(.a(\a[8] ), .b(\b[7] ), .out0(new_n123));
  nanp03aa1n02x5               g028(.a(new_n121), .b(new_n123), .c(new_n122), .o1(new_n124));
  oao003aa1n02x5               g029(.a(new_n111), .b(new_n112), .c(new_n115), .carry(new_n125));
  nanb02aa1n06x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  nand42aa1n03x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n97), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n126), .c(new_n107), .d(new_n119), .o1(new_n129));
  nor002aa1n08x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n10x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  xnbna2aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n98), .out0(\s[10] ));
  nanp02aa1n02x5               g038(.a(new_n101), .b(new_n99), .o1(new_n134));
  norb02aa1n06x4               g039(.a(new_n103), .b(new_n102), .out0(new_n135));
  inv000aa1d42x5               g040(.a(new_n106), .o1(new_n136));
  aoi012aa1n02x5               g041(.a(new_n136), .b(new_n134), .c(new_n135), .o1(new_n137));
  nano22aa1n02x4               g042(.a(new_n109), .b(new_n108), .c(new_n120), .out0(new_n138));
  nano23aa1n02x4               g043(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n139));
  nano32aa1n02x5               g044(.a(new_n137), .b(new_n139), .c(new_n138), .d(new_n113), .out0(new_n140));
  nona23aa1n09x5               g045(.a(new_n131), .b(new_n127), .c(new_n97), .d(new_n130), .out0(new_n141));
  oabi12aa1n02x5               g046(.a(new_n141), .b(new_n140), .c(new_n126), .out0(new_n142));
  oaoi03aa1n02x5               g047(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n143));
  inv020aa1n02x5               g048(.a(new_n143), .o1(new_n144));
  xnrc02aa1n12x5               g049(.a(\b[10] ), .b(\a[11] ), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  xnbna2aa1n03x5               g051(.a(new_n146), .b(new_n142), .c(new_n144), .out0(\s[11] ));
  inv040aa1d32x5               g052(.a(\a[11] ), .o1(new_n148));
  inv020aa1n08x5               g053(.a(\b[10] ), .o1(new_n149));
  nand42aa1n02x5               g054(.a(new_n149), .b(new_n148), .o1(new_n150));
  aob012aa1n02x5               g055(.a(new_n146), .b(new_n142), .c(new_n144), .out0(new_n151));
  inv040aa1d32x5               g056(.a(\a[12] ), .o1(new_n152));
  inv040aa1d28x5               g057(.a(\b[11] ), .o1(new_n153));
  nand22aa1n09x5               g058(.a(new_n153), .b(new_n152), .o1(new_n154));
  nand02aa1n08x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nand02aa1d04x5               g060(.a(new_n154), .b(new_n155), .o1(new_n156));
  inv000aa1d42x5               g061(.a(new_n156), .o1(new_n157));
  xnbna2aa1n03x5               g062(.a(new_n157), .b(new_n151), .c(new_n150), .out0(\s[12] ));
  nand42aa1n06x5               g063(.a(new_n119), .b(new_n107), .o1(new_n159));
  aoi013aa1n09x5               g064(.a(new_n125), .b(new_n121), .c(new_n123), .d(new_n122), .o1(new_n160));
  nand22aa1n03x5               g065(.a(new_n159), .b(new_n160), .o1(new_n161));
  nor043aa1n02x5               g066(.a(new_n141), .b(new_n145), .c(new_n156), .o1(new_n162));
  oai112aa1n02x7               g067(.a(new_n154), .b(new_n155), .c(new_n149), .d(new_n148), .o1(new_n163));
  oai112aa1n03x5               g068(.a(new_n131), .b(new_n150), .c(new_n130), .d(new_n97), .o1(new_n164));
  aoi112aa1n03x4               g069(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n165));
  norb02aa1n03x5               g070(.a(new_n154), .b(new_n165), .out0(new_n166));
  tech160nm_fioai012aa1n05x5   g071(.a(new_n166), .b(new_n164), .c(new_n163), .o1(new_n167));
  nor002aa1d32x5               g072(.a(\b[12] ), .b(\a[13] ), .o1(new_n168));
  nand22aa1n06x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nanb02aa1n02x5               g074(.a(new_n168), .b(new_n169), .out0(new_n170));
  inv000aa1d42x5               g075(.a(new_n170), .o1(new_n171));
  aoai13aa1n02x5               g076(.a(new_n171), .b(new_n167), .c(new_n161), .d(new_n162), .o1(new_n172));
  aoi112aa1n02x5               g077(.a(new_n171), .b(new_n167), .c(new_n161), .d(new_n162), .o1(new_n173));
  norb02aa1n02x5               g078(.a(new_n172), .b(new_n173), .out0(\s[13] ));
  inv000aa1d42x5               g079(.a(new_n168), .o1(new_n175));
  nor002aa1d32x5               g080(.a(\b[13] ), .b(\a[14] ), .o1(new_n176));
  nanp02aa1n12x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  xobna2aa1n03x5               g083(.a(new_n178), .b(new_n172), .c(new_n175), .out0(\s[14] ));
  nona23aa1d16x5               g084(.a(new_n177), .b(new_n169), .c(new_n168), .d(new_n176), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n180), .o1(new_n181));
  aoai13aa1n03x5               g086(.a(new_n181), .b(new_n167), .c(new_n161), .d(new_n162), .o1(new_n182));
  oaoi03aa1n02x5               g087(.a(\a[14] ), .b(\b[13] ), .c(new_n175), .o1(new_n183));
  inv000aa1d42x5               g088(.a(new_n183), .o1(new_n184));
  nor042aa1d18x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nanp02aa1n09x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  norb02aa1n06x5               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  xnbna2aa1n03x5               g092(.a(new_n187), .b(new_n182), .c(new_n184), .out0(\s[15] ));
  aob012aa1n03x5               g093(.a(new_n187), .b(new_n182), .c(new_n184), .out0(new_n189));
  nor042aa1n04x5               g094(.a(\b[15] ), .b(\a[16] ), .o1(new_n190));
  nand02aa1d08x5               g095(.a(\b[15] ), .b(\a[16] ), .o1(new_n191));
  norb02aa1n02x5               g096(.a(new_n191), .b(new_n190), .out0(new_n192));
  norp02aa1n02x5               g097(.a(new_n192), .b(new_n185), .o1(new_n193));
  inv000aa1n02x5               g098(.a(new_n185), .o1(new_n194));
  inv000aa1d42x5               g099(.a(new_n187), .o1(new_n195));
  aoai13aa1n02x7               g100(.a(new_n194), .b(new_n195), .c(new_n182), .d(new_n184), .o1(new_n196));
  aoi022aa1n03x5               g101(.a(new_n196), .b(new_n192), .c(new_n189), .d(new_n193), .o1(\s[16] ));
  nanb03aa1n02x5               g102(.a(new_n141), .b(new_n157), .c(new_n146), .out0(new_n198));
  nona23aa1d18x5               g103(.a(new_n191), .b(new_n186), .c(new_n185), .d(new_n190), .out0(new_n199));
  nor042aa1n09x5               g104(.a(new_n199), .b(new_n180), .o1(new_n200));
  norb02aa1n03x5               g105(.a(new_n200), .b(new_n198), .out0(new_n201));
  tech160nm_fioai012aa1n03p5x5 g106(.a(new_n201), .b(new_n140), .c(new_n126), .o1(new_n202));
  xorc02aa1n02x5               g107(.a(\a[17] ), .b(\b[16] ), .out0(new_n203));
  nanb03aa1n02x5               g108(.a(new_n190), .b(new_n191), .c(new_n186), .out0(new_n204));
  oai112aa1n02x7               g109(.a(new_n194), .b(new_n177), .c(new_n176), .d(new_n168), .o1(new_n205));
  aoi012aa1n02x7               g110(.a(new_n190), .b(new_n185), .c(new_n191), .o1(new_n206));
  oai012aa1n06x5               g111(.a(new_n206), .b(new_n205), .c(new_n204), .o1(new_n207));
  aoi112aa1n02x5               g112(.a(new_n207), .b(new_n203), .c(new_n167), .d(new_n200), .o1(new_n208));
  nona32aa1n03x5               g113(.a(new_n200), .b(new_n141), .c(new_n156), .d(new_n145), .out0(new_n209));
  aoi012aa1n12x5               g114(.a(new_n207), .b(new_n167), .c(new_n200), .o1(new_n210));
  aoai13aa1n12x5               g115(.a(new_n210), .b(new_n209), .c(new_n159), .d(new_n160), .o1(new_n211));
  aoi022aa1n02x5               g116(.a(new_n211), .b(new_n203), .c(new_n202), .d(new_n208), .o1(\s[17] ));
  inv040aa1d32x5               g117(.a(\a[17] ), .o1(new_n213));
  inv040aa1d32x5               g118(.a(\b[16] ), .o1(new_n214));
  nand42aa1n08x5               g119(.a(new_n214), .b(new_n213), .o1(new_n215));
  oaib12aa1n06x5               g120(.a(new_n211), .b(new_n214), .c(\a[17] ), .out0(new_n216));
  nor002aa1d32x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  nand42aa1d28x5               g122(.a(\b[17] ), .b(\a[18] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  xnbna2aa1n03x5               g124(.a(new_n219), .b(new_n216), .c(new_n215), .out0(\s[18] ));
  nand42aa1n06x5               g125(.a(\b[16] ), .b(\a[17] ), .o1(new_n221));
  nano32aa1n03x7               g126(.a(new_n217), .b(new_n215), .c(new_n218), .d(new_n221), .out0(new_n222));
  aoai13aa1n12x5               g127(.a(new_n218), .b(new_n217), .c(new_n213), .d(new_n214), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  xorc02aa1n12x5               g129(.a(\a[19] ), .b(\b[18] ), .out0(new_n225));
  aoai13aa1n06x5               g130(.a(new_n225), .b(new_n224), .c(new_n211), .d(new_n222), .o1(new_n226));
  aoi112aa1n02x5               g131(.a(new_n225), .b(new_n224), .c(new_n211), .d(new_n222), .o1(new_n227));
  norb02aa1n03x4               g132(.a(new_n226), .b(new_n227), .out0(\s[19] ));
  xnrc02aa1n02x5               g133(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  xorc02aa1n12x5               g134(.a(\a[20] ), .b(\b[19] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(\a[19] ), .o1(new_n231));
  inv000aa1d42x5               g136(.a(\b[18] ), .o1(new_n232));
  inv000aa1d42x5               g137(.a(\a[20] ), .o1(new_n233));
  inv000aa1d42x5               g138(.a(\b[19] ), .o1(new_n234));
  nanp02aa1n02x5               g139(.a(new_n234), .b(new_n233), .o1(new_n235));
  nanp02aa1n02x5               g140(.a(\b[19] ), .b(\a[20] ), .o1(new_n236));
  aoi022aa1n02x5               g141(.a(new_n235), .b(new_n236), .c(new_n232), .d(new_n231), .o1(new_n237));
  norp02aa1n04x5               g142(.a(\b[18] ), .b(\a[19] ), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n238), .o1(new_n239));
  nand42aa1n02x5               g144(.a(new_n226), .b(new_n239), .o1(new_n240));
  aoi022aa1n02x7               g145(.a(new_n240), .b(new_n230), .c(new_n226), .d(new_n237), .o1(\s[20] ));
  nand23aa1n04x5               g146(.a(new_n222), .b(new_n225), .c(new_n230), .o1(new_n242));
  inv000aa1d42x5               g147(.a(new_n242), .o1(new_n243));
  oai112aa1n02x5               g148(.a(new_n235), .b(new_n236), .c(new_n232), .d(new_n231), .o1(new_n244));
  oaoi03aa1n03x5               g149(.a(new_n233), .b(new_n234), .c(new_n238), .o1(new_n245));
  oai013aa1n03x5               g150(.a(new_n245), .b(new_n244), .c(new_n223), .d(new_n238), .o1(new_n246));
  xorc02aa1n12x5               g151(.a(\a[21] ), .b(\b[20] ), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n246), .c(new_n211), .d(new_n243), .o1(new_n248));
  aoi112aa1n02x5               g153(.a(new_n247), .b(new_n246), .c(new_n211), .d(new_n243), .o1(new_n249));
  norb02aa1n03x4               g154(.a(new_n248), .b(new_n249), .out0(\s[21] ));
  xorc02aa1n12x5               g155(.a(\a[22] ), .b(\b[21] ), .out0(new_n251));
  nor042aa1n03x5               g156(.a(\b[20] ), .b(\a[21] ), .o1(new_n252));
  norp02aa1n02x5               g157(.a(new_n251), .b(new_n252), .o1(new_n253));
  inv000aa1n03x5               g158(.a(new_n252), .o1(new_n254));
  nand42aa1n02x5               g159(.a(new_n248), .b(new_n254), .o1(new_n255));
  aoi022aa1n02x7               g160(.a(new_n255), .b(new_n251), .c(new_n248), .d(new_n253), .o1(\s[22] ));
  nand22aa1n09x5               g161(.a(new_n251), .b(new_n247), .o1(new_n257));
  nona22aa1n03x5               g162(.a(new_n211), .b(new_n242), .c(new_n257), .out0(new_n258));
  nona22aa1n09x5               g163(.a(new_n239), .b(new_n244), .c(new_n223), .out0(new_n259));
  oaoi03aa1n02x5               g164(.a(\a[22] ), .b(\b[21] ), .c(new_n254), .o1(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  aoai13aa1n12x5               g166(.a(new_n261), .b(new_n257), .c(new_n259), .d(new_n245), .o1(new_n262));
  inv000aa1n02x5               g167(.a(new_n262), .o1(new_n263));
  xorc02aa1n02x5               g168(.a(\a[23] ), .b(\b[22] ), .out0(new_n264));
  xnbna2aa1n03x5               g169(.a(new_n264), .b(new_n258), .c(new_n263), .out0(\s[23] ));
  aob012aa1n03x5               g170(.a(new_n264), .b(new_n258), .c(new_n263), .out0(new_n266));
  xorc02aa1n02x5               g171(.a(\a[24] ), .b(\b[23] ), .out0(new_n267));
  norp02aa1n02x5               g172(.a(\b[22] ), .b(\a[23] ), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n267), .b(new_n268), .o1(new_n269));
  inv040aa1n02x5               g174(.a(new_n257), .o1(new_n270));
  aoi013aa1n03x5               g175(.a(new_n262), .b(new_n211), .c(new_n243), .d(new_n270), .o1(new_n271));
  oaoi03aa1n03x5               g176(.a(\a[23] ), .b(\b[22] ), .c(new_n271), .o1(new_n272));
  aoi022aa1n03x5               g177(.a(new_n272), .b(new_n267), .c(new_n266), .d(new_n269), .o1(\s[24] ));
  inv000aa1d42x5               g178(.a(\a[23] ), .o1(new_n274));
  inv040aa1d32x5               g179(.a(\a[24] ), .o1(new_n275));
  xroi22aa1d06x4               g180(.a(new_n274), .b(\b[22] ), .c(new_n275), .d(\b[23] ), .out0(new_n276));
  nano32aa1n02x5               g181(.a(new_n242), .b(new_n276), .c(new_n247), .d(new_n251), .out0(new_n277));
  nand02aa1d06x5               g182(.a(new_n211), .b(new_n277), .o1(new_n278));
  inv000aa1d42x5               g183(.a(\b[23] ), .o1(new_n279));
  tech160nm_fioaoi03aa1n03p5x5 g184(.a(new_n275), .b(new_n279), .c(new_n268), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n280), .o1(new_n281));
  tech160nm_fiaoi012aa1n04x5   g186(.a(new_n281), .b(new_n262), .c(new_n276), .o1(new_n282));
  norp02aa1n24x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  and002aa1n03x5               g188(.a(\b[24] ), .b(\a[25] ), .o(new_n284));
  nor042aa1n03x5               g189(.a(new_n284), .b(new_n283), .o1(new_n285));
  aob012aa1n03x5               g190(.a(new_n285), .b(new_n278), .c(new_n282), .out0(new_n286));
  aoi112aa1n02x5               g191(.a(new_n285), .b(new_n281), .c(new_n262), .d(new_n276), .o1(new_n287));
  aobi12aa1n02x7               g192(.a(new_n286), .b(new_n287), .c(new_n278), .out0(\s[25] ));
  xorc02aa1n12x5               g193(.a(\a[26] ), .b(\b[25] ), .out0(new_n289));
  norp02aa1n02x5               g194(.a(new_n289), .b(new_n283), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n283), .o1(new_n291));
  aoai13aa1n02x5               g196(.a(new_n291), .b(new_n284), .c(new_n278), .d(new_n282), .o1(new_n292));
  aoi022aa1n03x5               g197(.a(new_n292), .b(new_n289), .c(new_n286), .d(new_n290), .o1(\s[26] ));
  and002aa1n02x5               g198(.a(new_n289), .b(new_n285), .o(new_n294));
  aoai13aa1n09x5               g199(.a(new_n294), .b(new_n281), .c(new_n262), .d(new_n276), .o1(new_n295));
  nor042aa1n03x5               g200(.a(\b[26] ), .b(\a[27] ), .o1(new_n296));
  and002aa1n06x5               g201(.a(\b[26] ), .b(\a[27] ), .o(new_n297));
  nor042aa1n03x5               g202(.a(new_n297), .b(new_n296), .o1(new_n298));
  nano32aa1n02x5               g203(.a(new_n242), .b(new_n294), .c(new_n270), .d(new_n276), .out0(new_n299));
  oao003aa1n02x5               g204(.a(\a[26] ), .b(\b[25] ), .c(new_n291), .carry(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  aoi112aa1n02x5               g206(.a(new_n301), .b(new_n298), .c(new_n211), .d(new_n299), .o1(new_n302));
  aoi012aa1n09x5               g207(.a(new_n301), .b(new_n211), .c(new_n299), .o1(new_n303));
  nand42aa1n02x5               g208(.a(new_n303), .b(new_n295), .o1(new_n304));
  aoi022aa1n02x7               g209(.a(new_n304), .b(new_n298), .c(new_n295), .d(new_n302), .o1(\s[27] ));
  aoai13aa1n03x5               g210(.a(new_n276), .b(new_n260), .c(new_n246), .d(new_n270), .o1(new_n306));
  aobi12aa1n06x5               g211(.a(new_n294), .b(new_n306), .c(new_n280), .out0(new_n307));
  inv000aa1d42x5               g212(.a(new_n297), .o1(new_n308));
  nona23aa1n03x5               g213(.a(new_n294), .b(new_n276), .c(new_n242), .d(new_n257), .out0(new_n309));
  aoai13aa1n04x5               g214(.a(new_n300), .b(new_n309), .c(new_n202), .d(new_n210), .o1(new_n310));
  oai012aa1n02x5               g215(.a(new_n308), .b(new_n310), .c(new_n307), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n296), .o1(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n297), .c(new_n303), .d(new_n295), .o1(new_n313));
  xorc02aa1n02x5               g218(.a(\a[28] ), .b(\b[27] ), .out0(new_n314));
  norp02aa1n02x5               g219(.a(new_n314), .b(new_n296), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n313), .b(new_n314), .c(new_n311), .d(new_n315), .o1(\s[28] ));
  and002aa1n02x5               g221(.a(new_n314), .b(new_n298), .o(new_n317));
  oai012aa1n02x5               g222(.a(new_n317), .b(new_n310), .c(new_n307), .o1(new_n318));
  inv040aa1n03x5               g223(.a(new_n317), .o1(new_n319));
  oao003aa1n02x5               g224(.a(\a[28] ), .b(\b[27] ), .c(new_n312), .carry(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n303), .d(new_n295), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n320), .b(new_n322), .out0(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g230(.a(new_n314), .b(new_n322), .c(new_n298), .o(new_n326));
  oai012aa1n02x5               g231(.a(new_n326), .b(new_n310), .c(new_n307), .o1(new_n327));
  inv000aa1n02x5               g232(.a(new_n326), .o1(new_n328));
  oao003aa1n02x5               g233(.a(\a[29] ), .b(\b[28] ), .c(new_n320), .carry(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n328), .c(new_n303), .d(new_n295), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[30] ), .b(\b[29] ), .out0(new_n331));
  norb02aa1n02x5               g236(.a(new_n329), .b(new_n331), .out0(new_n332));
  aoi022aa1n03x5               g237(.a(new_n330), .b(new_n331), .c(new_n327), .d(new_n332), .o1(\s[30] ));
  nano22aa1n02x5               g238(.a(new_n319), .b(new_n322), .c(new_n331), .out0(new_n334));
  oai012aa1n02x5               g239(.a(new_n334), .b(new_n310), .c(new_n307), .o1(new_n335));
  xorc02aa1n02x5               g240(.a(\a[31] ), .b(\b[30] ), .out0(new_n336));
  and002aa1n02x5               g241(.a(\b[29] ), .b(\a[30] ), .o(new_n337));
  oabi12aa1n02x5               g242(.a(new_n336), .b(\a[30] ), .c(\b[29] ), .out0(new_n338));
  oab012aa1n02x4               g243(.a(new_n338), .b(new_n329), .c(new_n337), .out0(new_n339));
  inv000aa1n02x5               g244(.a(new_n334), .o1(new_n340));
  oao003aa1n02x5               g245(.a(\a[30] ), .b(\b[29] ), .c(new_n329), .carry(new_n341));
  aoai13aa1n03x5               g246(.a(new_n341), .b(new_n340), .c(new_n303), .d(new_n295), .o1(new_n342));
  aoi022aa1n03x5               g247(.a(new_n342), .b(new_n336), .c(new_n335), .d(new_n339), .o1(\s[31] ));
  xnbna2aa1n03x5               g248(.a(new_n135), .b(new_n101), .c(new_n99), .out0(\s[3] ));
  xorc02aa1n02x5               g249(.a(\a[4] ), .b(\b[3] ), .out0(new_n345));
  aoi112aa1n02x5               g250(.a(new_n102), .b(new_n345), .c(new_n134), .d(new_n135), .o1(new_n346));
  aob012aa1n02x5               g251(.a(new_n107), .b(\b[3] ), .c(\a[4] ), .out0(new_n347));
  oab012aa1n02x4               g252(.a(new_n346), .b(new_n347), .c(new_n105), .out0(\s[4] ));
  xnrb03aa1n02x5               g253(.a(new_n347), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  tech160nm_fioaoi03aa1n03p5x5 g254(.a(\a[5] ), .b(\b[4] ), .c(new_n347), .o1(new_n350));
  xorb03aa1n02x5               g255(.a(new_n350), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g256(.a(new_n117), .o1(new_n352));
  norb02aa1n02x5               g257(.a(new_n116), .b(new_n115), .out0(new_n353));
  norb02aa1n02x5               g258(.a(new_n120), .b(new_n117), .out0(new_n354));
  nanp02aa1n02x5               g259(.a(new_n350), .b(new_n354), .o1(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n353), .b(new_n355), .c(new_n352), .out0(\s[7] ));
  orn002aa1n02x5               g261(.a(\a[7] ), .b(\b[6] ), .o(new_n357));
  aoai13aa1n02x5               g262(.a(new_n353), .b(new_n117), .c(new_n350), .d(new_n120), .o1(new_n358));
  xnbna2aa1n03x5               g263(.a(new_n123), .b(new_n358), .c(new_n357), .out0(\s[8] ));
  xnbna2aa1n03x5               g264(.a(new_n128), .b(new_n159), .c(new_n160), .out0(\s[9] ));
endmodule


