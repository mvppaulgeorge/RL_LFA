// Benchmark "adder" written by ABC on Thu Jul 18 09:48:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n144, new_n145, new_n146, new_n147,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n168, new_n169, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n338, new_n339, new_n340, new_n342, new_n343, new_n345, new_n346,
    new_n347, new_n349, new_n350, new_n351, new_n353, new_n354, new_n356,
    new_n357;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nand02aa1d24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[6] ), .b(\a[7] ), .o1(new_n98));
  nor042aa1n04x5               g003(.a(\b[5] ), .b(\a[6] ), .o1(new_n99));
  nor002aa1d32x5               g004(.a(\b[4] ), .b(\a[5] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[5] ), .b(\a[6] ), .o1(new_n101));
  aoai13aa1n12x5               g006(.a(new_n98), .b(new_n99), .c(new_n100), .d(new_n101), .o1(new_n102));
  nor002aa1n20x5               g007(.a(\b[6] ), .b(\a[7] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[7] ), .b(\a[8] ), .o1(new_n104));
  norp02aa1n24x5               g009(.a(new_n104), .b(new_n103), .o1(new_n105));
  aoi022aa1d18x5               g010(.a(new_n102), .b(new_n105), .c(\b[7] ), .d(\a[8] ), .o1(new_n106));
  orn002aa1n24x5               g011(.a(\a[2] ), .b(\b[1] ), .o(new_n107));
  nand22aa1n12x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  aoi012aa1d24x5               g013(.a(new_n108), .b(\a[2] ), .c(\b[1] ), .o1(new_n109));
  nand02aa1d10x5               g014(.a(\b[1] ), .b(\a[2] ), .o1(new_n110));
  nand02aa1d28x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nor002aa1d32x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanb03aa1d24x5               g017(.a(new_n112), .b(new_n110), .c(new_n111), .out0(new_n113));
  inv040aa1d32x5               g018(.a(\a[4] ), .o1(new_n114));
  inv040aa1d30x5               g019(.a(\b[3] ), .o1(new_n115));
  aoi012aa1n09x5               g020(.a(new_n112), .b(new_n114), .c(new_n115), .o1(new_n116));
  aoai13aa1n12x5               g021(.a(new_n116), .b(new_n113), .c(new_n107), .d(new_n109), .o1(new_n117));
  nand42aa1n06x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  inv040aa1n02x5               g023(.a(new_n104), .o1(new_n119));
  oai112aa1n04x5               g024(.a(new_n119), .b(new_n118), .c(\b[6] ), .d(\a[7] ), .o1(new_n120));
  oai022aa1n09x5               g025(.a(new_n114), .b(new_n115), .c(\b[4] ), .d(\a[5] ), .o1(new_n121));
  nand02aa1n08x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  aoi022aa1d24x5               g027(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n123));
  oai112aa1n06x5               g028(.a(new_n123), .b(new_n122), .c(\b[5] ), .d(\a[6] ), .o1(new_n124));
  nor043aa1n09x5               g029(.a(new_n124), .b(new_n120), .c(new_n121), .o1(new_n125));
  nor042aa1n04x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n06x4               g031(.a(new_n97), .b(new_n126), .out0(new_n127));
  inv040aa1n02x5               g032(.a(new_n127), .o1(new_n128));
  aoi112aa1n09x5               g033(.a(new_n128), .b(new_n106), .c(new_n125), .d(new_n117), .o1(new_n129));
  inv000aa1n06x5               g034(.a(new_n129), .o1(new_n130));
  xnrc02aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n130), .c(new_n97), .out0(\s[10] ));
  inv000aa1n02x5               g037(.a(new_n131), .o1(new_n133));
  aoai13aa1n06x5               g038(.a(new_n133), .b(new_n129), .c(\a[9] ), .d(\b[8] ), .o1(new_n134));
  nor002aa1d32x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand42aa1d28x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  inv000aa1d42x5               g042(.a(\b[9] ), .o1(new_n138));
  oaib12aa1n03x5               g043(.a(new_n134), .b(new_n138), .c(\a[10] ), .out0(new_n139));
  inv000aa1d42x5               g044(.a(\a[10] ), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n135), .o1(new_n141));
  oai112aa1n02x5               g046(.a(new_n141), .b(new_n136), .c(new_n138), .d(new_n140), .o1(new_n142));
  aboi22aa1n03x5               g047(.a(new_n142), .b(new_n134), .c(new_n139), .d(new_n137), .out0(\s[11] ));
  nanb02aa1n03x5               g048(.a(new_n142), .b(new_n134), .out0(new_n144));
  norp02aa1n24x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand42aa1n20x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  norb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n147), .b(new_n144), .c(new_n141), .out0(\s[12] ));
  nona23aa1n09x5               g053(.a(new_n146), .b(new_n136), .c(new_n135), .d(new_n145), .out0(new_n149));
  nor043aa1n02x5               g054(.a(new_n149), .b(new_n128), .c(new_n131), .o1(new_n150));
  aoai13aa1n06x5               g055(.a(new_n150), .b(new_n106), .c(new_n125), .d(new_n117), .o1(new_n151));
  oaoi03aa1n02x5               g056(.a(new_n140), .b(new_n138), .c(new_n126), .o1(new_n152));
  tech160nm_fiaoi012aa1n05x5   g057(.a(new_n145), .b(new_n135), .c(new_n146), .o1(new_n153));
  oai012aa1n02x7               g058(.a(new_n153), .b(new_n149), .c(new_n152), .o1(new_n154));
  nanb02aa1n06x5               g059(.a(new_n154), .b(new_n151), .out0(new_n155));
  nor002aa1n20x5               g060(.a(\b[12] ), .b(\a[13] ), .o1(new_n156));
  nand02aa1d24x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  norb02aa1n09x5               g062(.a(new_n157), .b(new_n156), .out0(new_n158));
  nano23aa1n03x7               g063(.a(new_n135), .b(new_n145), .c(new_n146), .d(new_n136), .out0(new_n159));
  oao003aa1n02x5               g064(.a(new_n140), .b(new_n138), .c(new_n126), .carry(new_n160));
  nand42aa1n02x5               g065(.a(new_n159), .b(new_n160), .o1(new_n161));
  inv000aa1n02x5               g066(.a(new_n158), .o1(new_n162));
  and003aa1n02x5               g067(.a(new_n161), .b(new_n162), .c(new_n153), .o(new_n163));
  aoi022aa1n02x5               g068(.a(new_n155), .b(new_n158), .c(new_n151), .d(new_n163), .o1(\s[13] ));
  nor002aa1n06x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nand02aa1d24x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  norb02aa1n03x5               g071(.a(new_n166), .b(new_n165), .out0(new_n167));
  aoi112aa1n02x5               g072(.a(new_n156), .b(new_n167), .c(new_n155), .d(new_n158), .o1(new_n168));
  aoai13aa1n02x5               g073(.a(new_n167), .b(new_n156), .c(new_n155), .d(new_n157), .o1(new_n169));
  norb02aa1n03x4               g074(.a(new_n169), .b(new_n168), .out0(\s[14] ));
  nano23aa1n06x5               g075(.a(new_n156), .b(new_n165), .c(new_n166), .d(new_n157), .out0(new_n171));
  ao0012aa1n12x5               g076(.a(new_n165), .b(new_n156), .c(new_n166), .o(new_n172));
  nor002aa1n20x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nand42aa1n10x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n12x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  aoai13aa1n06x5               g080(.a(new_n175), .b(new_n172), .c(new_n155), .d(new_n171), .o1(new_n176));
  aoi112aa1n02x7               g081(.a(new_n175), .b(new_n172), .c(new_n155), .d(new_n171), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(\s[15] ));
  nor042aa1n09x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  nand42aa1d28x5               g084(.a(\b[15] ), .b(\a[16] ), .o1(new_n180));
  norb02aa1n03x5               g085(.a(new_n180), .b(new_n179), .out0(new_n181));
  aoib12aa1n02x5               g086(.a(new_n173), .b(new_n180), .c(new_n179), .out0(new_n182));
  oaih12aa1n02x5               g087(.a(new_n176), .b(\b[14] ), .c(\a[15] ), .o1(new_n183));
  aoi022aa1n02x7               g088(.a(new_n183), .b(new_n181), .c(new_n176), .d(new_n182), .o1(\s[16] ));
  aoi012aa1d18x5               g089(.a(new_n106), .b(new_n125), .c(new_n117), .o1(new_n185));
  nano32aa1n03x7               g090(.a(new_n162), .b(new_n181), .c(new_n167), .d(new_n175), .out0(new_n186));
  nand02aa1n03x5               g091(.a(new_n186), .b(new_n150), .o1(new_n187));
  nano23aa1d15x5               g092(.a(new_n173), .b(new_n179), .c(new_n180), .d(new_n174), .out0(new_n188));
  nand02aa1n04x5               g093(.a(new_n188), .b(new_n172), .o1(new_n189));
  aoi012aa1d24x5               g094(.a(new_n179), .b(new_n173), .c(new_n180), .o1(new_n190));
  nanp02aa1n02x5               g095(.a(new_n189), .b(new_n190), .o1(new_n191));
  aoi012aa1n06x5               g096(.a(new_n191), .b(new_n154), .c(new_n186), .o1(new_n192));
  oai012aa1d24x5               g097(.a(new_n192), .b(new_n185), .c(new_n187), .o1(new_n193));
  xorc02aa1n12x5               g098(.a(\a[17] ), .b(\b[16] ), .out0(new_n194));
  inv000aa1n06x5               g099(.a(new_n106), .o1(new_n195));
  nanp02aa1n02x5               g100(.a(new_n109), .b(new_n107), .o1(new_n196));
  nano22aa1n02x4               g101(.a(new_n112), .b(new_n110), .c(new_n111), .out0(new_n197));
  aobi12aa1n02x5               g102(.a(new_n116), .b(new_n196), .c(new_n197), .out0(new_n198));
  norb03aa1n02x7               g103(.a(new_n118), .b(new_n104), .c(new_n103), .out0(new_n199));
  oai012aa1n02x5               g104(.a(new_n122), .b(\b[5] ), .c(\a[6] ), .o1(new_n200));
  nona23aa1n03x5               g105(.a(new_n199), .b(new_n123), .c(new_n121), .d(new_n200), .out0(new_n201));
  tech160nm_fioai012aa1n05x5   g106(.a(new_n195), .b(new_n198), .c(new_n201), .o1(new_n202));
  nanp02aa1n02x5               g107(.a(new_n188), .b(new_n171), .o1(new_n203));
  nano32aa1n03x7               g108(.a(new_n203), .b(new_n133), .c(new_n159), .d(new_n127), .out0(new_n204));
  nanb03aa1n02x5               g109(.a(new_n194), .b(new_n189), .c(new_n190), .out0(new_n205));
  aoi122aa1n02x5               g110(.a(new_n205), .b(new_n154), .c(new_n186), .d(new_n202), .e(new_n204), .o1(new_n206));
  aoi012aa1n02x5               g111(.a(new_n206), .b(new_n193), .c(new_n194), .o1(\s[17] ));
  inv000aa1d42x5               g112(.a(\a[17] ), .o1(new_n208));
  nanb02aa1n02x5               g113(.a(\b[16] ), .b(new_n208), .out0(new_n209));
  aobi12aa1n06x5               g114(.a(new_n190), .b(new_n188), .c(new_n172), .out0(new_n210));
  aoai13aa1n03x5               g115(.a(new_n210), .b(new_n203), .c(new_n161), .d(new_n153), .o1(new_n211));
  aoai13aa1n02x5               g116(.a(new_n194), .b(new_n211), .c(new_n202), .d(new_n204), .o1(new_n212));
  xorc02aa1n12x5               g117(.a(\a[18] ), .b(\b[17] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n212), .c(new_n209), .out0(\s[18] ));
  inv000aa1d42x5               g119(.a(\a[18] ), .o1(new_n215));
  xroi22aa1d04x5               g120(.a(new_n208), .b(\b[16] ), .c(new_n215), .d(\b[17] ), .out0(new_n216));
  oaoi03aa1n02x5               g121(.a(\a[18] ), .b(\b[17] ), .c(new_n209), .o1(new_n217));
  nor042aa1d18x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nand02aa1d24x5               g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  norb02aa1n15x5               g124(.a(new_n219), .b(new_n218), .out0(new_n220));
  aoai13aa1n09x5               g125(.a(new_n220), .b(new_n217), .c(new_n193), .d(new_n216), .o1(new_n221));
  aoi112aa1n02x5               g126(.a(new_n220), .b(new_n217), .c(new_n193), .d(new_n216), .o1(new_n222));
  norb02aa1n03x4               g127(.a(new_n221), .b(new_n222), .out0(\s[19] ));
  xnrc02aa1n02x5               g128(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1d18x5               g129(.a(\b[19] ), .b(\a[20] ), .o1(new_n225));
  nand02aa1d28x5               g130(.a(\b[19] ), .b(\a[20] ), .o1(new_n226));
  norb02aa1n06x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  aoib12aa1n02x5               g132(.a(new_n218), .b(new_n226), .c(new_n225), .out0(new_n228));
  tech160nm_fioai012aa1n03p5x5 g133(.a(new_n221), .b(\b[18] ), .c(\a[19] ), .o1(new_n229));
  aoi022aa1n02x7               g134(.a(new_n229), .b(new_n227), .c(new_n221), .d(new_n228), .o1(\s[20] ));
  nano23aa1n06x5               g135(.a(new_n218), .b(new_n225), .c(new_n226), .d(new_n219), .out0(new_n231));
  nand23aa1n09x5               g136(.a(new_n231), .b(new_n194), .c(new_n213), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n232), .o1(new_n233));
  nor042aa1n02x5               g138(.a(\b[17] ), .b(\a[18] ), .o1(new_n234));
  aoi112aa1n09x5               g139(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n235));
  oai112aa1n06x5               g140(.a(new_n220), .b(new_n227), .c(new_n235), .d(new_n234), .o1(new_n236));
  tech160nm_fiaoi012aa1n03p5x5 g141(.a(new_n225), .b(new_n218), .c(new_n226), .o1(new_n237));
  nanp02aa1n02x5               g142(.a(new_n236), .b(new_n237), .o1(new_n238));
  xorc02aa1n12x5               g143(.a(\a[21] ), .b(\b[20] ), .out0(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n238), .c(new_n193), .d(new_n233), .o1(new_n240));
  nano22aa1n02x4               g145(.a(new_n239), .b(new_n236), .c(new_n237), .out0(new_n241));
  aobi12aa1n02x5               g146(.a(new_n241), .b(new_n193), .c(new_n233), .out0(new_n242));
  norb02aa1n03x4               g147(.a(new_n240), .b(new_n242), .out0(\s[21] ));
  xorc02aa1n03x5               g148(.a(\a[22] ), .b(\b[21] ), .out0(new_n244));
  inv000aa1d42x5               g149(.a(\a[21] ), .o1(new_n245));
  aoib12aa1n02x5               g150(.a(new_n244), .b(new_n245), .c(\b[20] ), .out0(new_n246));
  oaib12aa1n06x5               g151(.a(new_n240), .b(\b[20] ), .c(new_n245), .out0(new_n247));
  aoi022aa1n02x7               g152(.a(new_n247), .b(new_n244), .c(new_n240), .d(new_n246), .o1(\s[22] ));
  nand02aa1n03x5               g153(.a(new_n244), .b(new_n239), .o1(new_n249));
  nano32aa1n02x4               g154(.a(new_n249), .b(new_n231), .c(new_n213), .d(new_n194), .out0(new_n250));
  inv000aa1d42x5               g155(.a(\a[22] ), .o1(new_n251));
  aoi112aa1n02x5               g156(.a(\b[20] ), .b(\a[21] ), .c(\a[22] ), .d(\b[21] ), .o1(new_n252));
  aoib12aa1n06x5               g157(.a(new_n252), .b(new_n251), .c(\b[21] ), .out0(new_n253));
  aoai13aa1n06x5               g158(.a(new_n253), .b(new_n249), .c(new_n236), .d(new_n237), .o1(new_n254));
  xorc02aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n254), .c(new_n193), .d(new_n250), .o1(new_n256));
  xroi22aa1d04x5               g161(.a(new_n245), .b(\b[20] ), .c(new_n251), .d(\b[21] ), .out0(new_n257));
  nanb02aa1n02x5               g162(.a(new_n255), .b(new_n253), .out0(new_n258));
  aoi012aa1n02x5               g163(.a(new_n258), .b(new_n238), .c(new_n257), .o1(new_n259));
  aobi12aa1n02x5               g164(.a(new_n259), .b(new_n193), .c(new_n250), .out0(new_n260));
  norb02aa1n03x4               g165(.a(new_n256), .b(new_n260), .out0(\s[23] ));
  xorc02aa1n02x5               g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  norp02aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  norp02aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  inv000aa1d48x5               g169(.a(\a[23] ), .o1(new_n265));
  oaib12aa1n06x5               g170(.a(new_n256), .b(\b[22] ), .c(new_n265), .out0(new_n266));
  aoi022aa1n02x7               g171(.a(new_n266), .b(new_n262), .c(new_n256), .d(new_n264), .o1(\s[24] ));
  inv040aa1d32x5               g172(.a(\a[24] ), .o1(new_n268));
  xroi22aa1d06x4               g173(.a(new_n265), .b(\b[22] ), .c(new_n268), .d(\b[23] ), .out0(new_n269));
  nano22aa1n03x7               g174(.a(new_n232), .b(new_n257), .c(new_n269), .out0(new_n270));
  aob012aa1n02x5               g175(.a(new_n263), .b(\b[23] ), .c(\a[24] ), .out0(new_n271));
  oaib12aa1n02x5               g176(.a(new_n271), .b(\b[23] ), .c(new_n268), .out0(new_n272));
  tech160nm_fiao0012aa1n02p5x5 g177(.a(new_n272), .b(new_n254), .c(new_n269), .o(new_n273));
  xorc02aa1n02x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  aoai13aa1n09x5               g179(.a(new_n274), .b(new_n273), .c(new_n193), .d(new_n270), .o1(new_n275));
  aoi112aa1n02x5               g180(.a(new_n274), .b(new_n272), .c(new_n254), .d(new_n269), .o1(new_n276));
  aobi12aa1n02x5               g181(.a(new_n276), .b(new_n270), .c(new_n193), .out0(new_n277));
  norb02aa1n03x4               g182(.a(new_n275), .b(new_n277), .out0(\s[25] ));
  xorc02aa1n02x5               g183(.a(\a[26] ), .b(\b[25] ), .out0(new_n279));
  norp02aa1n02x5               g184(.a(\b[24] ), .b(\a[25] ), .o1(new_n280));
  norp02aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(\a[25] ), .o1(new_n282));
  oaib12aa1n06x5               g187(.a(new_n275), .b(\b[24] ), .c(new_n282), .out0(new_n283));
  aoi022aa1n02x7               g188(.a(new_n283), .b(new_n279), .c(new_n275), .d(new_n281), .o1(\s[26] ));
  inv000aa1d42x5               g189(.a(\a[26] ), .o1(new_n285));
  xroi22aa1d04x5               g190(.a(new_n282), .b(\b[24] ), .c(new_n285), .d(\b[25] ), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n272), .c(new_n254), .d(new_n269), .o1(new_n287));
  nano32aa1n03x7               g192(.a(new_n232), .b(new_n286), .c(new_n257), .d(new_n269), .out0(new_n288));
  aoai13aa1n06x5               g193(.a(new_n288), .b(new_n211), .c(new_n202), .d(new_n204), .o1(new_n289));
  inv000aa1d42x5               g194(.a(\b[25] ), .o1(new_n290));
  oaoi03aa1n12x5               g195(.a(new_n285), .b(new_n290), .c(new_n280), .o1(new_n291));
  nanp03aa1n06x5               g196(.a(new_n289), .b(new_n287), .c(new_n291), .o1(new_n292));
  xorc02aa1n12x5               g197(.a(\a[27] ), .b(\b[26] ), .out0(new_n293));
  inv000aa1d42x5               g198(.a(new_n291), .o1(new_n294));
  aoi112aa1n02x7               g199(.a(new_n293), .b(new_n294), .c(new_n193), .d(new_n288), .o1(new_n295));
  aoi022aa1n02x5               g200(.a(new_n295), .b(new_n287), .c(new_n292), .d(new_n293), .o1(\s[27] ));
  nanp02aa1n03x5               g201(.a(new_n292), .b(new_n293), .o1(new_n297));
  xorc02aa1n02x5               g202(.a(\a[28] ), .b(\b[27] ), .out0(new_n298));
  nor042aa1n09x5               g203(.a(\b[26] ), .b(\a[27] ), .o1(new_n299));
  norp02aa1n02x5               g204(.a(new_n298), .b(new_n299), .o1(new_n300));
  tech160nm_fiaoi012aa1n05x5   g205(.a(new_n294), .b(new_n193), .c(new_n288), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n299), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n293), .o1(new_n303));
  aoai13aa1n03x5               g208(.a(new_n302), .b(new_n303), .c(new_n301), .d(new_n287), .o1(new_n304));
  aoi022aa1n03x5               g209(.a(new_n304), .b(new_n298), .c(new_n297), .d(new_n300), .o1(\s[28] ));
  inv000aa1d42x5               g210(.a(\a[27] ), .o1(new_n306));
  inv000aa1d42x5               g211(.a(\a[28] ), .o1(new_n307));
  xroi22aa1d04x5               g212(.a(new_n306), .b(\b[26] ), .c(new_n307), .d(\b[27] ), .out0(new_n308));
  inv000aa1d42x5               g213(.a(new_n308), .o1(new_n309));
  aoi013aa1n02x4               g214(.a(new_n309), .b(new_n289), .c(new_n287), .d(new_n291), .o1(new_n310));
  tech160nm_fixorc02aa1n03p5x5 g215(.a(\a[29] ), .b(\b[28] ), .out0(new_n311));
  aob012aa1n02x5               g216(.a(new_n299), .b(\b[27] ), .c(\a[28] ), .out0(new_n312));
  inv000aa1d42x5               g217(.a(new_n311), .o1(new_n313));
  oai112aa1n02x5               g218(.a(new_n313), .b(new_n312), .c(\b[27] ), .d(\a[28] ), .o1(new_n314));
  tech160nm_fiaoi012aa1n05x5   g219(.a(new_n314), .b(new_n292), .c(new_n308), .o1(new_n315));
  oaib12aa1n06x5               g220(.a(new_n312), .b(\b[27] ), .c(new_n307), .out0(new_n316));
  oaoi13aa1n02x7               g221(.a(new_n315), .b(new_n311), .c(new_n316), .d(new_n310), .o1(\s[29] ));
  xorb03aa1n02x5               g222(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n03x7               g223(.a(new_n313), .b(new_n293), .c(new_n298), .out0(new_n319));
  inv000aa1n02x5               g224(.a(new_n319), .o1(new_n320));
  aoi013aa1n03x5               g225(.a(new_n320), .b(new_n289), .c(new_n287), .d(new_n291), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  inv000aa1d42x5               g227(.a(\a[29] ), .o1(new_n323));
  oaib12aa1n06x5               g228(.a(new_n316), .b(new_n323), .c(\b[28] ), .out0(new_n324));
  aoib12aa1n02x5               g229(.a(new_n322), .b(new_n323), .c(\b[28] ), .out0(new_n325));
  nanp02aa1n02x5               g230(.a(new_n325), .b(new_n324), .o1(new_n326));
  tech160nm_fiaoi012aa1n05x5   g231(.a(new_n326), .b(new_n292), .c(new_n319), .o1(new_n327));
  oaib12aa1n02x5               g232(.a(new_n324), .b(\b[28] ), .c(new_n323), .out0(new_n328));
  oaoi13aa1n02x7               g233(.a(new_n327), .b(new_n322), .c(new_n328), .d(new_n321), .o1(\s[30] ));
  nanp03aa1n02x5               g234(.a(new_n308), .b(new_n311), .c(new_n322), .o1(new_n330));
  nanb02aa1n02x5               g235(.a(new_n330), .b(new_n292), .out0(new_n331));
  xorc02aa1n02x5               g236(.a(\a[31] ), .b(\b[30] ), .out0(new_n332));
  oai122aa1n06x5               g237(.a(new_n324), .b(\a[30] ), .c(\b[29] ), .d(\a[29] ), .e(\b[28] ), .o1(new_n333));
  aob012aa1n03x5               g238(.a(new_n333), .b(\b[29] ), .c(\a[30] ), .out0(new_n334));
  norb02aa1n02x5               g239(.a(new_n334), .b(new_n332), .out0(new_n335));
  aoai13aa1n03x5               g240(.a(new_n334), .b(new_n330), .c(new_n301), .d(new_n287), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n336), .b(new_n332), .c(new_n331), .d(new_n335), .o1(\s[31] ));
  aoi012aa1n02x5               g242(.a(new_n113), .b(new_n107), .c(new_n109), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n112), .o1(new_n339));
  aoi022aa1n02x5               g244(.a(new_n196), .b(new_n110), .c(new_n339), .d(new_n111), .o1(new_n340));
  norp02aa1n02x5               g245(.a(new_n340), .b(new_n338), .o1(\s[3] ));
  inv000aa1n03x5               g246(.a(new_n338), .o1(new_n342));
  xorc02aa1n02x5               g247(.a(\a[4] ), .b(\b[3] ), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n342), .c(new_n339), .out0(\s[4] ));
  nanb03aa1n06x5               g249(.a(new_n121), .b(new_n117), .c(new_n122), .out0(new_n345));
  oaib12aa1n02x5               g250(.a(new_n117), .b(new_n115), .c(\a[4] ), .out0(new_n346));
  nanb02aa1n02x5               g251(.a(new_n100), .b(new_n122), .out0(new_n347));
  aobi12aa1n02x5               g252(.a(new_n345), .b(new_n347), .c(new_n346), .out0(\s[5] ));
  inv000aa1d42x5               g253(.a(new_n100), .o1(new_n349));
  norb02aa1n02x5               g254(.a(new_n101), .b(new_n99), .out0(new_n350));
  nona23aa1n06x5               g255(.a(new_n345), .b(new_n101), .c(new_n99), .d(new_n100), .out0(new_n351));
  aoai13aa1n02x5               g256(.a(new_n351), .b(new_n350), .c(new_n349), .d(new_n345), .o1(\s[6] ));
  inv000aa1d42x5               g257(.a(new_n103), .o1(new_n353));
  aoi022aa1n02x5               g258(.a(new_n351), .b(new_n101), .c(new_n98), .d(new_n353), .o1(new_n354));
  aoi013aa1n02x4               g259(.a(new_n354), .b(new_n351), .c(new_n123), .d(new_n353), .o1(\s[7] ));
  nanp03aa1n03x5               g260(.a(new_n351), .b(new_n353), .c(new_n123), .o1(new_n356));
  norb02aa1n02x5               g261(.a(new_n118), .b(new_n104), .out0(new_n357));
  xnbna2aa1n03x5               g262(.a(new_n357), .b(new_n356), .c(new_n353), .out0(\s[8] ));
  oaib12aa1n02x5               g263(.a(new_n130), .b(new_n185), .c(new_n128), .out0(\s[9] ));
endmodule


