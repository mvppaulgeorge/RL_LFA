// Benchmark "adder" written by ABC on Wed Jul 17 16:16:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n326, new_n327, new_n329, new_n330, new_n331, new_n333,
    new_n334, new_n335, new_n337, new_n338;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\b[8] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\a[9] ), .b(new_n97), .out0(new_n98));
  nand02aa1d28x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(new_n99), .o1(new_n100));
  oaoi03aa1n09x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand02aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor002aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nano23aa1n06x5               g010(.a(new_n102), .b(new_n104), .c(new_n105), .d(new_n103), .out0(new_n106));
  oa0012aa1n06x5               g011(.a(new_n103), .b(new_n104), .c(new_n102), .o(new_n107));
  aoi012aa1n06x5               g012(.a(new_n107), .b(new_n106), .c(new_n101), .o1(new_n108));
  nor002aa1n03x5               g013(.a(\b[6] ), .b(\a[7] ), .o1(new_n109));
  nand42aa1n16x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nor042aa1n04x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand42aa1n03x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nano23aa1n02x4               g017(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n113));
  nor042aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand02aa1d28x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  norb02aa1n06x4               g020(.a(new_n115), .b(new_n114), .out0(new_n116));
  tech160nm_fixorc02aa1n04x5   g021(.a(\a[8] ), .b(\b[7] ), .out0(new_n117));
  nand23aa1n03x5               g022(.a(new_n113), .b(new_n116), .c(new_n117), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[8] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[7] ), .o1(new_n120));
  inv000aa1n02x5               g025(.a(new_n109), .o1(new_n121));
  aoai13aa1n06x5               g026(.a(new_n110), .b(new_n114), .c(new_n111), .d(new_n115), .o1(new_n122));
  nand22aa1n03x5               g027(.a(new_n122), .b(new_n121), .o1(new_n123));
  oaoi03aa1n12x5               g028(.a(new_n119), .b(new_n120), .c(new_n123), .o1(new_n124));
  oai012aa1n12x5               g029(.a(new_n124), .b(new_n108), .c(new_n118), .o1(new_n125));
  xnrc02aa1n12x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  inv000aa1d42x5               g031(.a(new_n126), .o1(new_n127));
  nanp02aa1n02x5               g032(.a(new_n125), .b(new_n127), .o1(new_n128));
  xorc02aa1n12x5               g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  xnbna2aa1n03x5               g034(.a(new_n129), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g035(.a(\a[10] ), .o1(new_n131));
  xroi22aa1d04x5               g036(.a(new_n131), .b(\b[9] ), .c(new_n97), .d(\a[9] ), .out0(new_n132));
  oaoi03aa1n02x5               g037(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n133));
  xorc02aa1n12x5               g038(.a(\a[11] ), .b(\b[10] ), .out0(new_n134));
  aoai13aa1n06x5               g039(.a(new_n134), .b(new_n133), .c(new_n125), .d(new_n132), .o1(new_n135));
  aoi112aa1n02x5               g040(.a(new_n134), .b(new_n133), .c(new_n125), .d(new_n132), .o1(new_n136));
  norb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(\s[11] ));
  inv000aa1d42x5               g042(.a(\a[11] ), .o1(new_n138));
  nanb02aa1d24x5               g043(.a(\b[10] ), .b(new_n138), .out0(new_n139));
  xorc02aa1n12x5               g044(.a(\a[12] ), .b(\b[11] ), .out0(new_n140));
  xnbna2aa1n03x5               g045(.a(new_n140), .b(new_n135), .c(new_n139), .out0(\s[12] ));
  nona23aa1n03x5               g046(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n142));
  nano22aa1n03x7               g047(.a(new_n142), .b(new_n117), .c(new_n116), .out0(new_n143));
  aoai13aa1n06x5               g048(.a(new_n143), .b(new_n107), .c(new_n101), .d(new_n106), .o1(new_n144));
  nano32aa1d12x5               g049(.a(new_n126), .b(new_n140), .c(new_n129), .d(new_n134), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  nor042aa1n02x5               g051(.a(\b[9] ), .b(\a[10] ), .o1(new_n147));
  aoi112aa1n09x5               g052(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n148));
  oai112aa1n06x5               g053(.a(new_n134), .b(new_n140), .c(new_n148), .d(new_n147), .o1(new_n149));
  oao003aa1n09x5               g054(.a(\a[12] ), .b(\b[11] ), .c(new_n139), .carry(new_n150));
  nand22aa1n12x5               g055(.a(new_n149), .b(new_n150), .o1(new_n151));
  inv000aa1d42x5               g056(.a(new_n151), .o1(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n146), .c(new_n144), .d(new_n124), .o1(new_n153));
  xorc02aa1n12x5               g058(.a(\a[13] ), .b(\b[12] ), .out0(new_n154));
  aoi112aa1n02x5               g059(.a(new_n154), .b(new_n151), .c(new_n125), .d(new_n145), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n155), .b(new_n153), .c(new_n154), .o1(\s[13] ));
  nor042aa1d18x5               g061(.a(\b[12] ), .b(\a[13] ), .o1(new_n157));
  inv030aa1n06x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n03x5               g063(.a(new_n154), .b(new_n151), .c(new_n125), .d(new_n145), .o1(new_n159));
  xorc02aa1n12x5               g064(.a(\a[14] ), .b(\b[13] ), .out0(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n159), .c(new_n158), .out0(\s[14] ));
  nand02aa1n06x5               g066(.a(new_n160), .b(new_n154), .o1(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n151), .c(new_n125), .d(new_n145), .o1(new_n164));
  oaoi03aa1n12x5               g069(.a(\a[14] ), .b(\b[13] ), .c(new_n158), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  xorc02aa1n12x5               g071(.a(\a[15] ), .b(\b[14] ), .out0(new_n167));
  xnbna2aa1n03x5               g072(.a(new_n167), .b(new_n164), .c(new_n166), .out0(\s[15] ));
  aoai13aa1n02x5               g073(.a(new_n167), .b(new_n165), .c(new_n153), .d(new_n163), .o1(new_n169));
  xorc02aa1n12x5               g074(.a(\a[16] ), .b(\b[15] ), .out0(new_n170));
  nor042aa1n06x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  norp02aa1n02x5               g076(.a(new_n170), .b(new_n171), .o1(new_n172));
  inv000aa1d42x5               g077(.a(new_n171), .o1(new_n173));
  inv000aa1d42x5               g078(.a(new_n167), .o1(new_n174));
  aoai13aa1n02x7               g079(.a(new_n173), .b(new_n174), .c(new_n164), .d(new_n166), .o1(new_n175));
  aoi022aa1n02x5               g080(.a(new_n175), .b(new_n170), .c(new_n169), .d(new_n172), .o1(\s[16] ));
  xnrc02aa1n02x5               g081(.a(\b[12] ), .b(\a[13] ), .out0(new_n177));
  xnrc02aa1n02x5               g082(.a(\b[13] ), .b(\a[14] ), .out0(new_n178));
  nona23aa1n08x5               g083(.a(new_n167), .b(new_n170), .c(new_n178), .d(new_n177), .out0(new_n179));
  nano32aa1n03x7               g084(.a(new_n179), .b(new_n132), .c(new_n134), .d(new_n140), .out0(new_n180));
  nanp02aa1n02x5               g085(.a(new_n125), .b(new_n180), .o1(new_n181));
  nano22aa1n03x7               g086(.a(new_n162), .b(new_n167), .c(new_n170), .out0(new_n182));
  nand02aa1d04x5               g087(.a(new_n145), .b(new_n182), .o1(new_n183));
  nand43aa1n02x5               g088(.a(new_n165), .b(new_n167), .c(new_n170), .o1(new_n184));
  oaoi03aa1n03x5               g089(.a(\a[16] ), .b(\b[15] ), .c(new_n173), .o1(new_n185));
  nanb02aa1n03x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  aoi012aa1n06x5               g091(.a(new_n186), .b(new_n151), .c(new_n182), .o1(new_n187));
  aoai13aa1n12x5               g092(.a(new_n187), .b(new_n183), .c(new_n144), .d(new_n124), .o1(new_n188));
  xorc02aa1n02x5               g093(.a(\a[17] ), .b(\b[16] ), .out0(new_n189));
  aoi112aa1n02x5               g094(.a(new_n189), .b(new_n186), .c(new_n151), .d(new_n182), .o1(new_n190));
  aoi022aa1n02x5               g095(.a(new_n188), .b(new_n189), .c(new_n181), .d(new_n190), .o1(\s[17] ));
  tech160nm_ficinv00aa1n08x5   g096(.clk(\a[17] ), .clkout(new_n192));
  nanb02aa1n12x5               g097(.a(\b[16] ), .b(new_n192), .out0(new_n193));
  aoi013aa1n03x5               g098(.a(new_n185), .b(new_n165), .c(new_n167), .d(new_n170), .o1(new_n194));
  aoai13aa1n06x5               g099(.a(new_n194), .b(new_n179), .c(new_n149), .d(new_n150), .o1(new_n195));
  aoai13aa1n03x5               g100(.a(new_n189), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n196));
  xorc02aa1n02x5               g101(.a(\a[18] ), .b(\b[17] ), .out0(new_n197));
  xnbna2aa1n03x5               g102(.a(new_n197), .b(new_n196), .c(new_n193), .out0(\s[18] ));
  inv000aa1d42x5               g103(.a(\a[18] ), .o1(new_n199));
  xroi22aa1d04x5               g104(.a(new_n192), .b(\b[16] ), .c(new_n199), .d(\b[17] ), .out0(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n201));
  oaoi03aa1n12x5               g106(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n202));
  inv000aa1d42x5               g107(.a(new_n202), .o1(new_n203));
  xorc02aa1n12x5               g108(.a(\a[19] ), .b(\b[18] ), .out0(new_n204));
  xnbna2aa1n03x5               g109(.a(new_n204), .b(new_n201), .c(new_n203), .out0(\s[19] ));
  xnrc02aa1n02x5               g110(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g111(.a(new_n204), .b(new_n202), .c(new_n188), .d(new_n200), .o1(new_n207));
  xorc02aa1n12x5               g112(.a(\a[20] ), .b(\b[19] ), .out0(new_n208));
  nor002aa1d32x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  norp02aa1n02x5               g114(.a(new_n208), .b(new_n209), .o1(new_n210));
  inv000aa1d42x5               g115(.a(new_n209), .o1(new_n211));
  inv000aa1d42x5               g116(.a(new_n204), .o1(new_n212));
  aoai13aa1n02x5               g117(.a(new_n211), .b(new_n212), .c(new_n201), .d(new_n203), .o1(new_n213));
  aoi022aa1n03x5               g118(.a(new_n213), .b(new_n208), .c(new_n207), .d(new_n210), .o1(\s[20] ));
  nano32aa1n02x4               g119(.a(new_n212), .b(new_n208), .c(new_n189), .d(new_n197), .out0(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n216));
  nand23aa1d12x5               g121(.a(new_n202), .b(new_n204), .c(new_n208), .o1(new_n217));
  oao003aa1n06x5               g122(.a(\a[20] ), .b(\b[19] ), .c(new_n211), .carry(new_n218));
  nand02aa1d16x5               g123(.a(new_n217), .b(new_n218), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n219), .o1(new_n220));
  xorc02aa1n12x5               g125(.a(\a[21] ), .b(\b[20] ), .out0(new_n221));
  xnbna2aa1n03x5               g126(.a(new_n221), .b(new_n216), .c(new_n220), .out0(\s[21] ));
  aoai13aa1n03x5               g127(.a(new_n221), .b(new_n219), .c(new_n188), .d(new_n215), .o1(new_n223));
  xorc02aa1n12x5               g128(.a(\a[22] ), .b(\b[21] ), .out0(new_n224));
  nor042aa1d18x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  norp02aa1n02x5               g130(.a(new_n224), .b(new_n225), .o1(new_n226));
  inv030aa1n02x5               g131(.a(new_n225), .o1(new_n227));
  xnrc02aa1n02x5               g132(.a(\b[20] ), .b(\a[21] ), .out0(new_n228));
  aoai13aa1n02x5               g133(.a(new_n227), .b(new_n228), .c(new_n216), .d(new_n220), .o1(new_n229));
  aoi022aa1n03x5               g134(.a(new_n229), .b(new_n224), .c(new_n223), .d(new_n226), .o1(\s[22] ));
  nand02aa1n04x5               g135(.a(new_n224), .b(new_n221), .o1(new_n231));
  nano32aa1n02x4               g136(.a(new_n231), .b(new_n200), .c(new_n204), .d(new_n208), .out0(new_n232));
  aoai13aa1n03x5               g137(.a(new_n232), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n231), .o1(new_n234));
  tech160nm_fioaoi03aa1n03p5x5 g139(.a(\a[22] ), .b(\b[21] ), .c(new_n227), .o1(new_n235));
  aoi012aa1n02x5               g140(.a(new_n235), .b(new_n219), .c(new_n234), .o1(new_n236));
  inv040aa1n02x5               g141(.a(new_n236), .o1(new_n237));
  xorc02aa1n12x5               g142(.a(\a[23] ), .b(\b[22] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n237), .c(new_n188), .d(new_n232), .o1(new_n239));
  aoi112aa1n02x5               g144(.a(new_n238), .b(new_n235), .c(new_n219), .d(new_n234), .o1(new_n240));
  aobi12aa1n03x7               g145(.a(new_n239), .b(new_n240), .c(new_n233), .out0(\s[23] ));
  xorc02aa1n12x5               g146(.a(\a[24] ), .b(\b[23] ), .out0(new_n242));
  nor002aa1d32x5               g147(.a(\b[22] ), .b(\a[23] ), .o1(new_n243));
  norp02aa1n02x5               g148(.a(new_n242), .b(new_n243), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n243), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n238), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n246), .c(new_n233), .d(new_n236), .o1(new_n247));
  aoi022aa1n03x5               g152(.a(new_n247), .b(new_n242), .c(new_n239), .d(new_n244), .o1(\s[24] ));
  xnrc02aa1n02x5               g153(.a(\b[21] ), .b(\a[22] ), .out0(new_n249));
  nona23aa1n09x5               g154(.a(new_n238), .b(new_n242), .c(new_n249), .d(new_n228), .out0(new_n250));
  nano32aa1n02x5               g155(.a(new_n250), .b(new_n200), .c(new_n204), .d(new_n208), .out0(new_n251));
  aoai13aa1n03x5               g156(.a(new_n251), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n252));
  oaoi03aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .c(new_n245), .o1(new_n253));
  aoi013aa1n06x4               g158(.a(new_n253), .b(new_n235), .c(new_n238), .d(new_n242), .o1(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n250), .c(new_n217), .d(new_n218), .o1(new_n255));
  xorc02aa1n12x5               g160(.a(\a[25] ), .b(\b[24] ), .out0(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n255), .c(new_n188), .d(new_n251), .o1(new_n257));
  nano22aa1n12x5               g162(.a(new_n231), .b(new_n238), .c(new_n242), .out0(new_n258));
  nand22aa1n12x5               g163(.a(new_n219), .b(new_n258), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n256), .o1(new_n260));
  and003aa1n02x5               g165(.a(new_n259), .b(new_n260), .c(new_n254), .o(new_n261));
  aobi12aa1n03x7               g166(.a(new_n257), .b(new_n261), .c(new_n252), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g167(.a(\a[26] ), .b(\b[25] ), .out0(new_n263));
  nor042aa1n03x5               g168(.a(\b[24] ), .b(\a[25] ), .o1(new_n264));
  norp02aa1n02x5               g169(.a(new_n263), .b(new_n264), .o1(new_n265));
  inv000aa1n02x5               g170(.a(new_n255), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n264), .o1(new_n267));
  aoai13aa1n03x5               g172(.a(new_n267), .b(new_n260), .c(new_n252), .d(new_n266), .o1(new_n268));
  aoi022aa1n03x5               g173(.a(new_n268), .b(new_n263), .c(new_n257), .d(new_n265), .o1(\s[26] ));
  nanp03aa1n02x5               g174(.a(new_n200), .b(new_n204), .c(new_n208), .o1(new_n270));
  and002aa1n12x5               g175(.a(new_n263), .b(new_n256), .o(new_n271));
  inv000aa1n04x5               g176(.a(new_n271), .o1(new_n272));
  nor043aa1n04x5               g177(.a(new_n270), .b(new_n250), .c(new_n272), .o1(new_n273));
  aoai13aa1n06x5               g178(.a(new_n273), .b(new_n195), .c(new_n125), .d(new_n180), .o1(new_n274));
  oao003aa1n02x5               g179(.a(\a[26] ), .b(\b[25] ), .c(new_n267), .carry(new_n275));
  aoai13aa1n12x5               g180(.a(new_n275), .b(new_n272), .c(new_n259), .d(new_n254), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[27] ), .b(\b[26] ), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n276), .c(new_n188), .d(new_n273), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n277), .o1(new_n279));
  nanp02aa1n02x5               g184(.a(new_n275), .b(new_n279), .o1(new_n280));
  aoi012aa1n02x5               g185(.a(new_n280), .b(new_n255), .c(new_n271), .o1(new_n281));
  aobi12aa1n03x7               g186(.a(new_n278), .b(new_n281), .c(new_n274), .out0(\s[27] ));
  xorc02aa1n02x5               g187(.a(\a[28] ), .b(\b[27] ), .out0(new_n283));
  nor042aa1n03x5               g188(.a(\b[26] ), .b(\a[27] ), .o1(new_n284));
  norp02aa1n02x5               g189(.a(new_n283), .b(new_n284), .o1(new_n285));
  aobi12aa1n06x5               g190(.a(new_n275), .b(new_n255), .c(new_n271), .out0(new_n286));
  inv000aa1n03x5               g191(.a(new_n284), .o1(new_n287));
  aoai13aa1n02x7               g192(.a(new_n287), .b(new_n279), .c(new_n274), .d(new_n286), .o1(new_n288));
  aoi022aa1n03x5               g193(.a(new_n288), .b(new_n283), .c(new_n278), .d(new_n285), .o1(\s[28] ));
  and002aa1n02x5               g194(.a(new_n283), .b(new_n277), .o(new_n290));
  aoai13aa1n06x5               g195(.a(new_n290), .b(new_n276), .c(new_n188), .d(new_n273), .o1(new_n291));
  inv000aa1d42x5               g196(.a(new_n290), .o1(new_n292));
  oaoi03aa1n09x5               g197(.a(\a[28] ), .b(\b[27] ), .c(new_n287), .o1(new_n293));
  inv000aa1d42x5               g198(.a(new_n293), .o1(new_n294));
  aoai13aa1n02x7               g199(.a(new_n294), .b(new_n292), .c(new_n274), .d(new_n286), .o1(new_n295));
  xorc02aa1n02x5               g200(.a(\a[29] ), .b(\b[28] ), .out0(new_n296));
  norp02aa1n02x5               g201(.a(new_n293), .b(new_n296), .o1(new_n297));
  aoi022aa1n03x5               g202(.a(new_n295), .b(new_n296), .c(new_n291), .d(new_n297), .o1(\s[29] ));
  xorb03aa1n02x5               g203(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g204(.a(new_n279), .b(new_n283), .c(new_n296), .out0(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n276), .c(new_n188), .d(new_n273), .o1(new_n301));
  inv000aa1d42x5               g206(.a(new_n300), .o1(new_n302));
  inv000aa1d42x5               g207(.a(\a[29] ), .o1(new_n303));
  inv000aa1d42x5               g208(.a(\b[28] ), .o1(new_n304));
  tech160nm_fioaoi03aa1n03p5x5 g209(.a(new_n303), .b(new_n304), .c(new_n293), .o1(new_n305));
  aoai13aa1n02x7               g210(.a(new_n305), .b(new_n302), .c(new_n274), .d(new_n286), .o1(new_n306));
  xorc02aa1n02x5               g211(.a(\a[30] ), .b(\b[29] ), .out0(new_n307));
  oabi12aa1n02x5               g212(.a(new_n307), .b(\a[29] ), .c(\b[28] ), .out0(new_n308));
  oaoi13aa1n02x5               g213(.a(new_n308), .b(new_n293), .c(new_n303), .d(new_n304), .o1(new_n309));
  aoi022aa1n03x5               g214(.a(new_n306), .b(new_n307), .c(new_n301), .d(new_n309), .o1(\s[30] ));
  nano32aa1n09x5               g215(.a(new_n279), .b(new_n307), .c(new_n283), .d(new_n296), .out0(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n276), .c(new_n188), .d(new_n273), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[31] ), .b(\b[30] ), .out0(new_n313));
  oao003aa1n02x5               g218(.a(\a[30] ), .b(\b[29] ), .c(new_n305), .carry(new_n314));
  norb02aa1n02x5               g219(.a(new_n314), .b(new_n313), .out0(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  aoai13aa1n02x7               g221(.a(new_n314), .b(new_n316), .c(new_n274), .d(new_n286), .o1(new_n317));
  aoi022aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n312), .d(new_n315), .o1(\s[31] ));
  inv000aa1d42x5               g223(.a(\b[1] ), .o1(new_n319));
  inv000aa1d42x5               g224(.a(\a[2] ), .o1(new_n320));
  aoi022aa1n02x5               g225(.a(new_n319), .b(new_n320), .c(\a[1] ), .d(\b[0] ), .o1(new_n321));
  oaib12aa1n02x5               g226(.a(new_n321), .b(new_n319), .c(\a[2] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n105), .b(new_n104), .out0(new_n323));
  aboi22aa1n03x5               g228(.a(new_n104), .b(new_n105), .c(new_n320), .d(new_n319), .out0(new_n324));
  aoi022aa1n02x5               g229(.a(new_n322), .b(new_n324), .c(new_n101), .d(new_n323), .o1(\s[3] ));
  obai22aa1n02x7               g230(.a(new_n103), .b(new_n102), .c(\a[3] ), .d(\b[2] ), .out0(new_n326));
  aoi012aa1n02x5               g231(.a(new_n326), .b(new_n101), .c(new_n323), .o1(new_n327));
  oab012aa1n02x4               g232(.a(new_n327), .b(new_n108), .c(new_n102), .out0(\s[4] ));
  norb02aa1n02x5               g233(.a(new_n112), .b(new_n111), .out0(new_n329));
  aoai13aa1n03x5               g234(.a(new_n329), .b(new_n107), .c(new_n106), .d(new_n101), .o1(new_n330));
  aoi112aa1n02x5               g235(.a(new_n107), .b(new_n329), .c(new_n106), .d(new_n101), .o1(new_n331));
  norb02aa1n02x5               g236(.a(new_n330), .b(new_n331), .out0(\s[5] ));
  inv000aa1d42x5               g237(.a(new_n115), .o1(new_n333));
  obai22aa1n02x7               g238(.a(new_n330), .b(new_n111), .c(new_n333), .d(new_n114), .out0(new_n334));
  nona32aa1n03x5               g239(.a(new_n330), .b(new_n333), .c(new_n114), .d(new_n111), .out0(new_n335));
  nanp02aa1n02x5               g240(.a(new_n334), .b(new_n335), .o1(\s[6] ));
  nona23aa1n03x5               g241(.a(new_n335), .b(new_n110), .c(new_n109), .d(new_n333), .out0(new_n337));
  aoi022aa1n02x5               g242(.a(new_n335), .b(new_n115), .c(new_n121), .d(new_n110), .o1(new_n338));
  norb02aa1n02x5               g243(.a(new_n337), .b(new_n338), .out0(\s[7] ));
  xnbna2aa1n03x5               g244(.a(new_n117), .b(new_n337), .c(new_n121), .out0(\s[8] ));
  xnbna2aa1n03x5               g245(.a(new_n127), .b(new_n144), .c(new_n124), .out0(\s[9] ));
endmodule


