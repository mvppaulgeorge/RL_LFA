// Benchmark "adder" written by ABC on Thu Jul 11 12:13:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n204, new_n205, new_n206, new_n207, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n349, new_n352, new_n354, new_n356;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  and002aa1n02x5               g001(.a(\b[8] ), .b(\a[9] ), .o(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  160nm_ficinv00aa1n08x5       g003(.clk(new_n98), .clkout(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  nanp02aa1n02x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  norp02aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  oai012aa1n02x5               g007(.a(new_n100), .b(new_n102), .c(new_n101), .o1(new_n103));
  160nm_ficinv00aa1n08x5       g008(.clk(\a[4] ), .clkout(new_n104));
  160nm_ficinv00aa1n08x5       g009(.clk(\b[3] ), .clkout(new_n105));
  nanp02aa1n02x5               g010(.a(new_n105), .b(new_n104), .o1(new_n106));
  nanp02aa1n02x5               g011(.a(\b[3] ), .b(\a[4] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(new_n106), .b(new_n107), .o1(new_n108));
  160nm_ficinv00aa1n08x5       g013(.clk(\a[3] ), .clkout(new_n109));
  160nm_ficinv00aa1n08x5       g014(.clk(\b[2] ), .clkout(new_n110));
  nanp02aa1n02x5               g015(.a(new_n110), .b(new_n109), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(new_n111), .b(new_n112), .o1(new_n113));
  norp03aa1n02x5               g018(.a(new_n103), .b(new_n108), .c(new_n113), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[2] ), .b(\a[3] ), .o1(new_n115));
  oaoi03aa1n02x5               g020(.a(new_n104), .b(new_n105), .c(new_n115), .o1(new_n116));
  160nm_ficinv00aa1n08x5       g021(.clk(new_n116), .clkout(new_n117));
  norp02aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[7] ), .b(\a[8] ), .o1(new_n119));
  norp02aa1n02x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nanp02aa1n02x5               g025(.a(\b[6] ), .b(\a[7] ), .o1(new_n121));
  nona23aa1n02x4               g026(.a(new_n121), .b(new_n119), .c(new_n118), .d(new_n120), .out0(new_n122));
  xnrc02aa1n02x5               g027(.a(\b[5] ), .b(\a[6] ), .out0(new_n123));
  norp02aa1n02x5               g028(.a(\b[4] ), .b(\a[5] ), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(\b[4] ), .b(\a[5] ), .o1(new_n125));
  nanb02aa1n02x5               g030(.a(new_n124), .b(new_n125), .out0(new_n126));
  norp03aa1n02x5               g031(.a(new_n122), .b(new_n123), .c(new_n126), .o1(new_n127));
  oai012aa1n02x5               g032(.a(new_n127), .b(new_n114), .c(new_n117), .o1(new_n128));
  nano23aa1n02x4               g033(.a(new_n118), .b(new_n120), .c(new_n121), .d(new_n119), .out0(new_n129));
  160nm_ficinv00aa1n08x5       g034(.clk(\a[6] ), .clkout(new_n130));
  160nm_ficinv00aa1n08x5       g035(.clk(\b[5] ), .clkout(new_n131));
  oao003aa1n02x5               g036(.a(new_n130), .b(new_n131), .c(new_n124), .carry(new_n132));
  oa0012aa1n02x5               g037(.a(new_n119), .b(new_n120), .c(new_n118), .o(new_n133));
  aoi012aa1n02x5               g038(.a(new_n133), .b(new_n129), .c(new_n132), .o1(new_n134));
  aoi013aa1n02x4               g039(.a(new_n97), .b(new_n128), .c(new_n134), .d(new_n99), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nanp02aa1n02x5               g041(.a(\b[9] ), .b(\a[10] ), .o1(new_n137));
  norp02aa1n02x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nanp02aa1n02x5               g043(.a(\b[10] ), .b(\a[11] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  norp02aa1n02x5               g045(.a(\b[9] ), .b(\a[10] ), .o1(new_n141));
  160nm_ficinv00aa1n08x5       g046(.clk(new_n141), .clkout(new_n142));
  oai013aa1n02x4               g047(.a(new_n116), .b(new_n108), .c(new_n103), .d(new_n113), .o1(new_n143));
  oaoi03aa1n02x5               g048(.a(new_n130), .b(new_n131), .c(new_n124), .o1(new_n144));
  oabi12aa1n02x5               g049(.a(new_n133), .b(new_n122), .c(new_n144), .out0(new_n145));
  aoi112aa1n02x5               g050(.a(new_n145), .b(new_n98), .c(new_n143), .d(new_n127), .o1(new_n146));
  oai012aa1n02x5               g051(.a(new_n142), .b(new_n146), .c(new_n97), .o1(new_n147));
  xobna2aa1n03x5               g052(.a(new_n140), .b(new_n147), .c(new_n137), .out0(\s[11] ));
  norp02aa1n02x5               g053(.a(\b[11] ), .b(\a[12] ), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(\b[11] ), .b(\a[12] ), .o1(new_n150));
  norb02aa1n02x5               g055(.a(new_n150), .b(new_n149), .out0(new_n151));
  aoi113aa1n02x5               g056(.a(new_n138), .b(new_n151), .c(new_n147), .d(new_n139), .e(new_n137), .o1(new_n152));
  160nm_ficinv00aa1n08x5       g057(.clk(new_n138), .clkout(new_n153));
  nanp03aa1n02x5               g058(.a(new_n147), .b(new_n137), .c(new_n140), .o1(new_n154));
  aobi12aa1n02x5               g059(.a(new_n151), .b(new_n154), .c(new_n153), .out0(new_n155));
  norp02aa1n02x5               g060(.a(new_n155), .b(new_n152), .o1(\s[12] ));
  norb02aa1n02x5               g061(.a(new_n137), .b(new_n141), .out0(new_n157));
  norp02aa1n02x5               g062(.a(new_n97), .b(new_n98), .o1(new_n158));
  nona23aa1n02x4               g063(.a(new_n150), .b(new_n139), .c(new_n138), .d(new_n149), .out0(new_n159));
  nano22aa1n02x4               g064(.a(new_n159), .b(new_n158), .c(new_n157), .out0(new_n160));
  160nm_ficinv00aa1n08x5       g065(.clk(new_n160), .clkout(new_n161));
  nano23aa1n02x4               g066(.a(new_n138), .b(new_n149), .c(new_n150), .d(new_n139), .out0(new_n162));
  aoi012aa1n02x5               g067(.a(new_n141), .b(new_n98), .c(new_n137), .o1(new_n163));
  160nm_ficinv00aa1n08x5       g068(.clk(new_n163), .clkout(new_n164));
  oai012aa1n02x5               g069(.a(new_n150), .b(new_n149), .c(new_n138), .o1(new_n165));
  aobi12aa1n02x5               g070(.a(new_n165), .b(new_n162), .c(new_n164), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n161), .c(new_n128), .d(new_n134), .o1(new_n167));
  xorb03aa1n02x5               g072(.a(new_n167), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n02x5               g073(.a(\b[12] ), .b(\a[13] ), .o1(new_n169));
  nanp02aa1n02x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  aoi012aa1n02x5               g075(.a(new_n169), .b(new_n167), .c(new_n170), .o1(new_n171));
  xnrb03aa1n02x5               g076(.a(new_n171), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  aoai13aa1n02x5               g077(.a(new_n160), .b(new_n145), .c(new_n143), .d(new_n127), .o1(new_n173));
  norp02aa1n02x5               g078(.a(\b[13] ), .b(\a[14] ), .o1(new_n174));
  nanp02aa1n02x5               g079(.a(\b[13] ), .b(\a[14] ), .o1(new_n175));
  nona23aa1n02x4               g080(.a(new_n175), .b(new_n170), .c(new_n169), .d(new_n174), .out0(new_n176));
  aoi012aa1n02x5               g081(.a(new_n174), .b(new_n169), .c(new_n175), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n177), .b(new_n176), .c(new_n173), .d(new_n166), .o1(new_n178));
  xorb03aa1n02x5               g083(.a(new_n178), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g084(.a(\b[14] ), .b(\a[15] ), .o1(new_n180));
  nanp02aa1n02x5               g085(.a(\b[14] ), .b(\a[15] ), .o1(new_n181));
  nanb02aa1n02x5               g086(.a(new_n180), .b(new_n181), .out0(new_n182));
  160nm_ficinv00aa1n08x5       g087(.clk(new_n182), .clkout(new_n183));
  norp02aa1n02x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  nanb02aa1n02x5               g090(.a(new_n184), .b(new_n185), .out0(new_n186));
  160nm_ficinv00aa1n08x5       g091(.clk(new_n186), .clkout(new_n187));
  aoi112aa1n02x5               g092(.a(new_n187), .b(new_n180), .c(new_n178), .d(new_n183), .o1(new_n188));
  160nm_ficinv00aa1n08x5       g093(.clk(new_n180), .clkout(new_n189));
  nano23aa1n02x4               g094(.a(new_n169), .b(new_n174), .c(new_n175), .d(new_n170), .out0(new_n190));
  160nm_ficinv00aa1n08x5       g095(.clk(new_n177), .clkout(new_n191));
  aoai13aa1n02x5               g096(.a(new_n183), .b(new_n191), .c(new_n167), .d(new_n190), .o1(new_n192));
  aoi012aa1n02x5               g097(.a(new_n186), .b(new_n192), .c(new_n189), .o1(new_n193));
  norp02aa1n02x5               g098(.a(new_n193), .b(new_n188), .o1(\s[16] ));
  nona23aa1n02x4               g099(.a(new_n185), .b(new_n181), .c(new_n180), .d(new_n184), .out0(new_n195));
  norp02aa1n02x5               g100(.a(new_n195), .b(new_n176), .o1(new_n196));
  nanp02aa1n02x5               g101(.a(new_n160), .b(new_n196), .o1(new_n197));
  oai012aa1n02x5               g102(.a(new_n165), .b(new_n159), .c(new_n163), .o1(new_n198));
  oai012aa1n02x5               g103(.a(new_n185), .b(new_n184), .c(new_n180), .o1(new_n199));
  oai012aa1n02x5               g104(.a(new_n199), .b(new_n195), .c(new_n177), .o1(new_n200));
  aoi012aa1n02x5               g105(.a(new_n200), .b(new_n198), .c(new_n196), .o1(new_n201));
  aoai13aa1n02x5               g106(.a(new_n201), .b(new_n197), .c(new_n128), .d(new_n134), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g108(.clk(\a[18] ), .clkout(new_n204));
  160nm_ficinv00aa1n08x5       g109(.clk(\a[17] ), .clkout(new_n205));
  160nm_ficinv00aa1n08x5       g110(.clk(\b[16] ), .clkout(new_n206));
  oaoi03aa1n02x5               g111(.a(new_n205), .b(new_n206), .c(new_n202), .o1(new_n207));
  xorb03aa1n02x5               g112(.a(new_n207), .b(\b[17] ), .c(new_n204), .out0(\s[18] ));
  nona22aa1n02x4               g113(.a(new_n190), .b(new_n186), .c(new_n182), .out0(new_n209));
  nano32aa1n02x4               g114(.a(new_n209), .b(new_n162), .c(new_n158), .d(new_n157), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n145), .c(new_n143), .d(new_n127), .o1(new_n211));
  xroi22aa1d04x5               g116(.a(new_n205), .b(\b[16] ), .c(new_n204), .d(\b[17] ), .out0(new_n212));
  160nm_ficinv00aa1n08x5       g117(.clk(new_n212), .clkout(new_n213));
  norp02aa1n02x5               g118(.a(\b[17] ), .b(\a[18] ), .o1(new_n214));
  aoi112aa1n02x5               g119(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n215));
  norp02aa1n02x5               g120(.a(new_n215), .b(new_n214), .o1(new_n216));
  aoai13aa1n02x5               g121(.a(new_n216), .b(new_n213), .c(new_n211), .d(new_n201), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g123(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  xorc02aa1n02x5               g125(.a(\a[19] ), .b(\b[18] ), .out0(new_n221));
  xorc02aa1n02x5               g126(.a(\a[20] ), .b(\b[19] ), .out0(new_n222));
  aoi112aa1n02x5               g127(.a(new_n220), .b(new_n222), .c(new_n217), .d(new_n221), .o1(new_n223));
  160nm_ficinv00aa1n08x5       g128(.clk(new_n220), .clkout(new_n224));
  160nm_ficinv00aa1n08x5       g129(.clk(new_n216), .clkout(new_n225));
  aoai13aa1n02x5               g130(.a(new_n221), .b(new_n225), .c(new_n202), .d(new_n212), .o1(new_n226));
  xnrc02aa1n02x5               g131(.a(\b[19] ), .b(\a[20] ), .out0(new_n227));
  aoi012aa1n02x5               g132(.a(new_n227), .b(new_n226), .c(new_n224), .o1(new_n228));
  norp02aa1n02x5               g133(.a(new_n228), .b(new_n223), .o1(\s[20] ));
  xnrc02aa1n02x5               g134(.a(\b[18] ), .b(\a[19] ), .out0(new_n230));
  norp02aa1n02x5               g135(.a(new_n227), .b(new_n230), .o1(new_n231));
  nanp02aa1n02x5               g136(.a(new_n212), .b(new_n231), .o1(new_n232));
  oaoi03aa1n02x5               g137(.a(\a[20] ), .b(\b[19] ), .c(new_n224), .o1(new_n233));
  aoi012aa1n02x5               g138(.a(new_n233), .b(new_n231), .c(new_n225), .o1(new_n234));
  aoai13aa1n02x5               g139(.a(new_n234), .b(new_n232), .c(new_n211), .d(new_n201), .o1(new_n235));
  xorb03aa1n02x5               g140(.a(new_n235), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g141(.a(\b[20] ), .b(\a[21] ), .o1(new_n237));
  nanp02aa1n02x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n238), .b(new_n237), .out0(new_n239));
  norp02aa1n02x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nanp02aa1n02x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  aoi112aa1n02x5               g147(.a(new_n237), .b(new_n242), .c(new_n235), .d(new_n239), .o1(new_n243));
  160nm_ficinv00aa1n08x5       g148(.clk(new_n237), .clkout(new_n244));
  160nm_ficinv00aa1n08x5       g149(.clk(new_n232), .clkout(new_n245));
  160nm_ficinv00aa1n08x5       g150(.clk(new_n234), .clkout(new_n246));
  aoai13aa1n02x5               g151(.a(new_n239), .b(new_n246), .c(new_n202), .d(new_n245), .o1(new_n247));
  160nm_ficinv00aa1n08x5       g152(.clk(new_n242), .clkout(new_n248));
  aoi012aa1n02x5               g153(.a(new_n248), .b(new_n247), .c(new_n244), .o1(new_n249));
  norp02aa1n02x5               g154(.a(new_n249), .b(new_n243), .o1(\s[22] ));
  nano23aa1n02x4               g155(.a(new_n237), .b(new_n240), .c(new_n241), .d(new_n238), .out0(new_n251));
  nanp03aa1n02x5               g156(.a(new_n212), .b(new_n231), .c(new_n251), .o1(new_n252));
  norp03aa1n02x5               g157(.a(new_n216), .b(new_n230), .c(new_n227), .o1(new_n253));
  oaoi03aa1n02x5               g158(.a(\a[22] ), .b(\b[21] ), .c(new_n244), .o1(new_n254));
  oaoi13aa1n02x5               g159(.a(new_n254), .b(new_n251), .c(new_n253), .d(new_n233), .o1(new_n255));
  aoai13aa1n02x5               g160(.a(new_n255), .b(new_n252), .c(new_n211), .d(new_n201), .o1(new_n256));
  xorb03aa1n02x5               g161(.a(new_n256), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g162(.a(\b[22] ), .b(\a[23] ), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n259), .b(new_n258), .out0(new_n260));
  xorc02aa1n02x5               g165(.a(\a[24] ), .b(\b[23] ), .out0(new_n261));
  aoi112aa1n02x5               g166(.a(new_n258), .b(new_n261), .c(new_n256), .d(new_n260), .o1(new_n262));
  160nm_ficinv00aa1n08x5       g167(.clk(new_n258), .clkout(new_n263));
  160nm_ficinv00aa1n08x5       g168(.clk(new_n252), .clkout(new_n264));
  160nm_ficinv00aa1n08x5       g169(.clk(new_n255), .clkout(new_n265));
  aoai13aa1n02x5               g170(.a(new_n260), .b(new_n265), .c(new_n202), .d(new_n264), .o1(new_n266));
  xnrc02aa1n02x5               g171(.a(\b[23] ), .b(\a[24] ), .out0(new_n267));
  aoi012aa1n02x5               g172(.a(new_n267), .b(new_n266), .c(new_n263), .o1(new_n268));
  norp02aa1n02x5               g173(.a(new_n268), .b(new_n262), .o1(\s[24] ));
  nano22aa1n02x4               g174(.a(new_n267), .b(new_n263), .c(new_n259), .out0(new_n270));
  nano22aa1n02x4               g175(.a(new_n232), .b(new_n251), .c(new_n270), .out0(new_n271));
  160nm_ficinv00aa1n08x5       g176(.clk(new_n271), .clkout(new_n272));
  oai112aa1n02x5               g177(.a(new_n221), .b(new_n222), .c(new_n215), .d(new_n214), .o1(new_n273));
  160nm_ficinv00aa1n08x5       g178(.clk(new_n233), .clkout(new_n274));
  nanp03aa1n02x5               g179(.a(new_n251), .b(new_n260), .c(new_n261), .o1(new_n275));
  aoi012aa1n02x5               g180(.a(new_n275), .b(new_n273), .c(new_n274), .o1(new_n276));
  norp02aa1n02x5               g181(.a(\b[23] ), .b(\a[24] ), .o1(new_n277));
  aoi112aa1n02x5               g182(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n278));
  nanp03aa1n02x5               g183(.a(new_n254), .b(new_n260), .c(new_n261), .o1(new_n279));
  nona22aa1n02x4               g184(.a(new_n279), .b(new_n278), .c(new_n277), .out0(new_n280));
  norp02aa1n02x5               g185(.a(new_n276), .b(new_n280), .o1(new_n281));
  aoai13aa1n02x5               g186(.a(new_n281), .b(new_n272), .c(new_n211), .d(new_n201), .o1(new_n282));
  xorb03aa1n02x5               g187(.a(new_n282), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g188(.a(\b[24] ), .b(\a[25] ), .o1(new_n284));
  xorc02aa1n02x5               g189(.a(\a[25] ), .b(\b[24] ), .out0(new_n285));
  xorc02aa1n02x5               g190(.a(\a[26] ), .b(\b[25] ), .out0(new_n286));
  aoi112aa1n02x5               g191(.a(new_n284), .b(new_n286), .c(new_n282), .d(new_n285), .o1(new_n287));
  160nm_ficinv00aa1n08x5       g192(.clk(new_n284), .clkout(new_n288));
  160nm_ficinv00aa1n08x5       g193(.clk(new_n281), .clkout(new_n289));
  aoai13aa1n02x5               g194(.a(new_n285), .b(new_n289), .c(new_n202), .d(new_n271), .o1(new_n290));
  160nm_ficinv00aa1n08x5       g195(.clk(new_n286), .clkout(new_n291));
  aoi012aa1n02x5               g196(.a(new_n291), .b(new_n290), .c(new_n288), .o1(new_n292));
  norp02aa1n02x5               g197(.a(new_n292), .b(new_n287), .o1(\s[26] ));
  xorc02aa1n02x5               g198(.a(\a[4] ), .b(\b[3] ), .out0(new_n294));
  norb02aa1n02x5               g199(.a(new_n112), .b(new_n115), .out0(new_n295));
  nanb03aa1n02x5               g200(.a(new_n103), .b(new_n294), .c(new_n295), .out0(new_n296));
  nona22aa1n02x4               g201(.a(new_n129), .b(new_n123), .c(new_n126), .out0(new_n297));
  aoai13aa1n02x5               g202(.a(new_n134), .b(new_n297), .c(new_n296), .d(new_n116), .o1(new_n298));
  oabi12aa1n02x5               g203(.a(new_n200), .b(new_n166), .c(new_n209), .out0(new_n299));
  and002aa1n02x5               g204(.a(new_n286), .b(new_n285), .o(new_n300));
  nano22aa1n02x4               g205(.a(new_n252), .b(new_n300), .c(new_n270), .out0(new_n301));
  aoai13aa1n02x5               g206(.a(new_n301), .b(new_n299), .c(new_n298), .d(new_n210), .o1(new_n302));
  oaoi03aa1n02x5               g207(.a(\a[26] ), .b(\b[25] ), .c(new_n288), .o1(new_n303));
  oaoi13aa1n02x5               g208(.a(new_n303), .b(new_n300), .c(new_n276), .d(new_n280), .o1(new_n304));
  norp02aa1n02x5               g209(.a(\b[26] ), .b(\a[27] ), .o1(new_n305));
  and002aa1n02x5               g210(.a(\b[26] ), .b(\a[27] ), .o(new_n306));
  norp02aa1n02x5               g211(.a(new_n306), .b(new_n305), .o1(new_n307));
  xnbna2aa1n03x5               g212(.a(new_n307), .b(new_n302), .c(new_n304), .out0(\s[27] ));
  160nm_ficinv00aa1n08x5       g213(.clk(new_n306), .clkout(new_n309));
  xorc02aa1n02x5               g214(.a(\a[28] ), .b(\b[27] ), .out0(new_n310));
  nano32aa1n02x4               g215(.a(new_n267), .b(new_n260), .c(new_n242), .d(new_n239), .out0(new_n311));
  oai012aa1n02x5               g216(.a(new_n311), .b(new_n253), .c(new_n233), .o1(new_n312));
  aoi113aa1n02x5               g217(.a(new_n278), .b(new_n277), .c(new_n254), .d(new_n261), .e(new_n260), .o1(new_n313));
  160nm_ficinv00aa1n08x5       g218(.clk(new_n300), .clkout(new_n314));
  160nm_ficinv00aa1n08x5       g219(.clk(new_n303), .clkout(new_n315));
  aoai13aa1n02x5               g220(.a(new_n315), .b(new_n314), .c(new_n312), .d(new_n313), .o1(new_n316));
  aoi112aa1n02x5               g221(.a(new_n316), .b(new_n305), .c(new_n202), .d(new_n301), .o1(new_n317));
  nano22aa1n02x4               g222(.a(new_n317), .b(new_n309), .c(new_n310), .out0(new_n318));
  160nm_ficinv00aa1n08x5       g223(.clk(new_n305), .clkout(new_n319));
  nanp03aa1n02x5               g224(.a(new_n302), .b(new_n304), .c(new_n319), .o1(new_n320));
  aoi012aa1n02x5               g225(.a(new_n310), .b(new_n320), .c(new_n309), .o1(new_n321));
  norp02aa1n02x5               g226(.a(new_n321), .b(new_n318), .o1(\s[28] ));
  and002aa1n02x5               g227(.a(new_n310), .b(new_n307), .o(new_n323));
  aoai13aa1n02x5               g228(.a(new_n323), .b(new_n316), .c(new_n202), .d(new_n301), .o1(new_n324));
  oao003aa1n02x5               g229(.a(\a[28] ), .b(\b[27] ), .c(new_n319), .carry(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[28] ), .b(\a[29] ), .out0(new_n326));
  aoi012aa1n02x5               g231(.a(new_n326), .b(new_n324), .c(new_n325), .o1(new_n327));
  aobi12aa1n02x5               g232(.a(new_n323), .b(new_n302), .c(new_n304), .out0(new_n328));
  nano22aa1n02x4               g233(.a(new_n328), .b(new_n325), .c(new_n326), .out0(new_n329));
  norp02aa1n02x5               g234(.a(new_n327), .b(new_n329), .o1(\s[29] ));
  xorb03aa1n02x5               g235(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g236(.a(new_n326), .b(new_n310), .c(new_n307), .out0(new_n332));
  aoai13aa1n02x5               g237(.a(new_n332), .b(new_n316), .c(new_n202), .d(new_n301), .o1(new_n333));
  oao003aa1n02x5               g238(.a(\a[29] ), .b(\b[28] ), .c(new_n325), .carry(new_n334));
  xnrc02aa1n02x5               g239(.a(\b[29] ), .b(\a[30] ), .out0(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n333), .c(new_n334), .o1(new_n336));
  aobi12aa1n02x5               g241(.a(new_n332), .b(new_n302), .c(new_n304), .out0(new_n337));
  nano22aa1n02x4               g242(.a(new_n337), .b(new_n334), .c(new_n335), .out0(new_n338));
  norp02aa1n02x5               g243(.a(new_n336), .b(new_n338), .o1(\s[30] ));
  nano23aa1n02x4               g244(.a(new_n335), .b(new_n326), .c(new_n310), .d(new_n307), .out0(new_n340));
  aobi12aa1n02x5               g245(.a(new_n340), .b(new_n302), .c(new_n304), .out0(new_n341));
  oao003aa1n02x5               g246(.a(\a[30] ), .b(\b[29] ), .c(new_n334), .carry(new_n342));
  xnrc02aa1n02x5               g247(.a(\b[30] ), .b(\a[31] ), .out0(new_n343));
  nano22aa1n02x4               g248(.a(new_n341), .b(new_n342), .c(new_n343), .out0(new_n344));
  aoai13aa1n02x5               g249(.a(new_n340), .b(new_n316), .c(new_n202), .d(new_n301), .o1(new_n345));
  aoi012aa1n02x5               g250(.a(new_n343), .b(new_n345), .c(new_n342), .o1(new_n346));
  norp02aa1n02x5               g251(.a(new_n346), .b(new_n344), .o1(\s[31] ));
  xnbna2aa1n03x5               g252(.a(new_n103), .b(new_n112), .c(new_n111), .out0(\s[3] ));
  oaoi03aa1n02x5               g253(.a(\a[3] ), .b(\b[2] ), .c(new_n103), .o1(new_n349));
  xorb03aa1n02x5               g254(.a(new_n349), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g255(.a(new_n143), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oai013aa1n02x4               g256(.a(new_n125), .b(new_n114), .c(new_n117), .d(new_n124), .o1(new_n352));
  xorb03aa1n02x5               g257(.a(new_n352), .b(\b[5] ), .c(new_n130), .out0(\s[6] ));
  oaoi03aa1n02x5               g258(.a(\a[6] ), .b(\b[5] ), .c(new_n352), .o1(new_n354));
  xorb03aa1n02x5               g259(.a(new_n354), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g260(.a(new_n120), .b(new_n354), .c(new_n121), .o1(new_n356));
  xnrb03aa1n02x5               g261(.a(new_n356), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g262(.a(new_n158), .b(new_n128), .c(new_n134), .out0(\s[9] ));
endmodule


