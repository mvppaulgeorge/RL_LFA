// Benchmark "adder" written by ABC on Thu Jul 18 06:27:25 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n321, new_n324, new_n326, new_n327,
    new_n329;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1d18x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv040aa1d32x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nand42aa1n03x5               g004(.a(new_n99), .b(new_n98), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand22aa1n09x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  aob012aa1n06x5               g007(.a(new_n100), .b(new_n101), .c(new_n102), .out0(new_n103));
  norp02aa1n24x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nand22aa1n12x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb02aa1n03x5               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nor002aa1d32x5               g011(.a(\b[2] ), .b(\a[3] ), .o1(new_n107));
  nand42aa1n04x5               g012(.a(\b[2] ), .b(\a[3] ), .o1(new_n108));
  norb02aa1n02x7               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nanp03aa1n04x5               g014(.a(new_n103), .b(new_n106), .c(new_n109), .o1(new_n110));
  aoi012aa1n06x5               g015(.a(new_n104), .b(new_n107), .c(new_n105), .o1(new_n111));
  nor022aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n09x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n16x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  tech160nm_finand02aa1n05x5   g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nano23aa1n02x4               g020(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n116));
  nand42aa1n04x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nor002aa1d24x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanb02aa1n02x5               g023(.a(new_n118), .b(new_n117), .out0(new_n119));
  inv040aa1d32x5               g024(.a(\a[5] ), .o1(new_n120));
  inv040aa1d32x5               g025(.a(\b[4] ), .o1(new_n121));
  nand22aa1n06x5               g026(.a(new_n121), .b(new_n120), .o1(new_n122));
  nand42aa1n02x5               g027(.a(\b[4] ), .b(\a[5] ), .o1(new_n123));
  nand02aa1n02x5               g028(.a(new_n122), .b(new_n123), .o1(new_n124));
  nona22aa1n02x4               g029(.a(new_n116), .b(new_n119), .c(new_n124), .out0(new_n125));
  oaih12aa1n02x5               g030(.a(new_n113), .b(new_n114), .c(new_n112), .o1(new_n126));
  oaoi03aa1n02x5               g031(.a(\a[6] ), .b(\b[5] ), .c(new_n122), .o1(new_n127));
  aobi12aa1n02x5               g032(.a(new_n126), .b(new_n116), .c(new_n127), .out0(new_n128));
  aoai13aa1n06x5               g033(.a(new_n128), .b(new_n125), .c(new_n110), .d(new_n111), .o1(new_n129));
  nanp02aa1n09x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  aoi012aa1n02x5               g035(.a(new_n97), .b(new_n129), .c(new_n130), .o1(new_n131));
  xnrb03aa1n02x5               g036(.a(new_n131), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n12x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  nand22aa1n04x5               g038(.a(\b[9] ), .b(\a[10] ), .o1(new_n134));
  nano23aa1d15x5               g039(.a(new_n97), .b(new_n133), .c(new_n134), .d(new_n130), .out0(new_n135));
  tech160nm_fioai012aa1n05x5   g040(.a(new_n134), .b(new_n133), .c(new_n97), .o1(new_n136));
  aob012aa1n03x5               g041(.a(new_n136), .b(new_n129), .c(new_n135), .out0(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  inv000aa1d42x5               g043(.a(\a[12] ), .o1(new_n139));
  nor022aa1n16x5               g044(.a(\b[10] ), .b(\a[11] ), .o1(new_n140));
  nand22aa1n09x5               g045(.a(\b[10] ), .b(\a[11] ), .o1(new_n141));
  tech160nm_fiaoi012aa1n05x5   g046(.a(new_n140), .b(new_n137), .c(new_n141), .o1(new_n142));
  xorb03aa1n02x5               g047(.a(new_n142), .b(\b[11] ), .c(new_n139), .out0(\s[12] ));
  tech160nm_fioaoi03aa1n02p5x5 g048(.a(new_n98), .b(new_n99), .c(new_n101), .o1(new_n144));
  nona23aa1n02x5               g049(.a(new_n108), .b(new_n105), .c(new_n104), .d(new_n107), .out0(new_n145));
  oaih12aa1n06x5               g050(.a(new_n111), .b(new_n145), .c(new_n144), .o1(new_n146));
  nona23aa1n06x5               g051(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n147));
  nor043aa1n04x5               g052(.a(new_n147), .b(new_n119), .c(new_n124), .o1(new_n148));
  aoai13aa1n02x7               g053(.a(new_n117), .b(new_n118), .c(new_n121), .d(new_n120), .o1(new_n149));
  tech160nm_fioai012aa1n05x5   g054(.a(new_n126), .b(new_n147), .c(new_n149), .o1(new_n150));
  norp02aa1n24x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nand02aa1d06x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  nona23aa1n03x5               g057(.a(new_n152), .b(new_n141), .c(new_n140), .d(new_n151), .out0(new_n153));
  norb02aa1n02x5               g058(.a(new_n135), .b(new_n153), .out0(new_n154));
  aoai13aa1n06x5               g059(.a(new_n154), .b(new_n150), .c(new_n146), .d(new_n148), .o1(new_n155));
  inv000aa1n02x5               g060(.a(new_n136), .o1(new_n156));
  nano23aa1n03x7               g061(.a(new_n140), .b(new_n151), .c(new_n152), .d(new_n141), .out0(new_n157));
  oai012aa1n02x5               g062(.a(new_n152), .b(new_n151), .c(new_n140), .o1(new_n158));
  aobi12aa1n06x5               g063(.a(new_n158), .b(new_n157), .c(new_n156), .out0(new_n159));
  nanp02aa1n03x5               g064(.a(new_n155), .b(new_n159), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  nand42aa1d28x5               g067(.a(\b[12] ), .b(\a[13] ), .o1(new_n163));
  tech160nm_fiaoi012aa1n05x5   g068(.a(new_n162), .b(new_n160), .c(new_n163), .o1(new_n164));
  xnrb03aa1n03x5               g069(.a(new_n164), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1d32x5               g070(.a(\b[13] ), .b(\a[14] ), .o1(new_n166));
  nand42aa1n20x5               g071(.a(\b[13] ), .b(\a[14] ), .o1(new_n167));
  nano23aa1d15x5               g072(.a(new_n162), .b(new_n166), .c(new_n167), .d(new_n163), .out0(new_n168));
  inv000aa1d42x5               g073(.a(new_n168), .o1(new_n169));
  tech160nm_fioai012aa1n05x5   g074(.a(new_n167), .b(new_n166), .c(new_n162), .o1(new_n170));
  aoai13aa1n06x5               g075(.a(new_n170), .b(new_n169), .c(new_n155), .d(new_n159), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .o1(new_n173));
  nanp02aa1n12x5               g078(.a(\b[14] ), .b(\a[15] ), .o1(new_n174));
  norb02aa1n02x5               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  nor042aa1n06x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  nand42aa1n08x5               g081(.a(\b[15] ), .b(\a[16] ), .o1(new_n177));
  nanb02aa1n02x5               g082(.a(new_n176), .b(new_n177), .out0(new_n178));
  aoai13aa1n03x5               g083(.a(new_n178), .b(new_n173), .c(new_n171), .d(new_n175), .o1(new_n179));
  aoi112aa1n03x4               g084(.a(new_n173), .b(new_n178), .c(new_n171), .d(new_n174), .o1(new_n180));
  nanb02aa1n03x5               g085(.a(new_n180), .b(new_n179), .out0(\s[16] ));
  nano23aa1n09x5               g086(.a(new_n173), .b(new_n176), .c(new_n177), .d(new_n174), .out0(new_n182));
  nand22aa1n09x5               g087(.a(new_n182), .b(new_n168), .o1(new_n183));
  nano22aa1d15x5               g088(.a(new_n183), .b(new_n135), .c(new_n157), .out0(new_n184));
  aoai13aa1n12x5               g089(.a(new_n184), .b(new_n150), .c(new_n146), .d(new_n148), .o1(new_n185));
  oai012aa1n02x7               g090(.a(new_n158), .b(new_n153), .c(new_n136), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n170), .o1(new_n187));
  oai012aa1n02x5               g092(.a(new_n177), .b(new_n176), .c(new_n173), .o1(new_n188));
  aob012aa1n02x5               g093(.a(new_n188), .b(new_n182), .c(new_n187), .out0(new_n189));
  aoib12aa1n12x5               g094(.a(new_n189), .b(new_n186), .c(new_n183), .out0(new_n190));
  xorc02aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n185), .c(new_n190), .out0(\s[17] ));
  inv040aa1d32x5               g097(.a(\a[18] ), .o1(new_n193));
  nanp02aa1n06x5               g098(.a(new_n185), .b(new_n190), .o1(new_n194));
  nor002aa1d32x5               g099(.a(\b[16] ), .b(\a[17] ), .o1(new_n195));
  tech160nm_fiaoi012aa1n05x5   g100(.a(new_n195), .b(new_n194), .c(new_n191), .o1(new_n196));
  xorb03aa1n02x5               g101(.a(new_n196), .b(\b[17] ), .c(new_n193), .out0(\s[18] ));
  inv000aa1d42x5               g102(.a(\a[17] ), .o1(new_n198));
  xroi22aa1d06x4               g103(.a(new_n198), .b(\b[16] ), .c(new_n193), .d(\b[17] ), .out0(new_n199));
  inv000aa1d42x5               g104(.a(new_n199), .o1(new_n200));
  nand02aa1d16x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  nor002aa1d32x5               g106(.a(\b[17] ), .b(\a[18] ), .o1(new_n202));
  nor042aa1n06x5               g107(.a(new_n202), .b(new_n195), .o1(new_n203));
  norb02aa1n02x5               g108(.a(new_n201), .b(new_n203), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  aoai13aa1n04x5               g110(.a(new_n205), .b(new_n200), .c(new_n185), .d(new_n190), .o1(new_n206));
  xorb03aa1n02x5               g111(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n09x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand02aa1d20x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nor022aa1n08x5               g115(.a(\b[19] ), .b(\a[20] ), .o1(new_n211));
  nand02aa1d08x5               g116(.a(\b[19] ), .b(\a[20] ), .o1(new_n212));
  nanb02aa1n02x5               g117(.a(new_n211), .b(new_n212), .out0(new_n213));
  aoai13aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n206), .d(new_n210), .o1(new_n214));
  aoi112aa1n03x4               g119(.a(new_n209), .b(new_n213), .c(new_n206), .d(new_n210), .o1(new_n215));
  nanb02aa1n03x5               g120(.a(new_n215), .b(new_n214), .out0(\s[20] ));
  nanb02aa1n02x5               g121(.a(new_n209), .b(new_n210), .out0(new_n217));
  nona22aa1n03x5               g122(.a(new_n199), .b(new_n217), .c(new_n213), .out0(new_n218));
  orn002aa1n03x5               g123(.a(\a[19] ), .b(\b[18] ), .o(new_n219));
  oai112aa1n06x5               g124(.a(new_n219), .b(new_n201), .c(new_n202), .d(new_n195), .o1(new_n220));
  nanb03aa1n09x5               g125(.a(new_n211), .b(new_n212), .c(new_n210), .out0(new_n221));
  oai012aa1n04x7               g126(.a(new_n212), .b(new_n211), .c(new_n209), .o1(new_n222));
  oai012aa1n18x5               g127(.a(new_n222), .b(new_n220), .c(new_n221), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n04x5               g129(.a(new_n224), .b(new_n218), .c(new_n185), .d(new_n190), .o1(new_n225));
  xorb03aa1n02x5               g130(.a(new_n225), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1d18x5               g131(.a(\b[20] ), .b(\a[21] ), .o1(new_n227));
  xorc02aa1n12x5               g132(.a(\a[21] ), .b(\b[20] ), .out0(new_n228));
  xorc02aa1n12x5               g133(.a(\a[22] ), .b(\b[21] ), .out0(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  aoai13aa1n03x5               g135(.a(new_n230), .b(new_n227), .c(new_n225), .d(new_n228), .o1(new_n231));
  aoi112aa1n03x4               g136(.a(new_n227), .b(new_n230), .c(new_n225), .d(new_n228), .o1(new_n232));
  nanb02aa1n03x5               g137(.a(new_n232), .b(new_n231), .out0(\s[22] ));
  inv000aa1d42x5               g138(.a(\a[21] ), .o1(new_n234));
  inv040aa1d28x5               g139(.a(\a[22] ), .o1(new_n235));
  xroi22aa1d06x4               g140(.a(new_n234), .b(\b[20] ), .c(new_n235), .d(\b[21] ), .out0(new_n236));
  nona23aa1n02x4               g141(.a(new_n199), .b(new_n236), .c(new_n213), .d(new_n217), .out0(new_n237));
  oai012aa1n03x5               g142(.a(new_n201), .b(\b[18] ), .c(\a[19] ), .o1(new_n238));
  nano22aa1n02x4               g143(.a(new_n211), .b(new_n210), .c(new_n212), .out0(new_n239));
  nona22aa1n02x4               g144(.a(new_n239), .b(new_n203), .c(new_n238), .out0(new_n240));
  nanp02aa1n09x5               g145(.a(new_n229), .b(new_n228), .o1(new_n241));
  inv040aa1d32x5               g146(.a(\b[21] ), .o1(new_n242));
  oao003aa1n03x5               g147(.a(new_n235), .b(new_n242), .c(new_n227), .carry(new_n243));
  inv000aa1n02x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n04x5               g149(.a(new_n244), .b(new_n241), .c(new_n240), .d(new_n222), .o1(new_n245));
  inv000aa1n02x5               g150(.a(new_n245), .o1(new_n246));
  aoai13aa1n04x5               g151(.a(new_n246), .b(new_n237), .c(new_n185), .d(new_n190), .o1(new_n247));
  xorb03aa1n02x5               g152(.a(new_n247), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor002aa1n02x5               g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  xorc02aa1n02x5               g154(.a(\a[23] ), .b(\b[22] ), .out0(new_n250));
  xorc02aa1n02x5               g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  inv000aa1d42x5               g156(.a(new_n251), .o1(new_n252));
  aoai13aa1n03x5               g157(.a(new_n252), .b(new_n249), .c(new_n247), .d(new_n250), .o1(new_n253));
  aoi112aa1n03x4               g158(.a(new_n249), .b(new_n252), .c(new_n247), .d(new_n250), .o1(new_n254));
  nanb02aa1n03x5               g159(.a(new_n254), .b(new_n253), .out0(\s[24] ));
  inv000aa1d42x5               g160(.a(\a[23] ), .o1(new_n256));
  inv000aa1d42x5               g161(.a(\a[24] ), .o1(new_n257));
  xroi22aa1d06x4               g162(.a(new_n256), .b(\b[22] ), .c(new_n257), .d(\b[23] ), .out0(new_n258));
  nanb03aa1n06x5               g163(.a(new_n218), .b(new_n258), .c(new_n236), .out0(new_n259));
  inv000aa1d42x5               g164(.a(\b[23] ), .o1(new_n260));
  oao003aa1n06x5               g165(.a(new_n257), .b(new_n260), .c(new_n249), .carry(new_n261));
  aoi012aa1n02x7               g166(.a(new_n261), .b(new_n245), .c(new_n258), .o1(new_n262));
  aoai13aa1n04x5               g167(.a(new_n262), .b(new_n259), .c(new_n185), .d(new_n190), .o1(new_n263));
  xorb03aa1n02x5               g168(.a(new_n263), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g169(.a(\b[24] ), .b(\a[25] ), .o1(new_n265));
  tech160nm_fixorc02aa1n05x5   g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  norp02aa1n04x5               g171(.a(\b[25] ), .b(\a[26] ), .o1(new_n267));
  nand42aa1n03x5               g172(.a(\b[25] ), .b(\a[26] ), .o1(new_n268));
  nanb02aa1n06x5               g173(.a(new_n267), .b(new_n268), .out0(new_n269));
  aoai13aa1n03x5               g174(.a(new_n269), .b(new_n265), .c(new_n263), .d(new_n266), .o1(new_n270));
  aoi112aa1n03x4               g175(.a(new_n265), .b(new_n269), .c(new_n263), .d(new_n266), .o1(new_n271));
  nanb02aa1n03x5               g176(.a(new_n271), .b(new_n270), .out0(\s[26] ));
  aobi12aa1n02x5               g177(.a(new_n188), .b(new_n182), .c(new_n187), .out0(new_n273));
  oai012aa1n02x5               g178(.a(new_n273), .b(new_n159), .c(new_n183), .o1(new_n274));
  norb02aa1n06x5               g179(.a(new_n266), .b(new_n269), .out0(new_n275));
  nano32aa1n03x7               g180(.a(new_n218), .b(new_n275), .c(new_n236), .d(new_n258), .out0(new_n276));
  aoai13aa1n06x5               g181(.a(new_n276), .b(new_n274), .c(new_n129), .d(new_n184), .o1(new_n277));
  aoai13aa1n03x5               g182(.a(new_n275), .b(new_n261), .c(new_n245), .d(new_n258), .o1(new_n278));
  oai012aa1n02x5               g183(.a(new_n268), .b(new_n267), .c(new_n265), .o1(new_n279));
  nand43aa1n03x5               g184(.a(new_n277), .b(new_n278), .c(new_n279), .o1(new_n280));
  xorb03aa1n03x5               g185(.a(new_n280), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1n03x5               g186(.a(\b[26] ), .b(\a[27] ), .o1(new_n282));
  xorc02aa1n02x5               g187(.a(\a[27] ), .b(\b[26] ), .out0(new_n283));
  xnrc02aa1n02x5               g188(.a(\b[27] ), .b(\a[28] ), .out0(new_n284));
  aoai13aa1n03x5               g189(.a(new_n284), .b(new_n282), .c(new_n280), .d(new_n283), .o1(new_n285));
  inv000aa1n02x5               g190(.a(new_n261), .o1(new_n286));
  aoai13aa1n04x5               g191(.a(new_n258), .b(new_n243), .c(new_n223), .d(new_n236), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n275), .o1(new_n288));
  aoai13aa1n06x5               g193(.a(new_n279), .b(new_n288), .c(new_n287), .d(new_n286), .o1(new_n289));
  aoai13aa1n03x5               g194(.a(new_n283), .b(new_n289), .c(new_n194), .d(new_n276), .o1(new_n290));
  nona22aa1n02x5               g195(.a(new_n290), .b(new_n284), .c(new_n282), .out0(new_n291));
  nanp02aa1n03x5               g196(.a(new_n285), .b(new_n291), .o1(\s[28] ));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  norb02aa1n02x5               g198(.a(new_n283), .b(new_n284), .out0(new_n294));
  inv000aa1n03x5               g199(.a(new_n282), .o1(new_n295));
  oaoi03aa1n02x5               g200(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .o1(new_n296));
  aoai13aa1n03x5               g201(.a(new_n293), .b(new_n296), .c(new_n280), .d(new_n294), .o1(new_n297));
  aoai13aa1n03x5               g202(.a(new_n294), .b(new_n289), .c(new_n194), .d(new_n276), .o1(new_n298));
  nona22aa1n02x5               g203(.a(new_n298), .b(new_n296), .c(new_n293), .out0(new_n299));
  nanp02aa1n03x5               g204(.a(new_n297), .b(new_n299), .o1(\s[29] ));
  xorb03aa1n02x5               g205(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g206(.a(new_n283), .b(new_n293), .c(new_n284), .out0(new_n302));
  oao003aa1n03x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n295), .carry(new_n303));
  oaoi03aa1n02x5               g208(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .o1(new_n304));
  nor002aa1n02x5               g209(.a(\b[29] ), .b(\a[30] ), .o1(new_n305));
  and002aa1n03x5               g210(.a(\b[29] ), .b(\a[30] ), .o(new_n306));
  nor042aa1n02x5               g211(.a(new_n306), .b(new_n305), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n307), .o1(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n304), .c(new_n280), .d(new_n302), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n302), .b(new_n289), .c(new_n194), .d(new_n276), .o1(new_n310));
  nona32aa1n02x5               g215(.a(new_n310), .b(new_n306), .c(new_n305), .d(new_n304), .out0(new_n311));
  nanp02aa1n03x5               g216(.a(new_n309), .b(new_n311), .o1(\s[30] ));
  nano23aa1n02x4               g217(.a(new_n293), .b(new_n284), .c(new_n283), .d(new_n307), .out0(new_n313));
  tech160nm_fiao0012aa1n02p5x5 g218(.a(new_n305), .b(new_n304), .c(new_n307), .o(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[30] ), .b(\a[31] ), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n314), .c(new_n280), .d(new_n313), .o1(new_n316));
  aoai13aa1n03x5               g221(.a(new_n313), .b(new_n289), .c(new_n194), .d(new_n276), .o1(new_n317));
  nona22aa1n02x5               g222(.a(new_n317), .b(new_n314), .c(new_n315), .out0(new_n318));
  nanp02aa1n03x5               g223(.a(new_n316), .b(new_n318), .o1(\s[31] ));
  xorb03aa1n02x5               g224(.a(new_n103), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  aoi012aa1n02x5               g225(.a(new_n107), .b(new_n103), .c(new_n108), .o1(new_n321));
  xnrc02aa1n02x5               g226(.a(new_n321), .b(new_n106), .out0(\s[4] ));
  xorb03aa1n02x5               g227(.a(new_n146), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoai13aa1n02x5               g228(.a(new_n122), .b(new_n124), .c(new_n110), .d(new_n111), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  orn002aa1n02x5               g230(.a(new_n119), .b(new_n124), .o(new_n326));
  aoai13aa1n02x5               g231(.a(new_n149), .b(new_n326), .c(new_n110), .d(new_n111), .o1(new_n327));
  xorb03aa1n02x5               g232(.a(new_n327), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi012aa1n02x5               g233(.a(new_n114), .b(new_n327), .c(new_n115), .o1(new_n329));
  xnrb03aa1n02x5               g234(.a(new_n329), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g235(.a(new_n129), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


