// Benchmark "adder" written by ABC on Thu Jul 18 05:14:50 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n317,
    new_n318, new_n320, new_n321, new_n322, new_n323, new_n325, new_n326,
    new_n328, new_n329, new_n330;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  tech160nm_fixorc02aa1n03p5x5 g001(.a(\a[10] ), .b(\b[9] ), .out0(new_n97));
  inv000aa1d42x5               g002(.a(\b[8] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(\a[9] ), .b(new_n98), .out0(new_n99));
  and002aa1n12x5               g004(.a(\b[0] ), .b(\a[1] ), .o(new_n100));
  oaoi03aa1n12x5               g005(.a(\a[2] ), .b(\b[1] ), .c(new_n100), .o1(new_n101));
  xorc02aa1n12x5               g006(.a(\a[3] ), .b(\b[2] ), .out0(new_n102));
  oaih22aa1n04x5               g007(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n103));
  aoi012aa1n12x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .o1(new_n104));
  nor042aa1n06x5               g009(.a(\b[6] ), .b(\a[7] ), .o1(new_n105));
  nanp02aa1n04x5               g010(.a(\b[7] ), .b(\a[8] ), .o1(new_n106));
  nand42aa1n08x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nano22aa1n03x7               g012(.a(new_n105), .b(new_n106), .c(new_n107), .out0(new_n108));
  nor002aa1d32x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  and002aa1n03x5               g014(.a(\b[4] ), .b(\a[5] ), .o(new_n110));
  aoi112aa1n06x5               g015(.a(new_n110), .b(new_n109), .c(\a[4] ), .d(\b[3] ), .o1(new_n111));
  nor042aa1n03x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  and002aa1n12x5               g017(.a(\b[5] ), .b(\a[6] ), .o(new_n113));
  nor042aa1n04x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nor043aa1n02x5               g019(.a(new_n113), .b(new_n114), .c(new_n112), .o1(new_n115));
  nand23aa1n04x5               g020(.a(new_n111), .b(new_n108), .c(new_n115), .o1(new_n116));
  norb02aa1n09x5               g021(.a(new_n106), .b(new_n112), .out0(new_n117));
  norb02aa1n02x7               g022(.a(new_n107), .b(new_n105), .out0(new_n118));
  oab012aa1n04x5               g023(.a(new_n113), .b(new_n109), .c(new_n114), .out0(new_n119));
  inv000aa1n02x5               g024(.a(new_n105), .o1(new_n120));
  oaoi03aa1n02x5               g025(.a(\a[8] ), .b(\b[7] ), .c(new_n120), .o1(new_n121));
  aoi013aa1n06x4               g026(.a(new_n121), .b(new_n119), .c(new_n117), .d(new_n118), .o1(new_n122));
  oai012aa1d24x5               g027(.a(new_n122), .b(new_n104), .c(new_n116), .o1(new_n123));
  oaib12aa1n09x5               g028(.a(new_n123), .b(new_n98), .c(\a[9] ), .out0(new_n124));
  xnbna2aa1n03x5               g029(.a(new_n97), .b(new_n124), .c(new_n99), .out0(\s[10] ));
  nanp02aa1n04x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nor042aa1n09x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  nanb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  nanp02aa1n02x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  oai022aa1n03x5               g034(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n130));
  oaib12aa1n02x5               g035(.a(new_n129), .b(new_n130), .c(new_n124), .out0(new_n131));
  nano22aa1n02x4               g036(.a(new_n127), .b(new_n129), .c(new_n126), .out0(new_n132));
  oaib12aa1n03x5               g037(.a(new_n132), .b(new_n130), .c(new_n124), .out0(new_n133));
  aobi12aa1n02x5               g038(.a(new_n133), .b(new_n131), .c(new_n128), .out0(\s[11] ));
  inv000aa1d42x5               g039(.a(new_n127), .o1(new_n135));
  norp02aa1n04x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanp02aa1n04x5               g041(.a(\b[11] ), .b(\a[12] ), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(new_n138));
  norp02aa1n02x5               g043(.a(new_n136), .b(new_n127), .o1(new_n139));
  nanp03aa1n02x5               g044(.a(new_n133), .b(new_n137), .c(new_n139), .o1(new_n140));
  aoai13aa1n02x5               g045(.a(new_n140), .b(new_n138), .c(new_n135), .d(new_n133), .o1(\s[12] ));
  nano23aa1n06x5               g046(.a(new_n136), .b(new_n127), .c(new_n137), .d(new_n126), .out0(new_n142));
  xnrc02aa1n02x5               g047(.a(\b[8] ), .b(\a[9] ), .out0(new_n143));
  nanb03aa1n06x5               g048(.a(new_n143), .b(new_n142), .c(new_n97), .out0(new_n144));
  nanb02aa1n09x5               g049(.a(new_n144), .b(new_n123), .out0(new_n145));
  aoi022aa1n02x5               g050(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n146));
  aoi112aa1n03x5               g051(.a(new_n136), .b(new_n127), .c(new_n130), .d(new_n146), .o1(new_n147));
  nanb02aa1n02x5               g052(.a(new_n147), .b(new_n137), .out0(new_n148));
  nor002aa1d32x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  nand42aa1d28x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nanb02aa1n02x5               g055(.a(new_n149), .b(new_n150), .out0(new_n151));
  xobna2aa1n03x5               g056(.a(new_n151), .b(new_n145), .c(new_n148), .out0(\s[13] ));
  aoi012aa1n02x5               g057(.a(new_n151), .b(new_n145), .c(new_n148), .o1(new_n153));
  nor042aa1n06x5               g058(.a(\b[13] ), .b(\a[14] ), .o1(new_n154));
  nand42aa1d28x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  inv040aa1n08x5               g060(.a(new_n149), .o1(new_n156));
  aoai13aa1n02x5               g061(.a(new_n156), .b(new_n151), .c(new_n145), .d(new_n148), .o1(new_n157));
  oaib12aa1n02x5               g062(.a(new_n157), .b(new_n154), .c(new_n155), .out0(new_n158));
  norb03aa1n02x5               g063(.a(new_n155), .b(new_n149), .c(new_n154), .out0(new_n159));
  oaib12aa1n02x5               g064(.a(new_n158), .b(new_n153), .c(new_n159), .out0(\s[14] ));
  nano23aa1d15x5               g065(.a(new_n149), .b(new_n154), .c(new_n155), .d(new_n150), .out0(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  oaoi03aa1n12x5               g067(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n162), .c(new_n145), .d(new_n148), .o1(new_n165));
  xorb03aa1n02x5               g070(.a(new_n165), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1d32x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nanp02aa1n09x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  tech160nm_fixnrc02aa1n04x5   g073(.a(\b[15] ), .b(\a[16] ), .out0(new_n169));
  aoai13aa1n03x5               g074(.a(new_n169), .b(new_n167), .c(new_n165), .d(new_n168), .o1(new_n170));
  nanb02aa1d24x5               g075(.a(new_n167), .b(new_n168), .out0(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  norp02aa1n02x5               g077(.a(new_n169), .b(new_n167), .o1(new_n173));
  aob012aa1n03x5               g078(.a(new_n173), .b(new_n165), .c(new_n172), .out0(new_n174));
  nanp02aa1n03x5               g079(.a(new_n170), .b(new_n174), .o1(\s[16] ));
  inv040aa1d32x5               g080(.a(\a[17] ), .o1(new_n176));
  nona22aa1n02x4               g081(.a(new_n161), .b(new_n169), .c(new_n171), .out0(new_n177));
  nor042aa1n06x5               g082(.a(new_n144), .b(new_n177), .o1(new_n178));
  nor002aa1n06x5               g083(.a(\b[15] ), .b(\a[16] ), .o1(new_n179));
  aoi012aa1n02x7               g084(.a(new_n179), .b(\a[12] ), .c(\b[11] ), .o1(new_n180));
  nona23aa1d18x5               g085(.a(new_n161), .b(new_n180), .c(new_n169), .d(new_n171), .out0(new_n181));
  aoi022aa1n02x5               g086(.a(\b[15] ), .b(\a[16] ), .c(\a[15] ), .d(\b[14] ), .o1(new_n182));
  oaoi13aa1n12x5               g087(.a(new_n179), .b(new_n182), .c(new_n163), .d(new_n167), .o1(new_n183));
  oai012aa1n18x5               g088(.a(new_n183), .b(new_n181), .c(new_n147), .o1(new_n184));
  aoi012aa1n02x7               g089(.a(new_n184), .b(new_n123), .c(new_n178), .o1(new_n185));
  xorb03aa1n02x5               g090(.a(new_n185), .b(\b[16] ), .c(new_n176), .out0(\s[17] ));
  xnrc02aa1n12x5               g091(.a(\b[17] ), .b(\a[18] ), .out0(new_n187));
  oaoi03aa1n02x5               g092(.a(\a[17] ), .b(\b[16] ), .c(new_n185), .o1(new_n188));
  xnrc02aa1n02x5               g093(.a(\b[16] ), .b(\a[17] ), .out0(new_n189));
  inv040aa1n18x5               g094(.a(\b[16] ), .o1(new_n190));
  nand22aa1n12x5               g095(.a(new_n190), .b(new_n176), .o1(new_n191));
  norb02aa1n02x5               g096(.a(new_n191), .b(new_n187), .out0(new_n192));
  oai012aa1n02x5               g097(.a(new_n192), .b(new_n185), .c(new_n189), .o1(new_n193));
  aob012aa1n03x5               g098(.a(new_n193), .b(new_n188), .c(new_n187), .out0(\s[18] ));
  norp02aa1n02x5               g099(.a(new_n187), .b(new_n189), .o1(new_n195));
  aoai13aa1n06x5               g100(.a(new_n195), .b(new_n184), .c(new_n123), .d(new_n178), .o1(new_n196));
  oaoi03aa1n12x5               g101(.a(\a[18] ), .b(\b[17] ), .c(new_n191), .o1(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  nor002aa1d32x5               g103(.a(\b[18] ), .b(\a[19] ), .o1(new_n199));
  nand42aa1d28x5               g104(.a(\b[18] ), .b(\a[19] ), .o1(new_n200));
  norb02aa1n15x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n196), .c(new_n198), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1n08x5               g108(.a(new_n199), .o1(new_n204));
  aob012aa1n02x5               g109(.a(new_n201), .b(new_n196), .c(new_n198), .out0(new_n205));
  nor042aa1n04x5               g110(.a(\b[19] ), .b(\a[20] ), .o1(new_n206));
  nand42aa1n16x5               g111(.a(\b[19] ), .b(\a[20] ), .o1(new_n207));
  norb02aa1n03x5               g112(.a(new_n207), .b(new_n206), .out0(new_n208));
  inv000aa1d42x5               g113(.a(new_n201), .o1(new_n209));
  norb03aa1n02x5               g114(.a(new_n207), .b(new_n199), .c(new_n206), .out0(new_n210));
  aoai13aa1n02x5               g115(.a(new_n210), .b(new_n209), .c(new_n196), .d(new_n198), .o1(new_n211));
  aoai13aa1n02x5               g116(.a(new_n211), .b(new_n208), .c(new_n205), .d(new_n204), .o1(\s[20] ));
  nano23aa1n06x5               g117(.a(new_n199), .b(new_n206), .c(new_n207), .d(new_n200), .out0(new_n213));
  nona22aa1n09x5               g118(.a(new_n213), .b(new_n187), .c(new_n189), .out0(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  aoai13aa1n06x5               g120(.a(new_n215), .b(new_n184), .c(new_n123), .d(new_n178), .o1(new_n216));
  oaoi03aa1n06x5               g121(.a(\a[20] ), .b(\b[19] ), .c(new_n204), .o1(new_n217));
  aoi012aa1n02x5               g122(.a(new_n217), .b(new_n213), .c(new_n197), .o1(new_n218));
  tech160nm_fixnrc02aa1n05x5   g123(.a(\b[20] ), .b(\a[21] ), .out0(new_n219));
  xobna2aa1n03x5               g124(.a(new_n219), .b(new_n216), .c(new_n218), .out0(\s[21] ));
  aoi012aa1n03x5               g125(.a(new_n219), .b(new_n216), .c(new_n218), .o1(new_n221));
  tech160nm_fixorc02aa1n02p5x5 g126(.a(\a[22] ), .b(\b[21] ), .out0(new_n222));
  norp02aa1n02x5               g127(.a(\b[20] ), .b(\a[21] ), .o1(new_n223));
  nor002aa1n02x5               g128(.a(new_n221), .b(new_n223), .o1(new_n224));
  nanp02aa1n02x5               g129(.a(\b[21] ), .b(\a[22] ), .o1(new_n225));
  oai022aa1n02x5               g130(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n226));
  nanb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  oai022aa1n02x5               g132(.a(new_n224), .b(new_n222), .c(new_n227), .d(new_n221), .o1(\s[22] ));
  nanb02aa1n06x5               g133(.a(new_n219), .b(new_n222), .out0(new_n229));
  norp02aa1n02x5               g134(.a(new_n214), .b(new_n229), .o1(new_n230));
  aoai13aa1n06x5               g135(.a(new_n230), .b(new_n184), .c(new_n123), .d(new_n178), .o1(new_n231));
  nor042aa1n02x5               g136(.a(\b[17] ), .b(\a[18] ), .o1(new_n232));
  aoi112aa1n06x5               g137(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n233));
  oai112aa1n06x5               g138(.a(new_n201), .b(new_n208), .c(new_n233), .d(new_n232), .o1(new_n234));
  inv000aa1n04x5               g139(.a(new_n217), .o1(new_n235));
  nand02aa1d04x5               g140(.a(new_n226), .b(new_n225), .o1(new_n236));
  aoai13aa1n12x5               g141(.a(new_n236), .b(new_n229), .c(new_n234), .d(new_n235), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  xnrc02aa1n12x5               g143(.a(\b[22] ), .b(\a[23] ), .out0(new_n239));
  xobna2aa1n03x5               g144(.a(new_n239), .b(new_n231), .c(new_n238), .out0(\s[23] ));
  nor042aa1n03x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  inv000aa1n03x5               g146(.a(new_n241), .o1(new_n242));
  tech160nm_fiao0012aa1n02p5x5 g147(.a(new_n239), .b(new_n231), .c(new_n238), .o(new_n243));
  xorc02aa1n06x5               g148(.a(\a[24] ), .b(\b[23] ), .out0(new_n244));
  nanp02aa1n02x5               g149(.a(\b[23] ), .b(\a[24] ), .o1(new_n245));
  oai022aa1n02x5               g150(.a(\a[23] ), .b(\b[22] ), .c(\b[23] ), .d(\a[24] ), .o1(new_n246));
  norb02aa1n02x5               g151(.a(new_n245), .b(new_n246), .out0(new_n247));
  aoai13aa1n02x5               g152(.a(new_n247), .b(new_n239), .c(new_n231), .d(new_n238), .o1(new_n248));
  aoai13aa1n02x5               g153(.a(new_n248), .b(new_n244), .c(new_n243), .d(new_n242), .o1(\s[24] ));
  orn002aa1n02x5               g154(.a(\a[22] ), .b(\b[21] ), .o(new_n250));
  nano22aa1n03x7               g155(.a(new_n219), .b(new_n250), .c(new_n225), .out0(new_n251));
  norb02aa1n02x7               g156(.a(new_n244), .b(new_n239), .out0(new_n252));
  inv000aa1n02x5               g157(.a(new_n252), .o1(new_n253));
  nano32aa1n03x7               g158(.a(new_n253), .b(new_n251), .c(new_n195), .d(new_n213), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n184), .c(new_n123), .d(new_n178), .o1(new_n255));
  aoai13aa1n06x5               g160(.a(new_n251), .b(new_n217), .c(new_n213), .d(new_n197), .o1(new_n256));
  oaoi03aa1n02x5               g161(.a(\a[24] ), .b(\b[23] ), .c(new_n242), .o1(new_n257));
  inv000aa1n02x5               g162(.a(new_n257), .o1(new_n258));
  aoai13aa1n12x5               g163(.a(new_n258), .b(new_n253), .c(new_n256), .d(new_n236), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  xorc02aa1n12x5               g165(.a(\a[25] ), .b(\b[24] ), .out0(new_n261));
  xnbna2aa1n03x5               g166(.a(new_n261), .b(new_n255), .c(new_n260), .out0(\s[25] ));
  norp02aa1n02x5               g167(.a(\b[24] ), .b(\a[25] ), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n263), .o1(new_n264));
  aob012aa1n03x5               g169(.a(new_n261), .b(new_n255), .c(new_n260), .out0(new_n265));
  tech160nm_fixorc02aa1n02p5x5 g170(.a(\a[26] ), .b(\b[25] ), .out0(new_n266));
  nanp02aa1n02x5               g171(.a(\b[25] ), .b(\a[26] ), .o1(new_n267));
  oai022aa1n02x5               g172(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n268));
  norb02aa1n02x5               g173(.a(new_n267), .b(new_n268), .out0(new_n269));
  nanp02aa1n03x5               g174(.a(new_n265), .b(new_n269), .o1(new_n270));
  aoai13aa1n02x5               g175(.a(new_n270), .b(new_n266), .c(new_n265), .d(new_n264), .o1(\s[26] ));
  and002aa1n02x5               g176(.a(new_n266), .b(new_n261), .o(new_n272));
  nano32aa1n06x5               g177(.a(new_n214), .b(new_n272), .c(new_n251), .d(new_n252), .out0(new_n273));
  aoai13aa1n12x5               g178(.a(new_n273), .b(new_n184), .c(new_n123), .d(new_n178), .o1(new_n274));
  aoai13aa1n06x5               g179(.a(new_n272), .b(new_n257), .c(new_n237), .d(new_n252), .o1(new_n275));
  nanp02aa1n02x5               g180(.a(new_n268), .b(new_n267), .o1(new_n276));
  nand23aa1n06x5               g181(.a(new_n274), .b(new_n275), .c(new_n276), .o1(new_n277));
  xorb03aa1n02x5               g182(.a(new_n277), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  norp02aa1n02x5               g183(.a(\b[26] ), .b(\a[27] ), .o1(new_n279));
  xorc02aa1n12x5               g184(.a(\a[27] ), .b(\b[26] ), .out0(new_n280));
  xnrc02aa1n12x5               g185(.a(\b[27] ), .b(\a[28] ), .out0(new_n281));
  aoai13aa1n03x5               g186(.a(new_n281), .b(new_n279), .c(new_n277), .d(new_n280), .o1(new_n282));
  aoi022aa1n09x5               g187(.a(new_n259), .b(new_n272), .c(new_n267), .d(new_n268), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n280), .o1(new_n284));
  nor042aa1n03x5               g189(.a(new_n281), .b(new_n279), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n284), .c(new_n283), .d(new_n274), .o1(new_n286));
  nanp02aa1n03x5               g191(.a(new_n282), .b(new_n286), .o1(\s[28] ));
  norb02aa1n15x5               g192(.a(new_n280), .b(new_n281), .out0(new_n288));
  nand02aa1n02x5               g193(.a(new_n277), .b(new_n288), .o1(new_n289));
  inv000aa1d42x5               g194(.a(new_n288), .o1(new_n290));
  ao0012aa1n12x5               g195(.a(new_n285), .b(\a[28] ), .c(\b[27] ), .o(new_n291));
  aoai13aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n283), .d(new_n274), .o1(new_n292));
  xorc02aa1n02x5               g197(.a(\a[29] ), .b(\b[28] ), .out0(new_n293));
  norb02aa1n02x5               g198(.a(new_n291), .b(new_n293), .out0(new_n294));
  aoi022aa1n03x5               g199(.a(new_n292), .b(new_n293), .c(new_n289), .d(new_n294), .o1(\s[29] ));
  xnrb03aa1n02x5               g200(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g201(.a(new_n281), .b(new_n280), .c(new_n293), .out0(new_n297));
  nand02aa1n02x5               g202(.a(new_n277), .b(new_n297), .o1(new_n298));
  inv000aa1n02x5               g203(.a(new_n297), .o1(new_n299));
  oaoi03aa1n12x5               g204(.a(\a[29] ), .b(\b[28] ), .c(new_n291), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n300), .o1(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n299), .c(new_n283), .d(new_n274), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .out0(new_n303));
  norp02aa1n02x5               g208(.a(new_n300), .b(new_n303), .o1(new_n304));
  aoi022aa1n03x5               g209(.a(new_n302), .b(new_n303), .c(new_n298), .d(new_n304), .o1(\s[30] ));
  nanp03aa1n02x5               g210(.a(new_n288), .b(new_n293), .c(new_n303), .o1(new_n306));
  nanb02aa1n03x5               g211(.a(new_n306), .b(new_n277), .out0(new_n307));
  inv000aa1d42x5               g212(.a(\a[30] ), .o1(new_n308));
  inv000aa1d42x5               g213(.a(\b[29] ), .o1(new_n309));
  oaoi03aa1n03x5               g214(.a(new_n308), .b(new_n309), .c(new_n300), .o1(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n306), .c(new_n283), .d(new_n274), .o1(new_n311));
  xorc02aa1n02x5               g216(.a(\a[31] ), .b(\b[30] ), .out0(new_n312));
  norb02aa1n02x7               g217(.a(new_n310), .b(new_n312), .out0(new_n313));
  aoi022aa1n03x5               g218(.a(new_n311), .b(new_n312), .c(new_n307), .d(new_n313), .o1(\s[31] ));
  xorb03aa1n02x5               g219(.a(new_n101), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  nanp02aa1n02x5               g220(.a(new_n101), .b(new_n102), .o1(new_n316));
  xorc02aa1n02x5               g221(.a(\a[4] ), .b(\b[3] ), .out0(new_n317));
  oab012aa1n02x4               g222(.a(new_n317), .b(\a[3] ), .c(\b[2] ), .out0(new_n318));
  aboi22aa1n03x5               g223(.a(new_n104), .b(new_n317), .c(new_n318), .d(new_n316), .out0(\s[4] ));
  and002aa1n02x5               g224(.a(\b[3] ), .b(\a[4] ), .o(new_n320));
  aoai13aa1n12x5               g225(.a(new_n111), .b(new_n103), .c(new_n101), .d(new_n102), .o1(new_n321));
  inv000aa1d42x5               g226(.a(new_n321), .o1(new_n322));
  xnrc02aa1n02x5               g227(.a(\b[4] ), .b(\a[5] ), .out0(new_n323));
  oaoi13aa1n02x5               g228(.a(new_n322), .b(new_n323), .c(new_n104), .d(new_n320), .o1(\s[5] ));
  inv000aa1d42x5               g229(.a(new_n109), .o1(new_n325));
  xnrc02aa1n02x5               g230(.a(\b[5] ), .b(\a[6] ), .out0(new_n326));
  xobna2aa1n03x5               g231(.a(new_n326), .b(new_n321), .c(new_n325), .out0(\s[6] ));
  nona32aa1n06x5               g232(.a(new_n321), .b(new_n114), .c(new_n113), .d(new_n109), .out0(new_n328));
  aboi22aa1n03x5               g233(.a(new_n113), .b(new_n328), .c(new_n120), .d(new_n107), .out0(new_n329));
  nona23aa1n06x5               g234(.a(new_n328), .b(new_n107), .c(new_n105), .d(new_n113), .out0(new_n330));
  norb02aa1n02x5               g235(.a(new_n330), .b(new_n329), .out0(\s[7] ));
  xnbna2aa1n03x5               g236(.a(new_n117), .b(new_n330), .c(new_n120), .out0(\s[8] ));
  xorb03aa1n02x5               g237(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


