// Benchmark "adder" written by ABC on Wed Jul 17 23:27:36 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n267, new_n268, new_n269, new_n270, new_n271, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n344,
    new_n345, new_n347, new_n348, new_n349, new_n351, new_n352, new_n353,
    new_n355, new_n356, new_n358, new_n359, new_n361, new_n362;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nanp02aa1n04x5               g001(.a(\b[2] ), .b(\a[3] ), .o1(new_n97));
  nor042aa1d18x5               g002(.a(\b[2] ), .b(\a[3] ), .o1(new_n98));
  nand42aa1d28x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nano22aa1n03x7               g004(.a(new_n98), .b(new_n97), .c(new_n99), .out0(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nor002aa1n06x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nona22aa1n09x5               g007(.a(new_n99), .b(new_n102), .c(new_n101), .out0(new_n103));
  oai022aa1d24x5               g008(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n104));
  aoi012aa1n06x5               g009(.a(new_n104), .b(new_n100), .c(new_n103), .o1(new_n105));
  inv000aa1d42x5               g010(.a(\a[5] ), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\b[4] ), .o1(new_n107));
  nanp02aa1n09x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nand42aa1n10x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  oai112aa1n06x5               g014(.a(new_n108), .b(new_n109), .c(new_n107), .d(new_n106), .o1(new_n110));
  xorc02aa1n12x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  oai022aa1d24x5               g016(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n112));
  nand02aa1d08x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  tech160nm_fioai012aa1n03p5x5 g018(.a(new_n113), .b(\b[6] ), .c(\a[7] ), .o1(new_n114));
  nor042aa1n02x5               g019(.a(new_n114), .b(new_n112), .o1(new_n115));
  nanb03aa1n12x5               g020(.a(new_n110), .b(new_n115), .c(new_n111), .out0(new_n116));
  nor042aa1d18x5               g021(.a(\b[6] ), .b(\a[7] ), .o1(new_n117));
  nano22aa1n03x7               g022(.a(new_n117), .b(new_n108), .c(new_n113), .out0(new_n118));
  inv000aa1d42x5               g023(.a(\a[8] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[7] ), .o1(new_n120));
  tech160nm_fioaoi03aa1n02p5x5 g025(.a(new_n119), .b(new_n120), .c(new_n117), .o1(new_n121));
  inv030aa1n02x5               g026(.a(new_n121), .o1(new_n122));
  aoi013aa1n09x5               g027(.a(new_n122), .b(new_n118), .c(new_n111), .d(new_n112), .o1(new_n123));
  oai012aa1n18x5               g028(.a(new_n123), .b(new_n105), .c(new_n116), .o1(new_n124));
  nor002aa1d24x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nand02aa1d08x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n06x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  nor002aa1d32x5               g032(.a(\b[9] ), .b(\a[10] ), .o1(new_n128));
  nanp02aa1n04x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nanb02aa1n02x5               g034(.a(new_n128), .b(new_n129), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n130), .b(new_n125), .c(new_n124), .d(new_n126), .o1(new_n131));
  nona22aa1n02x4               g036(.a(new_n129), .b(new_n125), .c(new_n128), .out0(new_n132));
  aoai13aa1n02x5               g037(.a(new_n131), .b(new_n132), .c(new_n127), .d(new_n124), .o1(\s[10] ));
  nor002aa1n08x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  nand42aa1n04x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nanb02aa1n02x5               g040(.a(new_n134), .b(new_n135), .out0(new_n136));
  aoai13aa1n02x5               g041(.a(new_n129), .b(new_n132), .c(new_n124), .d(new_n127), .o1(new_n137));
  inv040aa1n02x5               g042(.a(new_n134), .o1(new_n138));
  aoai13aa1n06x5               g043(.a(new_n135), .b(new_n132), .c(new_n124), .d(new_n127), .o1(new_n139));
  nano22aa1n02x4               g044(.a(new_n139), .b(new_n129), .c(new_n138), .out0(new_n140));
  aoi012aa1n02x5               g045(.a(new_n140), .b(new_n136), .c(new_n137), .o1(\s[11] ));
  aoai13aa1n06x5               g046(.a(new_n138), .b(new_n139), .c(\b[9] ), .d(\a[10] ), .o1(new_n142));
  xorb03aa1n02x5               g047(.a(new_n142), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1d24x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n08x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nona23aa1n03x5               g050(.a(new_n145), .b(new_n129), .c(new_n128), .d(new_n144), .out0(new_n146));
  nano32aa1n03x7               g051(.a(new_n146), .b(new_n127), .c(new_n138), .d(new_n135), .out0(new_n147));
  aoi022aa1d24x5               g052(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n148));
  oai012aa1n12x5               g053(.a(new_n148), .b(new_n125), .c(new_n128), .o1(new_n149));
  nona22aa1n02x4               g054(.a(new_n149), .b(new_n144), .c(new_n134), .out0(new_n150));
  nanp02aa1n02x5               g055(.a(new_n150), .b(new_n145), .o1(new_n151));
  aob012aa1n03x5               g056(.a(new_n151), .b(new_n124), .c(new_n147), .out0(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor002aa1d32x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand42aa1n08x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  tech160nm_fiaoi012aa1n05x5   g060(.a(new_n154), .b(new_n152), .c(new_n155), .o1(new_n156));
  xnrb03aa1n03x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  inv000aa1d42x5               g062(.a(new_n144), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n145), .o1(new_n159));
  aoi013aa1n09x5               g064(.a(new_n159), .b(new_n149), .c(new_n138), .d(new_n158), .o1(new_n160));
  nor042aa1n06x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nand22aa1n12x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nano23aa1n09x5               g067(.a(new_n154), .b(new_n161), .c(new_n162), .d(new_n155), .out0(new_n163));
  aoai13aa1n06x5               g068(.a(new_n163), .b(new_n160), .c(new_n124), .d(new_n147), .o1(new_n164));
  aoi012aa1n02x5               g069(.a(new_n161), .b(new_n154), .c(new_n162), .o1(new_n165));
  nor042aa1d18x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nand42aa1n20x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  norb02aa1n02x5               g072(.a(new_n167), .b(new_n166), .out0(new_n168));
  xnbna2aa1n03x5               g073(.a(new_n168), .b(new_n164), .c(new_n165), .out0(\s[15] ));
  nanp02aa1n03x5               g074(.a(new_n164), .b(new_n165), .o1(new_n170));
  nor042aa1d18x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nand42aa1n20x5               g076(.a(\b[15] ), .b(\a[16] ), .o1(new_n172));
  nanb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(new_n173));
  aoai13aa1n03x5               g078(.a(new_n173), .b(new_n166), .c(new_n170), .d(new_n167), .o1(new_n174));
  aoi112aa1n03x5               g079(.a(new_n166), .b(new_n173), .c(new_n170), .d(new_n167), .o1(new_n175));
  nanb02aa1n03x5               g080(.a(new_n175), .b(new_n174), .out0(\s[16] ));
  nanb03aa1n06x5               g081(.a(new_n98), .b(new_n99), .c(new_n97), .out0(new_n177));
  norb03aa1n03x5               g082(.a(new_n99), .b(new_n102), .c(new_n101), .out0(new_n178));
  oabi12aa1n06x5               g083(.a(new_n104), .b(new_n178), .c(new_n177), .out0(new_n179));
  xnrc02aa1n06x5               g084(.a(\b[7] ), .b(\a[8] ), .out0(new_n180));
  nor002aa1n04x5               g085(.a(\b[5] ), .b(\a[6] ), .o1(new_n181));
  nor002aa1d32x5               g086(.a(\b[4] ), .b(\a[5] ), .o1(new_n182));
  tech160nm_finor002aa1n03p5x5 g087(.a(new_n182), .b(new_n181), .o1(new_n183));
  aoi012aa1n02x5               g088(.a(new_n117), .b(\a[6] ), .c(\b[5] ), .o1(new_n184));
  nand42aa1n02x5               g089(.a(new_n183), .b(new_n184), .o1(new_n185));
  nor043aa1n02x5               g090(.a(new_n185), .b(new_n180), .c(new_n110), .o1(new_n186));
  nanb03aa1n02x5               g091(.a(new_n117), .b(new_n113), .c(new_n108), .out0(new_n187));
  oai013aa1n02x4               g092(.a(new_n121), .b(new_n187), .c(new_n180), .d(new_n183), .o1(new_n188));
  nano23aa1n02x5               g093(.a(new_n128), .b(new_n144), .c(new_n145), .d(new_n129), .out0(new_n189));
  nano23aa1n02x4               g094(.a(new_n125), .b(new_n134), .c(new_n135), .d(new_n126), .out0(new_n190));
  nano23aa1n02x5               g095(.a(new_n166), .b(new_n171), .c(new_n172), .d(new_n167), .out0(new_n191));
  nand02aa1d04x5               g096(.a(new_n191), .b(new_n163), .o1(new_n192));
  nano22aa1n03x7               g097(.a(new_n192), .b(new_n189), .c(new_n190), .out0(new_n193));
  aoai13aa1n06x5               g098(.a(new_n193), .b(new_n188), .c(new_n179), .d(new_n186), .o1(new_n194));
  nand02aa1n02x5               g099(.a(new_n186), .b(new_n179), .o1(new_n195));
  nona23aa1n03x5               g100(.a(new_n162), .b(new_n155), .c(new_n154), .d(new_n161), .out0(new_n196));
  nona23aa1n03x5               g101(.a(new_n172), .b(new_n167), .c(new_n166), .d(new_n171), .out0(new_n197));
  nor042aa1n03x5               g102(.a(new_n197), .b(new_n196), .o1(new_n198));
  nand22aa1n03x5               g103(.a(new_n147), .b(new_n198), .o1(new_n199));
  inv000aa1d42x5               g104(.a(new_n166), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n171), .o1(new_n201));
  inv000aa1d42x5               g106(.a(new_n172), .o1(new_n202));
  aoai13aa1n04x5               g107(.a(new_n167), .b(new_n161), .c(new_n154), .d(new_n162), .o1(new_n203));
  aoai13aa1n06x5               g108(.a(new_n201), .b(new_n202), .c(new_n203), .d(new_n200), .o1(new_n204));
  aoi012aa1n12x5               g109(.a(new_n204), .b(new_n160), .c(new_n198), .o1(new_n205));
  aoai13aa1n12x5               g110(.a(new_n205), .b(new_n199), .c(new_n195), .d(new_n123), .o1(new_n206));
  xorc02aa1n02x5               g111(.a(\a[17] ), .b(\b[16] ), .out0(new_n207));
  aoi112aa1n02x5               g112(.a(new_n204), .b(new_n207), .c(new_n160), .d(new_n198), .o1(new_n208));
  aoi022aa1n02x5               g113(.a(new_n206), .b(new_n207), .c(new_n194), .d(new_n208), .o1(\s[17] ));
  inv000aa1d42x5               g114(.a(\a[18] ), .o1(new_n210));
  nor042aa1n06x5               g115(.a(\b[16] ), .b(\a[17] ), .o1(new_n211));
  tech160nm_fiaoi012aa1n05x5   g116(.a(new_n211), .b(new_n206), .c(new_n207), .o1(new_n212));
  xorb03aa1n02x5               g117(.a(new_n212), .b(\b[17] ), .c(new_n210), .out0(\s[18] ));
  nand42aa1n03x5               g118(.a(\b[16] ), .b(\a[17] ), .o1(new_n214));
  nor002aa1n02x5               g119(.a(\b[17] ), .b(\a[18] ), .o1(new_n215));
  nand02aa1d06x5               g120(.a(\b[17] ), .b(\a[18] ), .o1(new_n216));
  nano23aa1n06x5               g121(.a(new_n211), .b(new_n215), .c(new_n216), .d(new_n214), .out0(new_n217));
  nand42aa1n02x5               g122(.a(new_n211), .b(new_n216), .o1(new_n218));
  oaib12aa1n06x5               g123(.a(new_n218), .b(\b[17] ), .c(new_n210), .out0(new_n219));
  nor002aa1n16x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nanp02aa1n04x5               g125(.a(\b[18] ), .b(\a[19] ), .o1(new_n221));
  norb02aa1n06x4               g126(.a(new_n221), .b(new_n220), .out0(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n219), .c(new_n206), .d(new_n217), .o1(new_n223));
  aoi112aa1n02x5               g128(.a(new_n222), .b(new_n219), .c(new_n206), .d(new_n217), .o1(new_n224));
  norb02aa1n02x5               g129(.a(new_n223), .b(new_n224), .out0(\s[19] ));
  xnrc02aa1n02x5               g130(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g131(.a(new_n220), .o1(new_n227));
  inv000aa1d42x5               g132(.a(\a[20] ), .o1(new_n228));
  inv000aa1d42x5               g133(.a(\b[19] ), .o1(new_n229));
  nanp02aa1n02x5               g134(.a(new_n229), .b(new_n228), .o1(new_n230));
  nand42aa1n02x5               g135(.a(\b[19] ), .b(\a[20] ), .o1(new_n231));
  nanp02aa1n02x5               g136(.a(new_n230), .b(new_n231), .o1(new_n232));
  aob012aa1n03x5               g137(.a(new_n232), .b(new_n223), .c(new_n227), .out0(new_n233));
  nona22aa1n02x4               g138(.a(new_n223), .b(new_n232), .c(new_n220), .out0(new_n234));
  nanp02aa1n03x5               g139(.a(new_n233), .b(new_n234), .o1(\s[20] ));
  nano22aa1n03x7               g140(.a(new_n232), .b(new_n217), .c(new_n222), .out0(new_n236));
  inv000aa1n03x5               g141(.a(new_n236), .o1(new_n237));
  inv000aa1n02x5               g142(.a(new_n231), .o1(new_n238));
  oai012aa1n02x5               g143(.a(new_n221), .b(\b[19] ), .c(\a[20] ), .o1(new_n239));
  nona32aa1n09x5               g144(.a(new_n219), .b(new_n239), .c(new_n238), .d(new_n220), .out0(new_n240));
  oaoi03aa1n12x5               g145(.a(new_n228), .b(new_n229), .c(new_n220), .o1(new_n241));
  and002aa1n02x5               g146(.a(new_n240), .b(new_n241), .o(new_n242));
  aoai13aa1n04x5               g147(.a(new_n242), .b(new_n237), .c(new_n194), .d(new_n205), .o1(new_n243));
  xorc02aa1n12x5               g148(.a(\a[21] ), .b(\b[20] ), .out0(new_n244));
  nanp02aa1n02x5               g149(.a(new_n240), .b(new_n241), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n244), .b(new_n245), .c(new_n206), .d(new_n236), .o1(new_n246));
  aoi012aa1n02x5               g151(.a(new_n246), .b(new_n243), .c(new_n244), .o1(\s[21] ));
  nor042aa1n04x5               g152(.a(\b[20] ), .b(\a[21] ), .o1(new_n248));
  tech160nm_fixnrc02aa1n04x5   g153(.a(\b[21] ), .b(\a[22] ), .out0(new_n249));
  aoai13aa1n02x5               g154(.a(new_n249), .b(new_n248), .c(new_n243), .d(new_n244), .o1(new_n250));
  aoi112aa1n03x4               g155(.a(new_n248), .b(new_n249), .c(new_n243), .d(new_n244), .o1(new_n251));
  nanb02aa1n03x5               g156(.a(new_n251), .b(new_n250), .out0(\s[22] ));
  oabi12aa1n06x5               g157(.a(new_n204), .b(new_n151), .c(new_n192), .out0(new_n253));
  nanb02aa1n06x5               g158(.a(new_n249), .b(new_n244), .out0(new_n254));
  nano23aa1n02x4               g159(.a(new_n254), .b(new_n232), .c(new_n217), .d(new_n222), .out0(new_n255));
  aoai13aa1n06x5               g160(.a(new_n255), .b(new_n253), .c(new_n124), .d(new_n193), .o1(new_n256));
  inv000aa1d42x5               g161(.a(\a[22] ), .o1(new_n257));
  inv000aa1d42x5               g162(.a(\b[21] ), .o1(new_n258));
  oao003aa1n02x5               g163(.a(new_n257), .b(new_n258), .c(new_n248), .carry(new_n259));
  inv000aa1n02x5               g164(.a(new_n259), .o1(new_n260));
  aoai13aa1n12x5               g165(.a(new_n260), .b(new_n254), .c(new_n240), .d(new_n241), .o1(new_n261));
  nanb02aa1n06x5               g166(.a(new_n261), .b(new_n256), .out0(new_n262));
  xorc02aa1n12x5               g167(.a(\a[23] ), .b(\b[22] ), .out0(new_n263));
  norb02aa1n02x7               g168(.a(new_n244), .b(new_n249), .out0(new_n264));
  aoi112aa1n02x5               g169(.a(new_n263), .b(new_n259), .c(new_n245), .d(new_n264), .o1(new_n265));
  aoi022aa1n02x5               g170(.a(new_n262), .b(new_n263), .c(new_n256), .d(new_n265), .o1(\s[23] ));
  nor042aa1n02x5               g171(.a(\b[22] ), .b(\a[23] ), .o1(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .out0(new_n268));
  aoai13aa1n03x5               g173(.a(new_n268), .b(new_n267), .c(new_n262), .d(new_n263), .o1(new_n269));
  aoai13aa1n02x5               g174(.a(new_n263), .b(new_n261), .c(new_n206), .d(new_n255), .o1(new_n270));
  nona22aa1n02x4               g175(.a(new_n270), .b(new_n268), .c(new_n267), .out0(new_n271));
  nanp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[24] ));
  norb02aa1n03x5               g177(.a(new_n263), .b(new_n268), .out0(new_n273));
  nano22aa1n03x5               g178(.a(new_n237), .b(new_n264), .c(new_n273), .out0(new_n274));
  aoai13aa1n06x5               g179(.a(new_n274), .b(new_n253), .c(new_n124), .d(new_n193), .o1(new_n275));
  nand42aa1n04x5               g180(.a(new_n261), .b(new_n273), .o1(new_n276));
  inv000aa1d42x5               g181(.a(\a[24] ), .o1(new_n277));
  inv000aa1d42x5               g182(.a(\b[23] ), .o1(new_n278));
  oao003aa1n02x5               g183(.a(new_n277), .b(new_n278), .c(new_n267), .carry(new_n279));
  inv000aa1d42x5               g184(.a(new_n279), .o1(new_n280));
  nand42aa1n04x5               g185(.a(new_n276), .b(new_n280), .o1(new_n281));
  nanb02aa1n03x5               g186(.a(new_n281), .b(new_n275), .out0(new_n282));
  tech160nm_fixorc02aa1n03p5x5 g187(.a(\a[25] ), .b(\b[24] ), .out0(new_n283));
  aoi112aa1n02x5               g188(.a(new_n283), .b(new_n279), .c(new_n261), .d(new_n273), .o1(new_n284));
  aoi022aa1n02x5               g189(.a(new_n282), .b(new_n283), .c(new_n275), .d(new_n284), .o1(\s[25] ));
  norp02aa1n02x5               g190(.a(\b[24] ), .b(\a[25] ), .o1(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[25] ), .b(\a[26] ), .out0(new_n287));
  aoai13aa1n03x5               g192(.a(new_n287), .b(new_n286), .c(new_n282), .d(new_n283), .o1(new_n288));
  aoai13aa1n02x5               g193(.a(new_n283), .b(new_n281), .c(new_n206), .d(new_n274), .o1(new_n289));
  nona22aa1n02x4               g194(.a(new_n289), .b(new_n287), .c(new_n286), .out0(new_n290));
  nanp02aa1n03x5               g195(.a(new_n288), .b(new_n290), .o1(\s[26] ));
  norb02aa1n02x5               g196(.a(new_n283), .b(new_n287), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n279), .c(new_n261), .d(new_n273), .o1(new_n293));
  nano32aa1n03x7               g198(.a(new_n237), .b(new_n292), .c(new_n264), .d(new_n273), .out0(new_n294));
  aoai13aa1n03x5               g199(.a(new_n294), .b(new_n253), .c(new_n124), .d(new_n193), .o1(new_n295));
  nanp02aa1n02x5               g200(.a(\b[25] ), .b(\a[26] ), .o1(new_n296));
  oai022aa1n02x5               g201(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n297));
  and002aa1n02x5               g202(.a(new_n297), .b(new_n296), .o(new_n298));
  inv000aa1d42x5               g203(.a(new_n298), .o1(new_n299));
  nand03aa1n02x5               g204(.a(new_n295), .b(new_n293), .c(new_n299), .o1(new_n300));
  xorc02aa1n12x5               g205(.a(\a[27] ), .b(\b[26] ), .out0(new_n301));
  aoi112aa1n02x5               g206(.a(new_n301), .b(new_n298), .c(new_n206), .d(new_n294), .o1(new_n302));
  aoi022aa1n02x5               g207(.a(new_n300), .b(new_n301), .c(new_n302), .d(new_n293), .o1(\s[27] ));
  norp02aa1n02x5               g208(.a(\b[26] ), .b(\a[27] ), .o1(new_n304));
  norp02aa1n02x5               g209(.a(\b[27] ), .b(\a[28] ), .o1(new_n305));
  nanp02aa1n02x5               g210(.a(\b[27] ), .b(\a[28] ), .o1(new_n306));
  nanb02aa1n02x5               g211(.a(new_n305), .b(new_n306), .out0(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n304), .c(new_n300), .d(new_n301), .o1(new_n308));
  nanb02aa1n02x5               g213(.a(new_n287), .b(new_n283), .out0(new_n309));
  aoi012aa1n06x5               g214(.a(new_n309), .b(new_n276), .c(new_n280), .o1(new_n310));
  nona23aa1n02x5               g215(.a(new_n236), .b(new_n273), .c(new_n309), .d(new_n254), .out0(new_n311));
  aoai13aa1n04x5               g216(.a(new_n299), .b(new_n311), .c(new_n194), .d(new_n205), .o1(new_n312));
  oai012aa1n03x5               g217(.a(new_n301), .b(new_n312), .c(new_n310), .o1(new_n313));
  nona22aa1n02x5               g218(.a(new_n313), .b(new_n307), .c(new_n304), .out0(new_n314));
  nanp02aa1n03x5               g219(.a(new_n308), .b(new_n314), .o1(\s[28] ));
  norb02aa1n03x5               g220(.a(new_n301), .b(new_n307), .out0(new_n316));
  oai012aa1n02x5               g221(.a(new_n316), .b(new_n312), .c(new_n310), .o1(new_n317));
  aoi022aa1n09x5               g222(.a(new_n206), .b(new_n294), .c(new_n296), .d(new_n297), .o1(new_n318));
  inv000aa1d42x5               g223(.a(new_n316), .o1(new_n319));
  aoi012aa1n03x5               g224(.a(new_n305), .b(new_n304), .c(new_n306), .o1(new_n320));
  aoai13aa1n03x5               g225(.a(new_n320), .b(new_n319), .c(new_n318), .d(new_n293), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .out0(new_n322));
  norb02aa1n02x5               g227(.a(new_n320), .b(new_n322), .out0(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n317), .d(new_n323), .o1(\s[29] ));
  xorb03aa1n02x5               g229(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g230(.a(new_n307), .b(new_n322), .c(new_n301), .out0(new_n326));
  oabi12aa1n02x5               g231(.a(new_n326), .b(new_n312), .c(new_n310), .out0(new_n327));
  oao003aa1n02x5               g232(.a(\a[29] ), .b(\b[28] ), .c(new_n320), .carry(new_n328));
  aoai13aa1n03x5               g233(.a(new_n328), .b(new_n326), .c(new_n318), .d(new_n293), .o1(new_n329));
  xorc02aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .out0(new_n330));
  norb02aa1n02x5               g235(.a(new_n328), .b(new_n330), .out0(new_n331));
  aoi022aa1n03x5               g236(.a(new_n329), .b(new_n330), .c(new_n327), .d(new_n331), .o1(\s[30] ));
  nand03aa1n02x5               g237(.a(new_n316), .b(new_n322), .c(new_n330), .o1(new_n333));
  oabi12aa1n02x5               g238(.a(new_n333), .b(new_n312), .c(new_n310), .out0(new_n334));
  xorc02aa1n02x5               g239(.a(\a[31] ), .b(\b[30] ), .out0(new_n335));
  inv000aa1d42x5               g240(.a(\a[30] ), .o1(new_n336));
  inv000aa1d42x5               g241(.a(\b[29] ), .o1(new_n337));
  inv000aa1n02x5               g242(.a(new_n328), .o1(new_n338));
  oabi12aa1n02x5               g243(.a(new_n335), .b(\a[30] ), .c(\b[29] ), .out0(new_n339));
  oaoi13aa1n02x5               g244(.a(new_n339), .b(new_n338), .c(new_n336), .d(new_n337), .o1(new_n340));
  oaoi03aa1n02x5               g245(.a(new_n336), .b(new_n337), .c(new_n338), .o1(new_n341));
  aoai13aa1n03x5               g246(.a(new_n341), .b(new_n333), .c(new_n318), .d(new_n293), .o1(new_n342));
  aoi022aa1n03x5               g247(.a(new_n342), .b(new_n335), .c(new_n334), .d(new_n340), .o1(\s[31] ));
  nanb02aa1n02x5               g248(.a(new_n98), .b(new_n97), .out0(new_n344));
  oai012aa1n02x5               g249(.a(new_n99), .b(new_n102), .c(new_n101), .o1(new_n345));
  aoi022aa1n02x5               g250(.a(new_n100), .b(new_n103), .c(new_n345), .d(new_n344), .o1(\s[3] ));
  xorc02aa1n02x5               g251(.a(\a[4] ), .b(\b[3] ), .out0(new_n347));
  aoi112aa1n02x5               g252(.a(new_n347), .b(new_n98), .c(new_n100), .d(new_n103), .o1(new_n348));
  norb02aa1n02x5               g253(.a(new_n109), .b(new_n105), .out0(new_n349));
  oaoi13aa1n02x5               g254(.a(new_n348), .b(new_n349), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  and002aa1n02x5               g255(.a(\b[4] ), .b(\a[5] ), .o(new_n351));
  norp02aa1n02x5               g256(.a(new_n351), .b(new_n182), .o1(new_n352));
  nona23aa1n06x5               g257(.a(new_n179), .b(new_n109), .c(new_n182), .d(new_n351), .out0(new_n353));
  oa0012aa1n02x5               g258(.a(new_n353), .b(new_n349), .c(new_n352), .o(\s[5] ));
  inv000aa1d42x5               g259(.a(new_n182), .o1(new_n355));
  norb02aa1n02x5               g260(.a(new_n113), .b(new_n181), .out0(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n356), .b(new_n353), .c(new_n355), .out0(\s[6] ));
  aob012aa1n02x5               g262(.a(new_n356), .b(new_n353), .c(new_n355), .out0(new_n358));
  tech160nm_fioai012aa1n03p5x5 g263(.a(new_n358), .b(\b[5] ), .c(\a[6] ), .o1(new_n359));
  xorb03aa1n02x5               g264(.a(new_n359), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoai13aa1n02x5               g265(.a(new_n180), .b(new_n117), .c(new_n359), .d(new_n108), .o1(new_n361));
  aoi112aa1n02x5               g266(.a(new_n117), .b(new_n180), .c(new_n359), .d(new_n108), .o1(new_n362));
  nanb02aa1n02x5               g267(.a(new_n362), .b(new_n361), .out0(\s[8] ));
  xorb03aa1n02x5               g268(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


