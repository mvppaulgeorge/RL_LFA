// Benchmark "adder" written by ABC on Thu Jul 18 03:56:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n331,
    new_n334, new_n336, new_n337, new_n338, new_n339, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n04x5               g001(.a(\b[7] ), .b(\a[8] ), .o1(new_n97));
  nanp02aa1n04x5               g002(.a(\b[7] ), .b(\a[8] ), .o1(new_n98));
  nor002aa1d24x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  nanp02aa1n04x5               g004(.a(\b[6] ), .b(\a[7] ), .o1(new_n100));
  nona23aa1n09x5               g005(.a(new_n100), .b(new_n98), .c(new_n97), .d(new_n99), .out0(new_n101));
  inv000aa1d42x5               g006(.a(\a[6] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[5] ), .o1(new_n103));
  nor042aa1n02x5               g008(.a(\b[4] ), .b(\a[5] ), .o1(new_n104));
  tech160nm_fioaoi03aa1n02p5x5 g009(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n105));
  inv000aa1d42x5               g010(.a(new_n99), .o1(new_n106));
  oaoi03aa1n02x5               g011(.a(\a[8] ), .b(\b[7] ), .c(new_n106), .o1(new_n107));
  oabi12aa1n12x5               g012(.a(new_n107), .b(new_n101), .c(new_n105), .out0(new_n108));
  norp02aa1n02x5               g013(.a(\b[3] ), .b(\a[4] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[3] ), .b(\a[4] ), .o1(new_n110));
  nor002aa1n02x5               g015(.a(\b[2] ), .b(\a[3] ), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[2] ), .b(\a[3] ), .o1(new_n112));
  nona23aa1n02x4               g017(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n113));
  inv000aa1d42x5               g018(.a(\a[2] ), .o1(new_n114));
  inv000aa1d42x5               g019(.a(\b[1] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[0] ), .b(\a[1] ), .o1(new_n116));
  tech160nm_fioaoi03aa1n05x5   g021(.a(new_n114), .b(new_n115), .c(new_n116), .o1(new_n117));
  tech160nm_fiao0012aa1n02p5x5 g022(.a(new_n109), .b(new_n111), .c(new_n110), .o(new_n118));
  oabi12aa1n06x5               g023(.a(new_n118), .b(new_n113), .c(new_n117), .out0(new_n119));
  xnrc02aa1n02x5               g024(.a(\b[5] ), .b(\a[6] ), .out0(new_n120));
  xnrc02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .out0(new_n121));
  nor043aa1n02x5               g026(.a(new_n101), .b(new_n120), .c(new_n121), .o1(new_n122));
  aoi012aa1n03x5               g027(.a(new_n108), .b(new_n119), .c(new_n122), .o1(new_n123));
  oaoi03aa1n02x5               g028(.a(\a[9] ), .b(\b[8] ), .c(new_n123), .o1(new_n124));
  xorb03aa1n02x5               g029(.a(new_n124), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor042aa1n06x5               g030(.a(\b[10] ), .b(\a[11] ), .o1(new_n126));
  nand02aa1n04x5               g031(.a(\b[10] ), .b(\a[11] ), .o1(new_n127));
  norb02aa1n02x5               g032(.a(new_n127), .b(new_n126), .out0(new_n128));
  inv000aa1d42x5               g033(.a(new_n128), .o1(new_n129));
  nor042aa1n04x5               g034(.a(\b[8] ), .b(\a[9] ), .o1(new_n130));
  nanp02aa1n02x5               g035(.a(\b[8] ), .b(\a[9] ), .o1(new_n131));
  nor042aa1n04x5               g036(.a(\b[9] ), .b(\a[10] ), .o1(new_n132));
  nand02aa1n04x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  nona23aa1n02x4               g038(.a(new_n133), .b(new_n131), .c(new_n130), .d(new_n132), .out0(new_n134));
  tech160nm_fioai012aa1n03p5x5 g039(.a(new_n133), .b(new_n132), .c(new_n130), .o1(new_n135));
  oaoi13aa1n03x5               g040(.a(new_n129), .b(new_n135), .c(new_n123), .d(new_n134), .o1(new_n136));
  oai112aa1n02x5               g041(.a(new_n135), .b(new_n129), .c(new_n123), .d(new_n134), .o1(new_n137));
  norb02aa1n02x5               g042(.a(new_n137), .b(new_n136), .out0(\s[11] ));
  norp02aa1n03x5               g043(.a(new_n136), .b(new_n126), .o1(new_n139));
  nor002aa1d32x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  inv000aa1d42x5               g045(.a(new_n140), .o1(new_n141));
  nand02aa1n04x5               g046(.a(\b[11] ), .b(\a[12] ), .o1(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n139), .b(new_n142), .c(new_n141), .out0(\s[12] ));
  nona23aa1d18x5               g048(.a(new_n142), .b(new_n127), .c(new_n126), .d(new_n140), .out0(new_n144));
  nor002aa1n02x5               g049(.a(new_n144), .b(new_n134), .o1(new_n145));
  aoai13aa1n06x5               g050(.a(new_n145), .b(new_n108), .c(new_n119), .d(new_n122), .o1(new_n146));
  nand42aa1n03x5               g051(.a(new_n126), .b(new_n142), .o1(new_n147));
  oai112aa1n06x5               g052(.a(new_n147), .b(new_n141), .c(new_n144), .d(new_n135), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  nor042aa1n06x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  nanp02aa1n02x5               g055(.a(\b[12] ), .b(\a[13] ), .o1(new_n151));
  norb02aa1n02x5               g056(.a(new_n151), .b(new_n150), .out0(new_n152));
  xnbna2aa1n03x5               g057(.a(new_n152), .b(new_n146), .c(new_n149), .out0(\s[13] ));
  inv000aa1d42x5               g058(.a(new_n150), .o1(new_n154));
  aob012aa1n02x5               g059(.a(new_n152), .b(new_n146), .c(new_n149), .out0(new_n155));
  norp02aa1n02x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nanp02aa1n02x5               g061(.a(\b[13] ), .b(\a[14] ), .o1(new_n157));
  norb02aa1n02x5               g062(.a(new_n157), .b(new_n156), .out0(new_n158));
  xnbna2aa1n03x5               g063(.a(new_n158), .b(new_n155), .c(new_n154), .out0(\s[14] ));
  nona23aa1n09x5               g064(.a(new_n157), .b(new_n151), .c(new_n150), .d(new_n156), .out0(new_n160));
  oai012aa1n02x5               g065(.a(new_n157), .b(new_n156), .c(new_n150), .o1(new_n161));
  aoai13aa1n02x5               g066(.a(new_n161), .b(new_n160), .c(new_n146), .d(new_n149), .o1(new_n162));
  xorb03aa1n02x5               g067(.a(new_n162), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor002aa1n02x5               g068(.a(\b[14] ), .b(\a[15] ), .o1(new_n164));
  nand42aa1n06x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  norp02aa1n02x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nand42aa1n03x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  aoi112aa1n02x5               g074(.a(new_n169), .b(new_n164), .c(new_n162), .d(new_n166), .o1(new_n170));
  aoai13aa1n03x5               g075(.a(new_n169), .b(new_n164), .c(new_n162), .d(new_n165), .o1(new_n171));
  norb02aa1n02x5               g076(.a(new_n171), .b(new_n170), .out0(\s[16] ));
  nano23aa1n02x4               g077(.a(new_n130), .b(new_n132), .c(new_n133), .d(new_n131), .out0(new_n173));
  nano23aa1n02x4               g078(.a(new_n164), .b(new_n167), .c(new_n168), .d(new_n165), .out0(new_n174));
  nano23aa1n06x5               g079(.a(new_n160), .b(new_n144), .c(new_n174), .d(new_n173), .out0(new_n175));
  aoai13aa1n12x5               g080(.a(new_n175), .b(new_n108), .c(new_n122), .d(new_n119), .o1(new_n176));
  nano22aa1n03x7               g081(.a(new_n160), .b(new_n166), .c(new_n169), .out0(new_n177));
  aoi112aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n178));
  obai22aa1n02x7               g083(.a(new_n174), .b(new_n161), .c(\a[16] ), .d(\b[15] ), .out0(new_n179));
  aoi112aa1n09x5               g084(.a(new_n179), .b(new_n178), .c(new_n148), .d(new_n177), .o1(new_n180));
  xorc02aa1n02x5               g085(.a(\a[17] ), .b(\b[16] ), .out0(new_n181));
  xnbna2aa1n03x5               g086(.a(new_n181), .b(new_n180), .c(new_n176), .out0(\s[17] ));
  inv000aa1d42x5               g087(.a(\a[17] ), .o1(new_n183));
  inv000aa1d42x5               g088(.a(\b[16] ), .o1(new_n184));
  nanp02aa1n02x5               g089(.a(new_n184), .b(new_n183), .o1(new_n185));
  inv000aa1d42x5               g090(.a(new_n108), .o1(new_n186));
  nano23aa1n02x4               g091(.a(new_n109), .b(new_n111), .c(new_n112), .d(new_n110), .out0(new_n187));
  oao003aa1n02x5               g092(.a(new_n114), .b(new_n115), .c(new_n116), .carry(new_n188));
  aoi012aa1n02x5               g093(.a(new_n118), .b(new_n187), .c(new_n188), .o1(new_n189));
  nano23aa1n02x4               g094(.a(new_n97), .b(new_n99), .c(new_n100), .d(new_n98), .out0(new_n190));
  nona22aa1n02x4               g095(.a(new_n190), .b(new_n120), .c(new_n121), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(new_n177), .b(new_n145), .o1(new_n192));
  oaoi13aa1n04x5               g097(.a(new_n192), .b(new_n186), .c(new_n189), .d(new_n191), .o1(new_n193));
  tech160nm_finand02aa1n03p5x5 g098(.a(new_n148), .b(new_n177), .o1(new_n194));
  nano22aa1n02x4               g099(.a(new_n161), .b(new_n166), .c(new_n169), .out0(new_n195));
  nona32aa1n02x5               g100(.a(new_n194), .b(new_n195), .c(new_n178), .d(new_n167), .out0(new_n196));
  oai012aa1n02x5               g101(.a(new_n181), .b(new_n196), .c(new_n193), .o1(new_n197));
  norp02aa1n02x5               g102(.a(\b[17] ), .b(\a[18] ), .o1(new_n198));
  nand42aa1n03x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nanb02aa1n09x5               g104(.a(new_n198), .b(new_n199), .out0(new_n200));
  xobna2aa1n03x5               g105(.a(new_n200), .b(new_n197), .c(new_n185), .out0(\s[18] ));
  nanp02aa1n02x5               g106(.a(\b[16] ), .b(\a[17] ), .o1(new_n202));
  nano22aa1d15x5               g107(.a(new_n200), .b(new_n185), .c(new_n202), .out0(new_n203));
  inv000aa1d42x5               g108(.a(new_n203), .o1(new_n204));
  aoai13aa1n06x5               g109(.a(new_n199), .b(new_n198), .c(new_n183), .d(new_n184), .o1(new_n205));
  aoai13aa1n06x5               g110(.a(new_n205), .b(new_n204), .c(new_n180), .d(new_n176), .o1(new_n206));
  xorb03aa1n03x5               g111(.a(new_n206), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g112(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n12x5               g113(.a(\b[18] ), .b(\a[19] ), .o1(new_n209));
  nand02aa1n03x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nanb02aa1d24x5               g115(.a(new_n209), .b(new_n210), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  inv000aa1d42x5               g117(.a(\a[20] ), .o1(new_n213));
  inv000aa1d42x5               g118(.a(\b[19] ), .o1(new_n214));
  nanp02aa1n02x5               g119(.a(new_n214), .b(new_n213), .o1(new_n215));
  nand42aa1n02x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nand02aa1d06x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoi112aa1n02x7               g123(.a(new_n209), .b(new_n218), .c(new_n206), .d(new_n212), .o1(new_n219));
  inv000aa1d42x5               g124(.a(new_n209), .o1(new_n220));
  nanp02aa1n06x5               g125(.a(new_n206), .b(new_n212), .o1(new_n221));
  aoi012aa1n03x5               g126(.a(new_n217), .b(new_n221), .c(new_n220), .o1(new_n222));
  nor002aa1n02x5               g127(.a(new_n222), .b(new_n219), .o1(\s[20] ));
  nona22aa1n02x4               g128(.a(new_n203), .b(new_n211), .c(new_n217), .out0(new_n224));
  nanp02aa1n02x5               g129(.a(new_n209), .b(new_n216), .o1(new_n225));
  norp03aa1n03x5               g130(.a(new_n205), .b(new_n211), .c(new_n217), .o1(new_n226));
  nano22aa1n03x5               g131(.a(new_n226), .b(new_n215), .c(new_n225), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n224), .c(new_n180), .d(new_n176), .o1(new_n228));
  xorb03aa1n02x5               g133(.a(new_n228), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  xorc02aa1n02x5               g135(.a(\a[21] ), .b(\b[20] ), .out0(new_n231));
  xorc02aa1n12x5               g136(.a(\a[22] ), .b(\b[21] ), .out0(new_n232));
  aoi112aa1n02x7               g137(.a(new_n230), .b(new_n232), .c(new_n228), .d(new_n231), .o1(new_n233));
  inv000aa1d42x5               g138(.a(new_n230), .o1(new_n234));
  nand42aa1n02x5               g139(.a(new_n228), .b(new_n231), .o1(new_n235));
  inv000aa1d42x5               g140(.a(new_n232), .o1(new_n236));
  aoi012aa1n03x5               g141(.a(new_n236), .b(new_n235), .c(new_n234), .o1(new_n237));
  norp02aa1n03x5               g142(.a(new_n237), .b(new_n233), .o1(\s[22] ));
  norp02aa1n02x5               g143(.a(\b[19] ), .b(\a[20] ), .o1(new_n239));
  nona23aa1n06x5               g144(.a(new_n216), .b(new_n210), .c(new_n209), .d(new_n239), .out0(new_n240));
  oai112aa1n02x5               g145(.a(new_n225), .b(new_n215), .c(new_n240), .d(new_n205), .o1(new_n241));
  and002aa1n02x5               g146(.a(new_n232), .b(new_n231), .o(new_n242));
  oaoi03aa1n02x5               g147(.a(\a[22] ), .b(\b[21] ), .c(new_n234), .o1(new_n243));
  aoi012aa1n02x5               g148(.a(new_n243), .b(new_n241), .c(new_n242), .o1(new_n244));
  nona23aa1n03x5               g149(.a(new_n231), .b(new_n203), .c(new_n236), .d(new_n240), .out0(new_n245));
  aoai13aa1n06x5               g150(.a(new_n244), .b(new_n245), .c(new_n180), .d(new_n176), .o1(new_n246));
  xorb03aa1n02x5               g151(.a(new_n246), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n06x5               g152(.a(\b[22] ), .b(\a[23] ), .o1(new_n248));
  tech160nm_finand02aa1n03p5x5 g153(.a(\b[22] ), .b(\a[23] ), .o1(new_n249));
  norb02aa1n02x5               g154(.a(new_n249), .b(new_n248), .out0(new_n250));
  nor042aa1n02x5               g155(.a(\b[23] ), .b(\a[24] ), .o1(new_n251));
  nand42aa1n02x5               g156(.a(\b[23] ), .b(\a[24] ), .o1(new_n252));
  norb02aa1n02x5               g157(.a(new_n252), .b(new_n251), .out0(new_n253));
  aoi112aa1n02x7               g158(.a(new_n248), .b(new_n253), .c(new_n246), .d(new_n250), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n248), .o1(new_n255));
  nand42aa1n02x5               g160(.a(new_n246), .b(new_n250), .o1(new_n256));
  inv000aa1d42x5               g161(.a(new_n253), .o1(new_n257));
  aoi012aa1n03x5               g162(.a(new_n257), .b(new_n256), .c(new_n255), .o1(new_n258));
  nor002aa1n02x5               g163(.a(new_n258), .b(new_n254), .o1(\s[24] ));
  nano23aa1d15x5               g164(.a(new_n248), .b(new_n251), .c(new_n252), .d(new_n249), .out0(new_n260));
  inv000aa1d42x5               g165(.a(new_n260), .o1(new_n261));
  nona23aa1n02x4               g166(.a(new_n242), .b(new_n203), .c(new_n261), .d(new_n240), .out0(new_n262));
  aoi112aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n263));
  aoi112aa1n02x7               g168(.a(new_n263), .b(new_n251), .c(new_n260), .d(new_n243), .o1(new_n264));
  nand03aa1n02x5               g169(.a(new_n260), .b(new_n231), .c(new_n232), .o1(new_n265));
  tech160nm_fioai012aa1n05x5   g170(.a(new_n264), .b(new_n227), .c(new_n265), .o1(new_n266));
  inv040aa1n03x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n262), .c(new_n180), .d(new_n176), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  xorc02aa1n12x5               g176(.a(\a[26] ), .b(\b[25] ), .out0(new_n272));
  aoi112aa1n03x4               g177(.a(new_n270), .b(new_n272), .c(new_n268), .d(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n270), .o1(new_n274));
  nand42aa1n02x5               g179(.a(new_n268), .b(new_n271), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n272), .o1(new_n276));
  aoi012aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .o1(new_n277));
  nor002aa1n02x5               g182(.a(new_n277), .b(new_n273), .o1(\s[26] ));
  and002aa1n02x5               g183(.a(new_n272), .b(new_n271), .o(new_n279));
  nano22aa1n03x7               g184(.a(new_n245), .b(new_n260), .c(new_n279), .out0(new_n280));
  oai012aa1n06x5               g185(.a(new_n280), .b(new_n196), .c(new_n193), .o1(new_n281));
  norp02aa1n02x5               g186(.a(\b[25] ), .b(\a[26] ), .o1(new_n282));
  aoi112aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .c(\a[26] ), .d(\b[25] ), .o1(new_n283));
  aoi112aa1n06x5               g188(.a(new_n282), .b(new_n283), .c(new_n266), .d(new_n279), .o1(new_n284));
  xorc02aa1n12x5               g189(.a(\a[27] ), .b(\b[26] ), .out0(new_n285));
  xnbna2aa1n03x5               g190(.a(new_n285), .b(new_n281), .c(new_n284), .out0(\s[27] ));
  nor042aa1n03x5               g191(.a(\b[26] ), .b(\a[27] ), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n287), .o1(new_n288));
  inv000aa1d42x5               g193(.a(new_n285), .o1(new_n289));
  tech160nm_fiaoi012aa1n02p5x5 g194(.a(new_n289), .b(new_n281), .c(new_n284), .o1(new_n290));
  xnrc02aa1n02x5               g195(.a(\b[27] ), .b(\a[28] ), .out0(new_n291));
  nano22aa1n03x5               g196(.a(new_n290), .b(new_n288), .c(new_n291), .out0(new_n292));
  nand02aa1d06x5               g197(.a(new_n180), .b(new_n176), .o1(new_n293));
  nanp02aa1n02x5               g198(.a(new_n260), .b(new_n243), .o1(new_n294));
  nona22aa1n02x4               g199(.a(new_n294), .b(new_n263), .c(new_n251), .out0(new_n295));
  inv040aa1n03x5               g200(.a(new_n265), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n279), .b(new_n295), .c(new_n241), .d(new_n296), .o1(new_n297));
  nona22aa1n02x5               g202(.a(new_n297), .b(new_n283), .c(new_n282), .out0(new_n298));
  aoai13aa1n03x5               g203(.a(new_n285), .b(new_n298), .c(new_n293), .d(new_n280), .o1(new_n299));
  aoi012aa1n03x5               g204(.a(new_n291), .b(new_n299), .c(new_n288), .o1(new_n300));
  nor002aa1n02x5               g205(.a(new_n300), .b(new_n292), .o1(\s[28] ));
  norb02aa1n02x5               g206(.a(new_n285), .b(new_n291), .out0(new_n302));
  aoai13aa1n06x5               g207(.a(new_n302), .b(new_n298), .c(new_n293), .d(new_n280), .o1(new_n303));
  oao003aa1n02x5               g208(.a(\a[28] ), .b(\b[27] ), .c(new_n288), .carry(new_n304));
  xnrc02aa1n02x5               g209(.a(\b[28] ), .b(\a[29] ), .out0(new_n305));
  tech160nm_fiaoi012aa1n05x5   g210(.a(new_n305), .b(new_n303), .c(new_n304), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n302), .o1(new_n307));
  tech160nm_fiaoi012aa1n05x5   g212(.a(new_n307), .b(new_n281), .c(new_n284), .o1(new_n308));
  nano22aa1n02x5               g213(.a(new_n308), .b(new_n304), .c(new_n305), .out0(new_n309));
  norp02aa1n03x5               g214(.a(new_n306), .b(new_n309), .o1(\s[29] ));
  xorb03aa1n02x5               g215(.a(new_n116), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n03x5               g216(.a(new_n285), .b(new_n305), .c(new_n291), .out0(new_n312));
  aoai13aa1n03x5               g217(.a(new_n312), .b(new_n298), .c(new_n293), .d(new_n280), .o1(new_n313));
  oao003aa1n02x5               g218(.a(\a[29] ), .b(\b[28] ), .c(new_n304), .carry(new_n314));
  xnrc02aa1n02x5               g219(.a(\b[29] ), .b(\a[30] ), .out0(new_n315));
  aoi012aa1n03x5               g220(.a(new_n315), .b(new_n313), .c(new_n314), .o1(new_n316));
  inv000aa1d42x5               g221(.a(new_n312), .o1(new_n317));
  aoi012aa1n02x7               g222(.a(new_n317), .b(new_n281), .c(new_n284), .o1(new_n318));
  nano22aa1n03x5               g223(.a(new_n318), .b(new_n314), .c(new_n315), .out0(new_n319));
  norp02aa1n03x5               g224(.a(new_n316), .b(new_n319), .o1(\s[30] ));
  norb02aa1n06x5               g225(.a(new_n312), .b(new_n315), .out0(new_n321));
  inv000aa1d42x5               g226(.a(new_n321), .o1(new_n322));
  tech160nm_fiaoi012aa1n02p5x5 g227(.a(new_n322), .b(new_n281), .c(new_n284), .o1(new_n323));
  oao003aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .c(new_n314), .carry(new_n324));
  xnrc02aa1n02x5               g229(.a(\b[30] ), .b(\a[31] ), .out0(new_n325));
  nano22aa1n02x4               g230(.a(new_n323), .b(new_n324), .c(new_n325), .out0(new_n326));
  aoai13aa1n03x5               g231(.a(new_n321), .b(new_n298), .c(new_n293), .d(new_n280), .o1(new_n327));
  aoi012aa1n03x5               g232(.a(new_n325), .b(new_n327), .c(new_n324), .o1(new_n328));
  norp02aa1n03x5               g233(.a(new_n328), .b(new_n326), .o1(\s[31] ));
  xnrb03aa1n02x5               g234(.a(new_n117), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g235(.a(\a[3] ), .b(\b[2] ), .c(new_n117), .o1(new_n331));
  xorb03aa1n02x5               g236(.a(new_n331), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g237(.a(new_n119), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  aoib12aa1n02x5               g238(.a(new_n104), .b(new_n119), .c(new_n121), .out0(new_n334));
  xorb03aa1n02x5               g239(.a(new_n334), .b(\b[5] ), .c(new_n102), .out0(\s[6] ));
  norb02aa1n02x5               g240(.a(new_n100), .b(new_n99), .out0(new_n336));
  nanb02aa1n02x5               g241(.a(new_n120), .b(new_n334), .out0(new_n337));
  oai112aa1n02x5               g242(.a(new_n337), .b(new_n336), .c(new_n103), .d(new_n102), .o1(new_n338));
  oaoi13aa1n02x5               g243(.a(new_n336), .b(new_n337), .c(new_n102), .d(new_n103), .o1(new_n339));
  norb02aa1n02x5               g244(.a(new_n338), .b(new_n339), .out0(\s[7] ));
  norb02aa1n02x5               g245(.a(new_n98), .b(new_n97), .out0(new_n341));
  xnbna2aa1n03x5               g246(.a(new_n341), .b(new_n338), .c(new_n106), .out0(\s[8] ));
  xnrb03aa1n02x5               g247(.a(new_n123), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


