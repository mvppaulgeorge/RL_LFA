// Benchmark "adder" written by ABC on Thu Jul 18 14:47:01 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n160, new_n161, new_n162, new_n163, new_n164, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n174,
    new_n175, new_n176, new_n177, new_n179, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n309, new_n312,
    new_n313, new_n315, new_n316, new_n317, new_n318, new_n319, new_n321;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nand42aa1n02x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand22aa1n06x5               g002(.a(\b[0] ), .b(\a[1] ), .o1(new_n98));
  nor002aa1n03x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  oai012aa1n09x5               g004(.a(new_n97), .b(new_n99), .c(new_n98), .o1(new_n100));
  tech160nm_fixnrc02aa1n04x5   g005(.a(\b[3] ), .b(\a[4] ), .out0(new_n101));
  inv000aa1d42x5               g006(.a(\a[3] ), .o1(new_n102));
  nanb02aa1n12x5               g007(.a(\b[2] ), .b(new_n102), .out0(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(new_n103), .b(new_n104), .o1(new_n105));
  oao003aa1n02x5               g010(.a(\a[4] ), .b(\b[3] ), .c(new_n103), .carry(new_n106));
  oai013aa1n09x5               g011(.a(new_n106), .b(new_n101), .c(new_n100), .d(new_n105), .o1(new_n107));
  xnrc02aa1n02x5               g012(.a(\b[5] ), .b(\a[6] ), .out0(new_n108));
  norp02aa1n09x5               g013(.a(\b[7] ), .b(\a[8] ), .o1(new_n109));
  nand02aa1n04x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nor002aa1d32x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nanp02aa1n04x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nona23aa1d18x5               g017(.a(new_n112), .b(new_n110), .c(new_n109), .d(new_n111), .out0(new_n113));
  xnrc02aa1n02x5               g018(.a(\b[4] ), .b(\a[5] ), .out0(new_n114));
  nor043aa1n03x5               g019(.a(new_n113), .b(new_n114), .c(new_n108), .o1(new_n115));
  tech160nm_fioai012aa1n03p5x5 g020(.a(new_n110), .b(new_n111), .c(new_n109), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\a[6] ), .o1(new_n117));
  oai022aa1n02x7               g022(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n118));
  oaib12aa1n06x5               g023(.a(new_n118), .b(new_n117), .c(\b[5] ), .out0(new_n119));
  oai012aa1d24x5               g024(.a(new_n116), .b(new_n113), .c(new_n119), .o1(new_n120));
  aoi012aa1n12x5               g025(.a(new_n120), .b(new_n107), .c(new_n115), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[9] ), .b(\b[8] ), .c(new_n121), .o1(new_n122));
  xorb03aa1n02x5               g027(.a(new_n122), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n06x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  nand02aa1n03x5               g029(.a(\b[10] ), .b(\a[11] ), .o1(new_n125));
  norb02aa1n02x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  inv000aa1n02x5               g031(.a(new_n126), .o1(new_n127));
  nor042aa1n04x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  nor002aa1n04x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  oai012aa1n12x5               g035(.a(new_n130), .b(new_n129), .c(new_n128), .o1(new_n131));
  nanp02aa1n02x5               g036(.a(\b[8] ), .b(\a[9] ), .o1(new_n132));
  nona23aa1n09x5               g037(.a(new_n130), .b(new_n132), .c(new_n128), .d(new_n129), .out0(new_n133));
  oaoi13aa1n02x5               g038(.a(new_n127), .b(new_n131), .c(new_n121), .d(new_n133), .o1(new_n134));
  oai112aa1n02x5               g039(.a(new_n131), .b(new_n127), .c(new_n121), .d(new_n133), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(\s[11] ));
  norp02aa1n02x5               g041(.a(new_n134), .b(new_n124), .o1(new_n137));
  xnrb03aa1n03x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor002aa1n03x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nand22aa1n03x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nona23aa1n09x5               g045(.a(new_n140), .b(new_n125), .c(new_n124), .d(new_n139), .out0(new_n141));
  norp02aa1n02x5               g046(.a(new_n141), .b(new_n133), .o1(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n120), .c(new_n107), .d(new_n115), .o1(new_n143));
  ao0012aa1n03x7               g048(.a(new_n139), .b(new_n124), .c(new_n140), .o(new_n144));
  oabi12aa1n18x5               g049(.a(new_n144), .b(new_n141), .c(new_n131), .out0(new_n145));
  inv000aa1d42x5               g050(.a(new_n145), .o1(new_n146));
  xnrc02aa1n12x5               g051(.a(\b[12] ), .b(\a[13] ), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n143), .c(new_n146), .out0(\s[13] ));
  orn002aa1n02x7               g054(.a(\a[13] ), .b(\b[12] ), .o(new_n150));
  aoai13aa1n02x5               g055(.a(new_n150), .b(new_n147), .c(new_n143), .d(new_n146), .o1(new_n151));
  xorb03aa1n02x5               g056(.a(new_n151), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  xnrc02aa1n02x5               g057(.a(\b[13] ), .b(\a[14] ), .out0(new_n153));
  nor042aa1n09x5               g058(.a(new_n153), .b(new_n147), .o1(new_n154));
  inv000aa1d42x5               g059(.a(new_n154), .o1(new_n155));
  tech160nm_fioaoi03aa1n02p5x5 g060(.a(\a[14] ), .b(\b[13] ), .c(new_n150), .o1(new_n156));
  inv000aa1n02x5               g061(.a(new_n156), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n155), .c(new_n143), .d(new_n146), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  inv000aa1d42x5               g064(.a(\a[16] ), .o1(new_n160));
  norp02aa1n02x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  xnrc02aa1n12x5               g066(.a(\b[14] ), .b(\a[15] ), .out0(new_n162));
  inv000aa1d42x5               g067(.a(new_n162), .o1(new_n163));
  aoi012aa1n02x5               g068(.a(new_n161), .b(new_n158), .c(new_n163), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[15] ), .c(new_n160), .out0(\s[16] ));
  xnrc02aa1n02x5               g070(.a(\b[15] ), .b(\a[16] ), .out0(new_n166));
  nor042aa1n02x5               g071(.a(new_n166), .b(new_n162), .o1(new_n167));
  nona23aa1n09x5               g072(.a(new_n154), .b(new_n167), .c(new_n141), .d(new_n133), .out0(new_n168));
  aoai13aa1n06x5               g073(.a(new_n167), .b(new_n156), .c(new_n145), .d(new_n154), .o1(new_n169));
  aoi112aa1n02x5               g074(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n170));
  aoib12aa1n02x5               g075(.a(new_n170), .b(new_n160), .c(\b[15] ), .out0(new_n171));
  oai112aa1n06x5               g076(.a(new_n169), .b(new_n171), .c(new_n121), .d(new_n168), .o1(new_n172));
  xorb03aa1n02x5               g077(.a(new_n172), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g078(.a(\a[18] ), .o1(new_n174));
  inv000aa1d42x5               g079(.a(\a[17] ), .o1(new_n175));
  inv000aa1d42x5               g080(.a(\b[16] ), .o1(new_n176));
  oaoi03aa1n03x5               g081(.a(new_n175), .b(new_n176), .c(new_n172), .o1(new_n177));
  xorb03aa1n02x5               g082(.a(new_n177), .b(\b[17] ), .c(new_n174), .out0(\s[18] ));
  nanp02aa1n02x5               g083(.a(new_n107), .b(new_n115), .o1(new_n179));
  inv000aa1d42x5               g084(.a(new_n120), .o1(new_n180));
  aoi012aa1n09x5               g085(.a(new_n168), .b(new_n179), .c(new_n180), .o1(new_n181));
  inv000aa1n02x5               g086(.a(new_n167), .o1(new_n182));
  inv030aa1n02x5               g087(.a(new_n131), .o1(new_n183));
  nano23aa1n03x7               g088(.a(new_n124), .b(new_n139), .c(new_n140), .d(new_n125), .out0(new_n184));
  aoai13aa1n04x5               g089(.a(new_n154), .b(new_n144), .c(new_n184), .d(new_n183), .o1(new_n185));
  aoai13aa1n06x5               g090(.a(new_n171), .b(new_n182), .c(new_n185), .d(new_n157), .o1(new_n186));
  xroi22aa1d06x4               g091(.a(new_n175), .b(\b[16] ), .c(new_n174), .d(\b[17] ), .out0(new_n187));
  tech160nm_fioai012aa1n03p5x5 g092(.a(new_n187), .b(new_n186), .c(new_n181), .o1(new_n188));
  oai022aa1n02x7               g093(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n189));
  oaib12aa1n06x5               g094(.a(new_n189), .b(new_n174), .c(\b[17] ), .out0(new_n190));
  nor042aa1n09x5               g095(.a(\b[18] ), .b(\a[19] ), .o1(new_n191));
  nand22aa1n03x5               g096(.a(\b[18] ), .b(\a[19] ), .o1(new_n192));
  nanb02aa1n02x5               g097(.a(new_n191), .b(new_n192), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  xnbna2aa1n03x5               g099(.a(new_n194), .b(new_n188), .c(new_n190), .out0(\s[19] ));
  xnrc02aa1n02x5               g100(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g101(.a(new_n191), .o1(new_n197));
  aoi012aa1n02x7               g102(.a(new_n193), .b(new_n188), .c(new_n190), .o1(new_n198));
  nor002aa1n04x5               g103(.a(\b[19] ), .b(\a[20] ), .o1(new_n199));
  nand02aa1d04x5               g104(.a(\b[19] ), .b(\a[20] ), .o1(new_n200));
  nanb02aa1n02x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  nano22aa1n03x5               g106(.a(new_n198), .b(new_n197), .c(new_n201), .out0(new_n202));
  nanp02aa1n02x5               g107(.a(new_n176), .b(new_n175), .o1(new_n203));
  oaoi03aa1n02x5               g108(.a(\a[18] ), .b(\b[17] ), .c(new_n203), .o1(new_n204));
  aoai13aa1n03x5               g109(.a(new_n194), .b(new_n204), .c(new_n172), .d(new_n187), .o1(new_n205));
  aoi012aa1n03x5               g110(.a(new_n201), .b(new_n205), .c(new_n197), .o1(new_n206));
  nor002aa1n02x5               g111(.a(new_n206), .b(new_n202), .o1(\s[20] ));
  nano23aa1n06x5               g112(.a(new_n191), .b(new_n199), .c(new_n200), .d(new_n192), .out0(new_n208));
  nand02aa1d04x5               g113(.a(new_n187), .b(new_n208), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  oaih12aa1n02x5               g115(.a(new_n210), .b(new_n186), .c(new_n181), .o1(new_n211));
  nona23aa1d18x5               g116(.a(new_n200), .b(new_n192), .c(new_n191), .d(new_n199), .out0(new_n212));
  aoi012aa1n09x5               g117(.a(new_n199), .b(new_n191), .c(new_n200), .o1(new_n213));
  oai012aa1d24x5               g118(.a(new_n213), .b(new_n212), .c(new_n190), .o1(new_n214));
  inv000aa1d42x5               g119(.a(new_n214), .o1(new_n215));
  nor002aa1d32x5               g120(.a(\b[20] ), .b(\a[21] ), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(\b[20] ), .b(\a[21] ), .o1(new_n217));
  norb02aa1n02x5               g122(.a(new_n217), .b(new_n216), .out0(new_n218));
  xnbna2aa1n03x5               g123(.a(new_n218), .b(new_n211), .c(new_n215), .out0(\s[21] ));
  inv000aa1d42x5               g124(.a(new_n216), .o1(new_n220));
  aobi12aa1n02x5               g125(.a(new_n218), .b(new_n211), .c(new_n215), .out0(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[21] ), .b(\a[22] ), .out0(new_n222));
  nano22aa1n02x4               g127(.a(new_n221), .b(new_n220), .c(new_n222), .out0(new_n223));
  aoai13aa1n03x5               g128(.a(new_n218), .b(new_n214), .c(new_n172), .d(new_n210), .o1(new_n224));
  aoi012aa1n03x5               g129(.a(new_n222), .b(new_n224), .c(new_n220), .o1(new_n225));
  nor002aa1n02x5               g130(.a(new_n225), .b(new_n223), .o1(\s[22] ));
  nano22aa1n03x7               g131(.a(new_n222), .b(new_n220), .c(new_n217), .out0(new_n227));
  and003aa1n02x5               g132(.a(new_n187), .b(new_n227), .c(new_n208), .o(new_n228));
  oaih12aa1n02x5               g133(.a(new_n228), .b(new_n186), .c(new_n181), .o1(new_n229));
  oao003aa1n06x5               g134(.a(\a[22] ), .b(\b[21] ), .c(new_n220), .carry(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  aoi012aa1n06x5               g136(.a(new_n231), .b(new_n214), .c(new_n227), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[22] ), .b(\a[23] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnbna2aa1n03x5               g139(.a(new_n234), .b(new_n229), .c(new_n232), .out0(\s[23] ));
  nor042aa1n03x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi012aa1n03x5               g142(.a(new_n233), .b(new_n229), .c(new_n232), .o1(new_n238));
  xnrc02aa1n02x5               g143(.a(\b[23] ), .b(\a[24] ), .out0(new_n239));
  nano22aa1n02x4               g144(.a(new_n238), .b(new_n237), .c(new_n239), .out0(new_n240));
  inv000aa1n02x5               g145(.a(new_n232), .o1(new_n241));
  aoai13aa1n03x5               g146(.a(new_n234), .b(new_n241), .c(new_n172), .d(new_n228), .o1(new_n242));
  aoi012aa1n03x5               g147(.a(new_n239), .b(new_n242), .c(new_n237), .o1(new_n243));
  nor002aa1n02x5               g148(.a(new_n243), .b(new_n240), .o1(\s[24] ));
  nor002aa1n02x5               g149(.a(new_n239), .b(new_n233), .o1(new_n245));
  nano22aa1n03x7               g150(.a(new_n209), .b(new_n227), .c(new_n245), .out0(new_n246));
  oaih12aa1n02x5               g151(.a(new_n246), .b(new_n186), .c(new_n181), .o1(new_n247));
  inv040aa1n02x5               g152(.a(new_n213), .o1(new_n248));
  aoai13aa1n06x5               g153(.a(new_n227), .b(new_n248), .c(new_n208), .d(new_n204), .o1(new_n249));
  inv000aa1n02x5               g154(.a(new_n245), .o1(new_n250));
  oao003aa1n02x5               g155(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .carry(new_n251));
  aoai13aa1n06x5               g156(.a(new_n251), .b(new_n250), .c(new_n249), .d(new_n230), .o1(new_n252));
  xnrc02aa1n12x5               g157(.a(\b[24] ), .b(\a[25] ), .out0(new_n253));
  aoib12aa1n06x5               g158(.a(new_n253), .b(new_n247), .c(new_n252), .out0(new_n254));
  inv000aa1d42x5               g159(.a(new_n253), .o1(new_n255));
  aoi112aa1n02x5               g160(.a(new_n255), .b(new_n252), .c(new_n172), .d(new_n246), .o1(new_n256));
  norp02aa1n02x5               g161(.a(new_n254), .b(new_n256), .o1(\s[25] ));
  nor042aa1n03x5               g162(.a(\b[24] ), .b(\a[25] ), .o1(new_n258));
  inv000aa1d42x5               g163(.a(new_n258), .o1(new_n259));
  xnrc02aa1n02x5               g164(.a(\b[25] ), .b(\a[26] ), .out0(new_n260));
  nano22aa1n03x7               g165(.a(new_n254), .b(new_n259), .c(new_n260), .out0(new_n261));
  aoai13aa1n03x5               g166(.a(new_n255), .b(new_n252), .c(new_n172), .d(new_n246), .o1(new_n262));
  aoi012aa1n03x5               g167(.a(new_n260), .b(new_n262), .c(new_n259), .o1(new_n263));
  nor002aa1n02x5               g168(.a(new_n263), .b(new_n261), .o1(\s[26] ));
  nor042aa1n03x5               g169(.a(new_n260), .b(new_n253), .o1(new_n265));
  nano32aa1n03x7               g170(.a(new_n209), .b(new_n265), .c(new_n227), .d(new_n245), .out0(new_n266));
  oai012aa1n06x5               g171(.a(new_n266), .b(new_n186), .c(new_n181), .o1(new_n267));
  oao003aa1n03x5               g172(.a(\a[26] ), .b(\b[25] ), .c(new_n259), .carry(new_n268));
  aobi12aa1n06x5               g173(.a(new_n268), .b(new_n252), .c(new_n265), .out0(new_n269));
  xorc02aa1n02x5               g174(.a(\a[27] ), .b(\b[26] ), .out0(new_n270));
  xnbna2aa1n03x5               g175(.a(new_n270), .b(new_n267), .c(new_n269), .out0(\s[27] ));
  norp02aa1n02x5               g176(.a(\b[26] ), .b(\a[27] ), .o1(new_n272));
  inv040aa1n03x5               g177(.a(new_n272), .o1(new_n273));
  aobi12aa1n03x5               g178(.a(new_n270), .b(new_n267), .c(new_n269), .out0(new_n274));
  xnrc02aa1n02x5               g179(.a(\b[27] ), .b(\a[28] ), .out0(new_n275));
  nano22aa1n03x5               g180(.a(new_n274), .b(new_n273), .c(new_n275), .out0(new_n276));
  aoai13aa1n03x5               g181(.a(new_n245), .b(new_n231), .c(new_n214), .d(new_n227), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n265), .o1(new_n278));
  aoai13aa1n04x5               g183(.a(new_n268), .b(new_n278), .c(new_n277), .d(new_n251), .o1(new_n279));
  aoai13aa1n03x5               g184(.a(new_n270), .b(new_n279), .c(new_n172), .d(new_n266), .o1(new_n280));
  aoi012aa1n03x5               g185(.a(new_n275), .b(new_n280), .c(new_n273), .o1(new_n281));
  nor002aa1n02x5               g186(.a(new_n281), .b(new_n276), .o1(\s[28] ));
  norb02aa1n02x5               g187(.a(new_n270), .b(new_n275), .out0(new_n283));
  aobi12aa1n03x5               g188(.a(new_n283), .b(new_n267), .c(new_n269), .out0(new_n284));
  oao003aa1n02x5               g189(.a(\a[28] ), .b(\b[27] ), .c(new_n273), .carry(new_n285));
  xnrc02aa1n02x5               g190(.a(\b[28] ), .b(\a[29] ), .out0(new_n286));
  nano22aa1n03x5               g191(.a(new_n284), .b(new_n285), .c(new_n286), .out0(new_n287));
  aoai13aa1n02x7               g192(.a(new_n283), .b(new_n279), .c(new_n172), .d(new_n266), .o1(new_n288));
  aoi012aa1n03x5               g193(.a(new_n286), .b(new_n288), .c(new_n285), .o1(new_n289));
  norp02aa1n03x5               g194(.a(new_n289), .b(new_n287), .o1(\s[29] ));
  xorb03aa1n02x5               g195(.a(new_n98), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g196(.a(new_n270), .b(new_n286), .c(new_n275), .out0(new_n292));
  aobi12aa1n06x5               g197(.a(new_n292), .b(new_n267), .c(new_n269), .out0(new_n293));
  oao003aa1n03x5               g198(.a(\a[29] ), .b(\b[28] ), .c(new_n285), .carry(new_n294));
  xnrc02aa1n02x5               g199(.a(\b[29] ), .b(\a[30] ), .out0(new_n295));
  nano22aa1n03x7               g200(.a(new_n293), .b(new_n294), .c(new_n295), .out0(new_n296));
  aoai13aa1n03x5               g201(.a(new_n292), .b(new_n279), .c(new_n172), .d(new_n266), .o1(new_n297));
  aoi012aa1n03x5               g202(.a(new_n295), .b(new_n297), .c(new_n294), .o1(new_n298));
  nor002aa1n02x5               g203(.a(new_n298), .b(new_n296), .o1(\s[30] ));
  xnrc02aa1n02x5               g204(.a(\b[30] ), .b(\a[31] ), .out0(new_n300));
  norb02aa1n02x5               g205(.a(new_n292), .b(new_n295), .out0(new_n301));
  aobi12aa1n03x5               g206(.a(new_n301), .b(new_n267), .c(new_n269), .out0(new_n302));
  oao003aa1n02x5               g207(.a(\a[30] ), .b(\b[29] ), .c(new_n294), .carry(new_n303));
  nano22aa1n03x5               g208(.a(new_n302), .b(new_n300), .c(new_n303), .out0(new_n304));
  aoai13aa1n02x7               g209(.a(new_n301), .b(new_n279), .c(new_n172), .d(new_n266), .o1(new_n305));
  aoi012aa1n02x5               g210(.a(new_n300), .b(new_n305), .c(new_n303), .o1(new_n306));
  nor002aa1n02x5               g211(.a(new_n306), .b(new_n304), .o1(\s[31] ));
  xnbna2aa1n03x5               g212(.a(new_n100), .b(new_n104), .c(new_n103), .out0(\s[3] ));
  oaoi03aa1n02x5               g213(.a(\a[3] ), .b(\b[2] ), .c(new_n100), .o1(new_n309));
  xorb03aa1n02x5               g214(.a(new_n309), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g215(.a(new_n107), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norp02aa1n02x5               g216(.a(\b[4] ), .b(\a[5] ), .o1(new_n312));
  aoib12aa1n06x5               g217(.a(new_n312), .b(new_n107), .c(new_n114), .out0(new_n313));
  xorb03aa1n02x5               g218(.a(new_n313), .b(\b[5] ), .c(new_n117), .out0(\s[6] ));
  and002aa1n02x5               g219(.a(\b[5] ), .b(\a[6] ), .o(new_n315));
  nanb02aa1n02x5               g220(.a(new_n108), .b(new_n313), .out0(new_n316));
  nona23aa1n03x5               g221(.a(new_n316), .b(new_n112), .c(new_n315), .d(new_n111), .out0(new_n317));
  inv000aa1d42x5               g222(.a(new_n111), .o1(new_n318));
  aboi22aa1n03x5               g223(.a(new_n315), .b(new_n316), .c(new_n318), .d(new_n112), .out0(new_n319));
  norb02aa1n02x5               g224(.a(new_n317), .b(new_n319), .out0(\s[7] ));
  norb02aa1n02x5               g225(.a(new_n110), .b(new_n109), .out0(new_n321));
  xnbna2aa1n03x5               g226(.a(new_n321), .b(new_n317), .c(new_n318), .out0(\s[8] ));
  xnrb03aa1n02x5               g227(.a(new_n121), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


