// Benchmark "adder" written by ABC on Thu Jul 18 02:13:00 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n327, new_n329, new_n332, new_n333,
    new_n335, new_n337;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  inv040aa1d30x5               g002(.a(\b[8] ), .o1(new_n98));
  nanp02aa1n02x5               g003(.a(new_n98), .b(new_n97), .o1(new_n99));
  nand22aa1n06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  nand42aa1n02x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  nor042aa1n04x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  oai112aa1n04x5               g008(.a(new_n103), .b(new_n101), .c(new_n102), .d(new_n100), .o1(new_n104));
  oa0022aa1n09x5               g009(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n105));
  aoi022aa1n12x5               g010(.a(new_n104), .b(new_n105), .c(\b[3] ), .d(\a[4] ), .o1(new_n106));
  nor042aa1n02x5               g011(.a(\b[5] ), .b(\a[6] ), .o1(new_n107));
  nand42aa1n03x5               g012(.a(\b[5] ), .b(\a[6] ), .o1(new_n108));
  norb02aa1n02x7               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  nor042aa1n03x5               g014(.a(\b[7] ), .b(\a[8] ), .o1(new_n110));
  nand02aa1n03x5               g015(.a(\b[7] ), .b(\a[8] ), .o1(new_n111));
  nor042aa1n03x5               g016(.a(\b[6] ), .b(\a[7] ), .o1(new_n112));
  nand02aa1n03x5               g017(.a(\b[6] ), .b(\a[7] ), .o1(new_n113));
  nona23aa1n12x5               g018(.a(new_n113), .b(new_n111), .c(new_n110), .d(new_n112), .out0(new_n114));
  nor002aa1n03x5               g019(.a(\b[4] ), .b(\a[5] ), .o1(new_n115));
  nand42aa1n02x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  norb02aa1n03x4               g021(.a(new_n116), .b(new_n115), .out0(new_n117));
  nano22aa1n03x7               g022(.a(new_n114), .b(new_n109), .c(new_n117), .out0(new_n118));
  oa0012aa1n02x5               g023(.a(new_n111), .b(new_n112), .c(new_n110), .o(new_n119));
  oai012aa1n02x5               g024(.a(new_n108), .b(new_n115), .c(new_n107), .o1(new_n120));
  oabi12aa1n06x5               g025(.a(new_n119), .b(new_n120), .c(new_n114), .out0(new_n121));
  tech160nm_fixorc02aa1n03p5x5 g026(.a(\a[9] ), .b(\b[8] ), .out0(new_n122));
  aoai13aa1n06x5               g027(.a(new_n122), .b(new_n121), .c(new_n106), .d(new_n118), .o1(new_n123));
  nor002aa1d32x5               g028(.a(\b[9] ), .b(\a[10] ), .o1(new_n124));
  nand42aa1n08x5               g029(.a(\b[9] ), .b(\a[10] ), .o1(new_n125));
  norb02aa1n06x5               g030(.a(new_n125), .b(new_n124), .out0(new_n126));
  xnbna2aa1n03x5               g031(.a(new_n126), .b(new_n123), .c(new_n99), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(new_n124), .o1(new_n128));
  inv000aa1d42x5               g033(.a(new_n126), .o1(new_n129));
  aoai13aa1n04x5               g034(.a(new_n128), .b(new_n129), .c(new_n123), .d(new_n99), .o1(new_n130));
  xorb03aa1n02x5               g035(.a(new_n130), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor022aa1n08x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nanp02aa1n04x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nor022aa1n06x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  nanp02aa1n04x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n135), .b(new_n134), .out0(new_n136));
  aoi112aa1n02x5               g041(.a(new_n132), .b(new_n136), .c(new_n130), .d(new_n133), .o1(new_n137));
  aoai13aa1n02x5               g042(.a(new_n136), .b(new_n132), .c(new_n130), .d(new_n133), .o1(new_n138));
  norb02aa1n02x5               g043(.a(new_n138), .b(new_n137), .out0(\s[12] ));
  nona23aa1n09x5               g044(.a(new_n135), .b(new_n133), .c(new_n132), .d(new_n134), .out0(new_n140));
  nano22aa1n03x7               g045(.a(new_n140), .b(new_n122), .c(new_n126), .out0(new_n141));
  aoai13aa1n06x5               g046(.a(new_n141), .b(new_n121), .c(new_n106), .d(new_n118), .o1(new_n142));
  nano23aa1n03x7               g047(.a(new_n132), .b(new_n134), .c(new_n135), .d(new_n133), .out0(new_n143));
  oai012aa1n02x7               g048(.a(new_n135), .b(new_n134), .c(new_n132), .o1(new_n144));
  aoai13aa1n12x5               g049(.a(new_n125), .b(new_n124), .c(new_n97), .d(new_n98), .o1(new_n145));
  inv000aa1n02x5               g050(.a(new_n145), .o1(new_n146));
  aobi12aa1n06x5               g051(.a(new_n144), .b(new_n143), .c(new_n146), .out0(new_n147));
  nor002aa1d24x5               g052(.a(\b[12] ), .b(\a[13] ), .o1(new_n148));
  nanp02aa1n04x5               g053(.a(\b[12] ), .b(\a[13] ), .o1(new_n149));
  norb02aa1n02x5               g054(.a(new_n149), .b(new_n148), .out0(new_n150));
  xnbna2aa1n03x5               g055(.a(new_n150), .b(new_n142), .c(new_n147), .out0(\s[13] ));
  inv000aa1d42x5               g056(.a(new_n148), .o1(new_n152));
  nanp02aa1n02x5               g057(.a(\b[3] ), .b(\a[4] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(new_n104), .b(new_n105), .o1(new_n154));
  nanp02aa1n02x5               g059(.a(new_n154), .b(new_n153), .o1(new_n155));
  nano23aa1n09x5               g060(.a(new_n110), .b(new_n112), .c(new_n113), .d(new_n111), .out0(new_n156));
  nanp03aa1n02x5               g061(.a(new_n156), .b(new_n109), .c(new_n117), .o1(new_n157));
  aoib12aa1n12x5               g062(.a(new_n119), .b(new_n156), .c(new_n120), .out0(new_n158));
  oai012aa1n06x5               g063(.a(new_n158), .b(new_n155), .c(new_n157), .o1(new_n159));
  tech160nm_fioai012aa1n05x5   g064(.a(new_n144), .b(new_n140), .c(new_n145), .o1(new_n160));
  aoai13aa1n02x5               g065(.a(new_n150), .b(new_n160), .c(new_n159), .d(new_n141), .o1(new_n161));
  nor042aa1n04x5               g066(.a(\b[13] ), .b(\a[14] ), .o1(new_n162));
  nanp02aa1n04x5               g067(.a(\b[13] ), .b(\a[14] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  xnbna2aa1n03x5               g069(.a(new_n164), .b(new_n161), .c(new_n152), .out0(\s[14] ));
  nona23aa1n09x5               g070(.a(new_n163), .b(new_n149), .c(new_n148), .d(new_n162), .out0(new_n166));
  oaoi03aa1n02x5               g071(.a(\a[14] ), .b(\b[13] ), .c(new_n152), .o1(new_n167));
  inv000aa1d42x5               g072(.a(new_n167), .o1(new_n168));
  aoai13aa1n04x5               g073(.a(new_n168), .b(new_n166), .c(new_n142), .d(new_n147), .o1(new_n169));
  xorb03aa1n02x5               g074(.a(new_n169), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g075(.a(\b[14] ), .b(\a[15] ), .o1(new_n171));
  nanp02aa1n04x5               g076(.a(\b[14] ), .b(\a[15] ), .o1(new_n172));
  nor042aa1n03x5               g077(.a(\b[15] ), .b(\a[16] ), .o1(new_n173));
  nand02aa1d20x5               g078(.a(\b[15] ), .b(\a[16] ), .o1(new_n174));
  norb02aa1n02x7               g079(.a(new_n174), .b(new_n173), .out0(new_n175));
  aoi112aa1n02x5               g080(.a(new_n171), .b(new_n175), .c(new_n169), .d(new_n172), .o1(new_n176));
  aoai13aa1n02x5               g081(.a(new_n175), .b(new_n171), .c(new_n169), .d(new_n172), .o1(new_n177));
  norb02aa1n02x5               g082(.a(new_n177), .b(new_n176), .out0(\s[16] ));
  nand02aa1d04x5               g083(.a(new_n106), .b(new_n118), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n172), .b(new_n171), .out0(new_n180));
  nano22aa1n03x7               g085(.a(new_n166), .b(new_n180), .c(new_n175), .out0(new_n181));
  nanp02aa1n02x5               g086(.a(new_n141), .b(new_n181), .o1(new_n182));
  oai112aa1n02x5               g087(.a(new_n163), .b(new_n172), .c(new_n162), .d(new_n148), .o1(new_n183));
  nona22aa1n03x5               g088(.a(new_n183), .b(new_n173), .c(new_n171), .out0(new_n184));
  aoi022aa1d18x5               g089(.a(new_n160), .b(new_n181), .c(new_n174), .d(new_n184), .o1(new_n185));
  aoai13aa1n12x5               g090(.a(new_n185), .b(new_n182), .c(new_n179), .d(new_n158), .o1(new_n186));
  xorb03aa1n02x5               g091(.a(new_n186), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  nano23aa1n03x5               g092(.a(new_n148), .b(new_n162), .c(new_n163), .d(new_n149), .out0(new_n188));
  nanp03aa1n02x5               g093(.a(new_n188), .b(new_n180), .c(new_n175), .o1(new_n189));
  nano32aa1n03x7               g094(.a(new_n189), .b(new_n143), .c(new_n126), .d(new_n122), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n121), .c(new_n106), .d(new_n118), .o1(new_n191));
  nor042aa1n06x5               g096(.a(\b[16] ), .b(\a[17] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(new_n192), .o1(new_n193));
  tech160nm_fixnrc02aa1n04x5   g098(.a(\b[16] ), .b(\a[17] ), .out0(new_n194));
  aoai13aa1n03x5               g099(.a(new_n193), .b(new_n194), .c(new_n191), .d(new_n185), .o1(new_n195));
  xorb03aa1n02x5               g100(.a(new_n195), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  xnrc02aa1n02x5               g101(.a(\b[17] ), .b(\a[18] ), .out0(new_n197));
  nor042aa1n06x5               g102(.a(new_n197), .b(new_n194), .o1(new_n198));
  inv000aa1d42x5               g103(.a(new_n198), .o1(new_n199));
  oaoi03aa1n12x5               g104(.a(\a[18] ), .b(\b[17] ), .c(new_n193), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n06x5               g106(.a(new_n201), .b(new_n199), .c(new_n191), .d(new_n185), .o1(new_n202));
  xorb03aa1n02x5               g107(.a(new_n202), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g108(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n12x5               g109(.a(\b[18] ), .b(\a[19] ), .o1(new_n205));
  nanp02aa1n04x5               g110(.a(\b[18] ), .b(\a[19] ), .o1(new_n206));
  tech160nm_fixnrc02aa1n04x5   g111(.a(\b[19] ), .b(\a[20] ), .out0(new_n207));
  inv000aa1d42x5               g112(.a(new_n207), .o1(new_n208));
  aoi112aa1n02x5               g113(.a(new_n205), .b(new_n208), .c(new_n202), .d(new_n206), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n205), .o1(new_n210));
  nanb02aa1n18x5               g115(.a(new_n205), .b(new_n206), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  aoai13aa1n02x7               g117(.a(new_n212), .b(new_n200), .c(new_n186), .d(new_n198), .o1(new_n213));
  aoi012aa1n03x5               g118(.a(new_n207), .b(new_n213), .c(new_n210), .o1(new_n214));
  norp02aa1n03x5               g119(.a(new_n214), .b(new_n209), .o1(\s[20] ));
  nona22aa1n09x5               g120(.a(new_n198), .b(new_n211), .c(new_n207), .out0(new_n216));
  nanp02aa1n02x5               g121(.a(\b[17] ), .b(\a[18] ), .o1(new_n217));
  oai022aa1n02x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  nanp03aa1n02x5               g123(.a(new_n218), .b(new_n217), .c(new_n206), .o1(new_n219));
  oab012aa1n02x4               g124(.a(new_n205), .b(\a[20] ), .c(\b[19] ), .out0(new_n220));
  aoi022aa1n02x5               g125(.a(new_n219), .b(new_n220), .c(\b[19] ), .d(\a[20] ), .o1(new_n221));
  inv000aa1n02x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n216), .c(new_n191), .d(new_n185), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1d32x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  nand42aa1n04x5               g130(.a(\b[20] ), .b(\a[21] ), .o1(new_n226));
  norb02aa1n02x5               g131(.a(new_n226), .b(new_n225), .out0(new_n227));
  nor022aa1n16x5               g132(.a(\b[21] ), .b(\a[22] ), .o1(new_n228));
  nanp02aa1n04x5               g133(.a(\b[21] ), .b(\a[22] ), .o1(new_n229));
  norb02aa1n02x5               g134(.a(new_n229), .b(new_n228), .out0(new_n230));
  aoi112aa1n03x4               g135(.a(new_n225), .b(new_n230), .c(new_n223), .d(new_n227), .o1(new_n231));
  inv000aa1n03x5               g136(.a(new_n225), .o1(new_n232));
  inv000aa1d42x5               g137(.a(new_n216), .o1(new_n233));
  aoai13aa1n03x5               g138(.a(new_n227), .b(new_n221), .c(new_n186), .d(new_n233), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n230), .o1(new_n235));
  tech160nm_fiaoi012aa1n02p5x5 g140(.a(new_n235), .b(new_n234), .c(new_n232), .o1(new_n236));
  nor002aa1n02x5               g141(.a(new_n236), .b(new_n231), .o1(\s[22] ));
  nona23aa1d24x5               g142(.a(new_n229), .b(new_n226), .c(new_n225), .d(new_n228), .out0(new_n238));
  nona23aa1d18x5               g143(.a(new_n198), .b(new_n208), .c(new_n238), .d(new_n211), .out0(new_n239));
  and002aa1n02x5               g144(.a(\b[19] ), .b(\a[20] ), .o(new_n240));
  aoi112aa1n02x5               g145(.a(new_n238), .b(new_n240), .c(new_n219), .d(new_n220), .o1(new_n241));
  oaoi03aa1n02x5               g146(.a(\a[22] ), .b(\b[21] ), .c(new_n232), .o1(new_n242));
  norp02aa1n02x5               g147(.a(new_n241), .b(new_n242), .o1(new_n243));
  aoai13aa1n06x5               g148(.a(new_n243), .b(new_n239), .c(new_n191), .d(new_n185), .o1(new_n244));
  xorb03aa1n02x5               g149(.a(new_n244), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n12x5               g150(.a(\b[22] ), .b(\a[23] ), .o1(new_n246));
  nanp02aa1n02x5               g151(.a(\b[22] ), .b(\a[23] ), .o1(new_n247));
  norb02aa1n06x4               g152(.a(new_n247), .b(new_n246), .out0(new_n248));
  xorc02aa1n02x5               g153(.a(\a[24] ), .b(\b[23] ), .out0(new_n249));
  aoi112aa1n02x5               g154(.a(new_n246), .b(new_n249), .c(new_n244), .d(new_n248), .o1(new_n250));
  inv000aa1d42x5               g155(.a(new_n246), .o1(new_n251));
  inv000aa1d42x5               g156(.a(new_n239), .o1(new_n252));
  inv000aa1n02x5               g157(.a(new_n243), .o1(new_n253));
  aoai13aa1n03x5               g158(.a(new_n248), .b(new_n253), .c(new_n186), .d(new_n252), .o1(new_n254));
  xnrc02aa1n02x5               g159(.a(\b[23] ), .b(\a[24] ), .out0(new_n255));
  aoi012aa1n02x7               g160(.a(new_n255), .b(new_n254), .c(new_n251), .o1(new_n256));
  nor002aa1n02x5               g161(.a(new_n256), .b(new_n250), .o1(\s[24] ));
  inv000aa1d42x5               g162(.a(new_n238), .o1(new_n258));
  nano22aa1n03x7               g163(.a(new_n255), .b(new_n251), .c(new_n247), .out0(new_n259));
  nano22aa1n03x7               g164(.a(new_n216), .b(new_n258), .c(new_n259), .out0(new_n260));
  inv000aa1n02x5               g165(.a(new_n260), .o1(new_n261));
  nanp02aa1n02x5               g166(.a(new_n219), .b(new_n220), .o1(new_n262));
  nona23aa1n09x5               g167(.a(new_n262), .b(new_n259), .c(new_n238), .d(new_n240), .out0(new_n263));
  oaoi03aa1n02x5               g168(.a(\a[24] ), .b(\b[23] ), .c(new_n251), .o1(new_n264));
  aoi013aa1n06x4               g169(.a(new_n264), .b(new_n242), .c(new_n249), .d(new_n248), .o1(new_n265));
  nanp02aa1n02x5               g170(.a(new_n263), .b(new_n265), .o1(new_n266));
  inv000aa1n02x5               g171(.a(new_n266), .o1(new_n267));
  aoai13aa1n06x5               g172(.a(new_n267), .b(new_n261), .c(new_n191), .d(new_n185), .o1(new_n268));
  xorb03aa1n02x5               g173(.a(new_n268), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  nor042aa1n03x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  xorc02aa1n02x5               g175(.a(\a[25] ), .b(\b[24] ), .out0(new_n271));
  xorc02aa1n12x5               g176(.a(\a[26] ), .b(\b[25] ), .out0(new_n272));
  aoi112aa1n02x5               g177(.a(new_n270), .b(new_n272), .c(new_n268), .d(new_n271), .o1(new_n273));
  inv000aa1d42x5               g178(.a(new_n270), .o1(new_n274));
  aoai13aa1n03x5               g179(.a(new_n271), .b(new_n266), .c(new_n186), .d(new_n260), .o1(new_n275));
  inv000aa1d42x5               g180(.a(new_n272), .o1(new_n276));
  aoi012aa1n03x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .o1(new_n277));
  nor002aa1n02x5               g182(.a(new_n277), .b(new_n273), .o1(\s[26] ));
  nanp02aa1n02x5               g183(.a(new_n184), .b(new_n174), .o1(new_n279));
  oai012aa1n02x5               g184(.a(new_n279), .b(new_n147), .c(new_n189), .o1(new_n280));
  and002aa1n02x5               g185(.a(new_n272), .b(new_n271), .o(new_n281));
  nano22aa1d15x5               g186(.a(new_n239), .b(new_n281), .c(new_n259), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n280), .c(new_n159), .d(new_n190), .o1(new_n283));
  inv040aa1n02x5               g188(.a(new_n281), .o1(new_n284));
  oao003aa1n02x5               g189(.a(\a[26] ), .b(\b[25] ), .c(new_n274), .carry(new_n285));
  aoai13aa1n12x5               g190(.a(new_n285), .b(new_n284), .c(new_n263), .d(new_n265), .o1(new_n286));
  inv040aa1n06x5               g191(.a(new_n286), .o1(new_n287));
  nor002aa1n12x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  nanp02aa1n02x5               g193(.a(\b[26] ), .b(\a[27] ), .o1(new_n289));
  nanb02aa1n06x5               g194(.a(new_n288), .b(new_n289), .out0(new_n290));
  xobna2aa1n03x5               g195(.a(new_n290), .b(new_n283), .c(new_n287), .out0(\s[27] ));
  inv000aa1d42x5               g196(.a(new_n288), .o1(new_n292));
  aoai13aa1n03x5               g197(.a(new_n289), .b(new_n286), .c(new_n186), .d(new_n282), .o1(new_n293));
  xnrc02aa1n02x5               g198(.a(\b[27] ), .b(\a[28] ), .out0(new_n294));
  aoi012aa1n03x5               g199(.a(new_n294), .b(new_n293), .c(new_n292), .o1(new_n295));
  aoi022aa1n02x7               g200(.a(new_n283), .b(new_n287), .c(\b[26] ), .d(\a[27] ), .o1(new_n296));
  nano22aa1n03x5               g201(.a(new_n296), .b(new_n292), .c(new_n294), .out0(new_n297));
  norp02aa1n03x5               g202(.a(new_n295), .b(new_n297), .o1(\s[28] ));
  nor042aa1n04x5               g203(.a(new_n294), .b(new_n290), .o1(new_n299));
  aoai13aa1n03x5               g204(.a(new_n299), .b(new_n286), .c(new_n186), .d(new_n282), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .carry(new_n301));
  xnrc02aa1n12x5               g206(.a(\b[28] ), .b(\a[29] ), .out0(new_n302));
  aoi012aa1n03x5               g207(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n299), .o1(new_n304));
  tech160nm_fiaoi012aa1n02p5x5 g209(.a(new_n304), .b(new_n283), .c(new_n287), .o1(new_n305));
  nano22aa1n03x5               g210(.a(new_n305), .b(new_n301), .c(new_n302), .out0(new_n306));
  norp02aa1n03x5               g211(.a(new_n303), .b(new_n306), .o1(\s[29] ));
  xorb03aa1n02x5               g212(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norp03aa1n02x5               g213(.a(new_n302), .b(new_n294), .c(new_n290), .o1(new_n309));
  aoai13aa1n03x5               g214(.a(new_n309), .b(new_n286), .c(new_n186), .d(new_n282), .o1(new_n310));
  oao003aa1n02x5               g215(.a(\a[29] ), .b(\b[28] ), .c(new_n301), .carry(new_n311));
  xnrc02aa1n02x5               g216(.a(\b[29] ), .b(\a[30] ), .out0(new_n312));
  tech160nm_fiaoi012aa1n02p5x5 g217(.a(new_n312), .b(new_n310), .c(new_n311), .o1(new_n313));
  inv020aa1n02x5               g218(.a(new_n309), .o1(new_n314));
  tech160nm_fiaoi012aa1n02p5x5 g219(.a(new_n314), .b(new_n283), .c(new_n287), .o1(new_n315));
  nano22aa1n03x5               g220(.a(new_n315), .b(new_n311), .c(new_n312), .out0(new_n316));
  norp02aa1n03x5               g221(.a(new_n313), .b(new_n316), .o1(\s[30] ));
  xnrc02aa1n02x5               g222(.a(\b[30] ), .b(\a[31] ), .out0(new_n318));
  norb03aa1n03x5               g223(.a(new_n299), .b(new_n312), .c(new_n302), .out0(new_n319));
  aoai13aa1n06x5               g224(.a(new_n319), .b(new_n286), .c(new_n186), .d(new_n282), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n321));
  tech160nm_fiaoi012aa1n05x5   g226(.a(new_n318), .b(new_n320), .c(new_n321), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n319), .o1(new_n323));
  tech160nm_fiaoi012aa1n03p5x5 g228(.a(new_n323), .b(new_n283), .c(new_n287), .o1(new_n324));
  nano22aa1n03x5               g229(.a(new_n324), .b(new_n318), .c(new_n321), .out0(new_n325));
  norp02aa1n03x5               g230(.a(new_n322), .b(new_n325), .o1(\s[31] ));
  oai012aa1n02x5               g231(.a(new_n101), .b(new_n102), .c(new_n100), .o1(new_n327));
  xnrb03aa1n02x5               g232(.a(new_n327), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g233(.a(\a[3] ), .b(\b[2] ), .c(new_n327), .o1(new_n329));
  xorb03aa1n02x5               g234(.a(new_n329), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g235(.a(new_n106), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi13aa1n02x5               g236(.a(new_n109), .b(new_n116), .c(new_n106), .d(new_n115), .o1(new_n332));
  oai112aa1n02x5               g237(.a(new_n116), .b(new_n109), .c(new_n106), .d(new_n115), .o1(new_n333));
  norb02aa1n02x5               g238(.a(new_n333), .b(new_n332), .out0(\s[6] ));
  norb02aa1n02x5               g239(.a(new_n333), .b(new_n107), .out0(new_n335));
  xnrb03aa1n02x5               g240(.a(new_n335), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g241(.a(\a[7] ), .b(\b[6] ), .c(new_n335), .o1(new_n337));
  xorb03aa1n02x5               g242(.a(new_n337), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g243(.a(new_n122), .b(new_n179), .c(new_n158), .out0(\s[9] ));
endmodule


