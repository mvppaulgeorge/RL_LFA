// Benchmark "adder" written by ABC on Wed Jul 17 19:24:32 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n162, new_n163, new_n164, new_n165, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n176,
    new_n177, new_n178, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n186, new_n187, new_n188, new_n189, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n366,
    new_n367, new_n369, new_n370, new_n371, new_n372, new_n374, new_n376,
    new_n377, new_n378, new_n380;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  orn002aa1n24x5               g001(.a(\a[2] ), .b(\b[1] ), .o(new_n97));
  nand42aa1n02x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand02aa1n04x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  nand02aa1n04x5               g004(.a(new_n99), .b(new_n98), .o1(new_n100));
  nor002aa1d32x5               g005(.a(\b[2] ), .b(\a[3] ), .o1(new_n101));
  nand02aa1d06x5               g006(.a(\b[2] ), .b(\a[3] ), .o1(new_n102));
  nanb02aa1n02x5               g007(.a(new_n101), .b(new_n102), .out0(new_n103));
  nand42aa1n16x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  nor002aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  norb03aa1n03x5               g010(.a(new_n104), .b(new_n101), .c(new_n105), .out0(new_n106));
  aoai13aa1n04x5               g011(.a(new_n106), .b(new_n103), .c(new_n97), .d(new_n100), .o1(new_n107));
  nor002aa1n12x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  nor002aa1d32x5               g013(.a(\b[4] ), .b(\a[5] ), .o1(new_n109));
  nor002aa1n03x5               g014(.a(\b[5] ), .b(\a[6] ), .o1(new_n110));
  nor043aa1d12x5               g015(.a(new_n110), .b(new_n109), .c(new_n108), .o1(new_n111));
  oai012aa1n12x5               g016(.a(new_n104), .b(\b[7] ), .c(\a[8] ), .o1(new_n112));
  nanp02aa1n24x5               g017(.a(\b[5] ), .b(\a[6] ), .o1(new_n113));
  nand02aa1n04x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand02aa1n02x5               g019(.a(new_n114), .b(new_n113), .o1(new_n115));
  aoi022aa1n09x5               g020(.a(\b[7] ), .b(\a[8] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n116));
  norb03aa1n03x5               g021(.a(new_n116), .b(new_n115), .c(new_n112), .out0(new_n117));
  inv000aa1d42x5               g022(.a(new_n109), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[7] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[6] ), .o1(new_n120));
  nor042aa1n04x5               g025(.a(\b[7] ), .b(\a[8] ), .o1(new_n121));
  nand02aa1n06x5               g026(.a(\b[7] ), .b(\a[8] ), .o1(new_n122));
  aoai13aa1n04x5               g027(.a(new_n122), .b(new_n121), .c(new_n119), .d(new_n120), .o1(new_n123));
  norb02aa1n06x4               g028(.a(new_n113), .b(new_n110), .out0(new_n124));
  aoi022aa1n02x7               g029(.a(\b[6] ), .b(\a[7] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n125));
  nona23aa1n02x4               g030(.a(new_n125), .b(new_n122), .c(new_n121), .d(new_n108), .out0(new_n126));
  aoai13aa1n03x5               g031(.a(new_n123), .b(new_n126), .c(new_n124), .d(new_n118), .o1(new_n127));
  aoi013aa1n06x4               g032(.a(new_n127), .b(new_n107), .c(new_n111), .d(new_n117), .o1(new_n128));
  tech160nm_fioaoi03aa1n02p5x5 g033(.a(\a[9] ), .b(\b[8] ), .c(new_n128), .o1(new_n129));
  nor042aa1n06x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  and002aa1n12x5               g035(.a(\b[9] ), .b(\a[10] ), .o(new_n131));
  nor042aa1n04x5               g036(.a(new_n131), .b(new_n130), .o1(new_n132));
  nor042aa1n06x5               g037(.a(\b[8] ), .b(\a[9] ), .o1(new_n133));
  nand02aa1n08x5               g038(.a(new_n100), .b(new_n97), .o1(new_n134));
  norb02aa1n06x5               g039(.a(new_n102), .b(new_n101), .out0(new_n135));
  nona22aa1n09x5               g040(.a(new_n104), .b(new_n105), .c(new_n101), .out0(new_n136));
  aoi012aa1d18x5               g041(.a(new_n136), .b(new_n134), .c(new_n135), .o1(new_n137));
  nona23aa1d18x5               g042(.a(new_n111), .b(new_n116), .c(new_n115), .d(new_n112), .out0(new_n138));
  inv000aa1n02x5               g043(.a(new_n123), .o1(new_n139));
  inv040aa1n12x5               g044(.a(\a[6] ), .o1(new_n140));
  inv000aa1d48x5               g045(.a(\b[5] ), .o1(new_n141));
  nand42aa1n06x5               g046(.a(new_n141), .b(new_n140), .o1(new_n142));
  oai112aa1n06x5               g047(.a(new_n142), .b(new_n113), .c(\b[4] ), .d(\a[5] ), .o1(new_n143));
  nano22aa1n03x7               g048(.a(new_n108), .b(new_n113), .c(new_n114), .out0(new_n144));
  norb02aa1n06x5               g049(.a(new_n122), .b(new_n121), .out0(new_n145));
  aoi013aa1n06x4               g050(.a(new_n139), .b(new_n144), .c(new_n143), .d(new_n145), .o1(new_n146));
  oai012aa1d24x5               g051(.a(new_n146), .b(new_n137), .c(new_n138), .o1(new_n147));
  xorc02aa1n12x5               g052(.a(\a[9] ), .b(\b[8] ), .out0(new_n148));
  aoi112aa1n02x5               g053(.a(new_n132), .b(new_n133), .c(new_n147), .d(new_n148), .o1(new_n149));
  aoi012aa1n02x5               g054(.a(new_n149), .b(new_n129), .c(new_n132), .o1(\s[10] ));
  aoai13aa1n03x5               g055(.a(new_n132), .b(new_n133), .c(new_n147), .d(new_n148), .o1(new_n151));
  oabi12aa1n18x5               g056(.a(new_n131), .b(new_n133), .c(new_n130), .out0(new_n152));
  nor002aa1d32x5               g057(.a(\b[10] ), .b(\a[11] ), .o1(new_n153));
  nand02aa1d28x5               g058(.a(\b[10] ), .b(\a[11] ), .o1(new_n154));
  norb02aa1n09x5               g059(.a(new_n154), .b(new_n153), .out0(new_n155));
  xnbna2aa1n03x5               g060(.a(new_n155), .b(new_n151), .c(new_n152), .out0(\s[11] ));
  oab012aa1n06x5               g061(.a(new_n131), .b(new_n133), .c(new_n130), .out0(new_n157));
  aoai13aa1n02x5               g062(.a(new_n155), .b(new_n157), .c(new_n129), .d(new_n132), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n153), .o1(new_n159));
  inv000aa1d42x5               g064(.a(new_n155), .o1(new_n160));
  aoai13aa1n02x7               g065(.a(new_n159), .b(new_n160), .c(new_n151), .d(new_n152), .o1(new_n161));
  nor002aa1n16x5               g066(.a(\b[11] ), .b(\a[12] ), .o1(new_n162));
  nand02aa1d28x5               g067(.a(\b[11] ), .b(\a[12] ), .o1(new_n163));
  norb02aa1n02x5               g068(.a(new_n163), .b(new_n162), .out0(new_n164));
  aoib12aa1n02x5               g069(.a(new_n153), .b(new_n163), .c(new_n162), .out0(new_n165));
  aoi022aa1n02x7               g070(.a(new_n161), .b(new_n164), .c(new_n158), .d(new_n165), .o1(\s[12] ));
  nano23aa1n09x5               g071(.a(new_n153), .b(new_n162), .c(new_n163), .d(new_n154), .out0(new_n167));
  nand23aa1n03x5               g072(.a(new_n167), .b(new_n148), .c(new_n132), .o1(new_n168));
  nona23aa1d16x5               g073(.a(new_n163), .b(new_n154), .c(new_n153), .d(new_n162), .out0(new_n169));
  aoi012aa1n09x5               g074(.a(new_n162), .b(new_n153), .c(new_n163), .o1(new_n170));
  oai012aa1d24x5               g075(.a(new_n170), .b(new_n169), .c(new_n152), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  oaih12aa1n02x5               g077(.a(new_n172), .b(new_n128), .c(new_n168), .o1(new_n173));
  nor002aa1d32x5               g078(.a(\b[12] ), .b(\a[13] ), .o1(new_n174));
  nand02aa1d16x5               g079(.a(\b[12] ), .b(\a[13] ), .o1(new_n175));
  norb02aa1n03x5               g080(.a(new_n175), .b(new_n174), .out0(new_n176));
  nano22aa1n03x7               g081(.a(new_n169), .b(new_n148), .c(new_n132), .out0(new_n177));
  aoi112aa1n02x5               g082(.a(new_n176), .b(new_n171), .c(new_n147), .d(new_n177), .o1(new_n178));
  aoi012aa1n02x5               g083(.a(new_n178), .b(new_n173), .c(new_n176), .o1(\s[13] ));
  inv000aa1d42x5               g084(.a(new_n174), .o1(new_n180));
  aoai13aa1n03x5               g085(.a(new_n176), .b(new_n171), .c(new_n147), .d(new_n177), .o1(new_n181));
  nor022aa1n16x5               g086(.a(\b[13] ), .b(\a[14] ), .o1(new_n182));
  nand02aa1d16x5               g087(.a(\b[13] ), .b(\a[14] ), .o1(new_n183));
  norb02aa1n03x5               g088(.a(new_n183), .b(new_n182), .out0(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n184), .b(new_n181), .c(new_n180), .out0(\s[14] ));
  nano23aa1n06x5               g090(.a(new_n174), .b(new_n182), .c(new_n183), .d(new_n175), .out0(new_n186));
  aoai13aa1n06x5               g091(.a(new_n186), .b(new_n171), .c(new_n147), .d(new_n177), .o1(new_n187));
  oai012aa1n03x5               g092(.a(new_n183), .b(new_n182), .c(new_n174), .o1(new_n188));
  xorc02aa1n12x5               g093(.a(\a[15] ), .b(\b[14] ), .out0(new_n189));
  xnbna2aa1n03x5               g094(.a(new_n189), .b(new_n187), .c(new_n188), .out0(\s[15] ));
  inv000aa1d42x5               g095(.a(new_n188), .o1(new_n191));
  aoai13aa1n02x5               g096(.a(new_n189), .b(new_n191), .c(new_n173), .d(new_n186), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\a[15] ), .o1(new_n193));
  inv000aa1d42x5               g098(.a(\b[14] ), .o1(new_n194));
  nanp02aa1n06x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  inv040aa1n02x5               g100(.a(new_n189), .o1(new_n196));
  aoai13aa1n03x5               g101(.a(new_n195), .b(new_n196), .c(new_n187), .d(new_n188), .o1(new_n197));
  xorc02aa1n12x5               g102(.a(\a[16] ), .b(\b[15] ), .out0(new_n198));
  inv000aa1d42x5               g103(.a(\b[15] ), .o1(new_n199));
  nanb02aa1n12x5               g104(.a(\a[16] ), .b(new_n199), .out0(new_n200));
  nand42aa1n02x5               g105(.a(\b[15] ), .b(\a[16] ), .o1(new_n201));
  aoi022aa1n02x5               g106(.a(new_n200), .b(new_n201), .c(new_n194), .d(new_n193), .o1(new_n202));
  aoi022aa1n03x5               g107(.a(new_n197), .b(new_n198), .c(new_n192), .d(new_n202), .o1(\s[16] ));
  nand23aa1n04x5               g108(.a(new_n186), .b(new_n189), .c(new_n198), .o1(new_n204));
  nor042aa1n04x5               g109(.a(new_n204), .b(new_n168), .o1(new_n205));
  nanp02aa1n02x5               g110(.a(new_n147), .b(new_n205), .o1(new_n206));
  nano32aa1n03x7               g111(.a(new_n196), .b(new_n198), .c(new_n176), .d(new_n184), .out0(new_n207));
  nand02aa1n02x5               g112(.a(new_n207), .b(new_n177), .o1(new_n208));
  oai112aa1n06x5               g113(.a(new_n200), .b(new_n201), .c(new_n194), .d(new_n193), .o1(new_n209));
  oai112aa1n04x5               g114(.a(new_n183), .b(new_n195), .c(new_n182), .d(new_n174), .o1(new_n210));
  oaoi03aa1n02x5               g115(.a(\a[16] ), .b(\b[15] ), .c(new_n195), .o1(new_n211));
  oabi12aa1n02x5               g116(.a(new_n211), .b(new_n210), .c(new_n209), .out0(new_n212));
  aoi012aa1n12x5               g117(.a(new_n212), .b(new_n207), .c(new_n171), .o1(new_n213));
  oaih12aa1n12x5               g118(.a(new_n213), .b(new_n128), .c(new_n208), .o1(new_n214));
  xorc02aa1n02x5               g119(.a(\a[17] ), .b(\b[16] ), .out0(new_n215));
  aoi112aa1n02x5               g120(.a(new_n212), .b(new_n215), .c(new_n207), .d(new_n171), .o1(new_n216));
  aoi022aa1n02x5               g121(.a(new_n214), .b(new_n215), .c(new_n206), .d(new_n216), .o1(\s[17] ));
  inv000aa1d42x5               g122(.a(\a[17] ), .o1(new_n218));
  nanb02aa1d24x5               g123(.a(\b[16] ), .b(new_n218), .out0(new_n219));
  nanp02aa1n04x5               g124(.a(new_n167), .b(new_n157), .o1(new_n220));
  oab012aa1n06x5               g125(.a(new_n211), .b(new_n210), .c(new_n209), .out0(new_n221));
  aoai13aa1n12x5               g126(.a(new_n221), .b(new_n204), .c(new_n220), .d(new_n170), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n215), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n223));
  xorc02aa1n02x5               g128(.a(\a[18] ), .b(\b[17] ), .out0(new_n224));
  xnbna2aa1n03x5               g129(.a(new_n224), .b(new_n223), .c(new_n219), .out0(\s[18] ));
  inv000aa1d42x5               g130(.a(\a[18] ), .o1(new_n226));
  xroi22aa1d04x5               g131(.a(new_n218), .b(\b[16] ), .c(new_n226), .d(\b[17] ), .out0(new_n227));
  aoai13aa1n06x5               g132(.a(new_n227), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n228));
  oaoi03aa1n12x5               g133(.a(\a[18] ), .b(\b[17] ), .c(new_n219), .o1(new_n229));
  inv000aa1d42x5               g134(.a(new_n229), .o1(new_n230));
  nor002aa1d32x5               g135(.a(\b[18] ), .b(\a[19] ), .o1(new_n231));
  nanp02aa1n06x5               g136(.a(\b[18] ), .b(\a[19] ), .o1(new_n232));
  norb02aa1n09x5               g137(.a(new_n232), .b(new_n231), .out0(new_n233));
  xnbna2aa1n03x5               g138(.a(new_n233), .b(new_n228), .c(new_n230), .out0(\s[19] ));
  xnrc02aa1n02x5               g139(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g140(.a(new_n233), .b(new_n229), .c(new_n214), .d(new_n227), .o1(new_n236));
  inv040aa1n02x5               g141(.a(new_n231), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n233), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n237), .b(new_n238), .c(new_n228), .d(new_n230), .o1(new_n239));
  xorc02aa1n02x5               g144(.a(\a[20] ), .b(\b[19] ), .out0(new_n240));
  inv040aa1d32x5               g145(.a(\a[20] ), .o1(new_n241));
  inv040aa1d28x5               g146(.a(\b[19] ), .o1(new_n242));
  nanp02aa1n06x5               g147(.a(new_n242), .b(new_n241), .o1(new_n243));
  nand22aa1n12x5               g148(.a(\b[19] ), .b(\a[20] ), .o1(new_n244));
  aoi012aa1n02x5               g149(.a(new_n231), .b(new_n243), .c(new_n244), .o1(new_n245));
  aoi022aa1n03x5               g150(.a(new_n239), .b(new_n240), .c(new_n236), .d(new_n245), .o1(\s[20] ));
  nano32aa1n03x7               g151(.a(new_n238), .b(new_n240), .c(new_n215), .d(new_n224), .out0(new_n247));
  aoai13aa1n06x5               g152(.a(new_n247), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n248));
  nanp03aa1n04x5               g153(.a(new_n243), .b(new_n232), .c(new_n244), .o1(new_n249));
  nanp02aa1n03x5               g154(.a(\b[17] ), .b(\a[18] ), .o1(new_n250));
  oai022aa1d24x5               g155(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n251));
  oai112aa1n06x5               g156(.a(new_n251), .b(new_n250), .c(\b[18] ), .d(\a[19] ), .o1(new_n252));
  oaoi03aa1n09x5               g157(.a(new_n241), .b(new_n242), .c(new_n231), .o1(new_n253));
  oai012aa1n12x5               g158(.a(new_n253), .b(new_n252), .c(new_n249), .o1(new_n254));
  inv000aa1d42x5               g159(.a(new_n254), .o1(new_n255));
  nor042aa1d18x5               g160(.a(\b[20] ), .b(\a[21] ), .o1(new_n256));
  nanp02aa1n09x5               g161(.a(\b[20] ), .b(\a[21] ), .o1(new_n257));
  norb02aa1n12x5               g162(.a(new_n257), .b(new_n256), .out0(new_n258));
  xnbna2aa1n03x5               g163(.a(new_n258), .b(new_n248), .c(new_n255), .out0(\s[21] ));
  aoai13aa1n03x5               g164(.a(new_n258), .b(new_n254), .c(new_n214), .d(new_n247), .o1(new_n260));
  inv000aa1d42x5               g165(.a(new_n256), .o1(new_n261));
  inv000aa1d42x5               g166(.a(new_n258), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n261), .b(new_n262), .c(new_n248), .d(new_n255), .o1(new_n263));
  nor002aa1n03x5               g168(.a(\b[21] ), .b(\a[22] ), .o1(new_n264));
  nand42aa1n06x5               g169(.a(\b[21] ), .b(\a[22] ), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n265), .b(new_n264), .out0(new_n266));
  aoib12aa1n02x5               g171(.a(new_n256), .b(new_n265), .c(new_n264), .out0(new_n267));
  aoi022aa1n03x5               g172(.a(new_n263), .b(new_n266), .c(new_n260), .d(new_n267), .o1(\s[22] ));
  inv000aa1n02x5               g173(.a(new_n244), .o1(new_n269));
  nano32aa1n03x7               g174(.a(new_n269), .b(new_n237), .c(new_n243), .d(new_n232), .out0(new_n270));
  nano23aa1n06x5               g175(.a(new_n256), .b(new_n264), .c(new_n265), .d(new_n257), .out0(new_n271));
  and003aa1n02x5               g176(.a(new_n227), .b(new_n271), .c(new_n270), .o(new_n272));
  aoai13aa1n06x5               g177(.a(new_n272), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n273));
  oai022aa1n04x5               g178(.a(\a[21] ), .b(\b[20] ), .c(\b[21] ), .d(\a[22] ), .o1(new_n274));
  aoi022aa1n02x5               g179(.a(new_n254), .b(new_n271), .c(new_n265), .d(new_n274), .o1(new_n275));
  xorc02aa1n12x5               g180(.a(\a[23] ), .b(\b[22] ), .out0(new_n276));
  xnbna2aa1n03x5               g181(.a(new_n276), .b(new_n273), .c(new_n275), .out0(\s[23] ));
  inv040aa1n03x5               g182(.a(new_n275), .o1(new_n278));
  aoai13aa1n03x5               g183(.a(new_n276), .b(new_n278), .c(new_n214), .d(new_n272), .o1(new_n279));
  inv000aa1d42x5               g184(.a(\a[23] ), .o1(new_n280));
  inv030aa1n04x5               g185(.a(\b[22] ), .o1(new_n281));
  nand02aa1n03x5               g186(.a(new_n281), .b(new_n280), .o1(new_n282));
  inv000aa1n02x5               g187(.a(new_n276), .o1(new_n283));
  aoai13aa1n02x5               g188(.a(new_n282), .b(new_n283), .c(new_n273), .d(new_n275), .o1(new_n284));
  xorc02aa1n03x5               g189(.a(\a[24] ), .b(\b[23] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(\b[23] ), .o1(new_n286));
  nanb02aa1n12x5               g191(.a(\a[24] ), .b(new_n286), .out0(new_n287));
  nanp02aa1n02x5               g192(.a(\b[23] ), .b(\a[24] ), .o1(new_n288));
  aoi022aa1n02x5               g193(.a(new_n287), .b(new_n288), .c(new_n281), .d(new_n280), .o1(new_n289));
  aoi022aa1n03x5               g194(.a(new_n284), .b(new_n285), .c(new_n279), .d(new_n289), .o1(\s[24] ));
  nand23aa1n04x5               g195(.a(new_n271), .b(new_n276), .c(new_n285), .o1(new_n291));
  nano22aa1n02x5               g196(.a(new_n291), .b(new_n227), .c(new_n270), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n293));
  oai012aa1n02x5               g198(.a(new_n232), .b(\b[19] ), .c(\a[20] ), .o1(new_n294));
  nona32aa1n06x5               g199(.a(new_n229), .b(new_n294), .c(new_n269), .d(new_n231), .out0(new_n295));
  oai112aa1n02x5               g200(.a(new_n287), .b(new_n288), .c(new_n281), .d(new_n280), .o1(new_n296));
  nanp03aa1n02x5               g201(.a(new_n274), .b(new_n282), .c(new_n265), .o1(new_n297));
  oaoi03aa1n02x5               g202(.a(\a[24] ), .b(\b[23] ), .c(new_n282), .o1(new_n298));
  oab012aa1n09x5               g203(.a(new_n298), .b(new_n297), .c(new_n296), .out0(new_n299));
  aoai13aa1n04x5               g204(.a(new_n299), .b(new_n291), .c(new_n295), .d(new_n253), .o1(new_n300));
  inv000aa1n02x5               g205(.a(new_n300), .o1(new_n301));
  nanp02aa1n02x5               g206(.a(new_n293), .b(new_n301), .o1(new_n302));
  xorc02aa1n02x5               g207(.a(\a[25] ), .b(\b[24] ), .out0(new_n303));
  nano32aa1n03x7               g208(.a(new_n283), .b(new_n285), .c(new_n258), .d(new_n266), .out0(new_n304));
  nand22aa1n03x5               g209(.a(new_n304), .b(new_n254), .o1(new_n305));
  inv000aa1n02x5               g210(.a(new_n303), .o1(new_n306));
  and003aa1n02x5               g211(.a(new_n305), .b(new_n306), .c(new_n299), .o(new_n307));
  aoi022aa1n02x5               g212(.a(new_n302), .b(new_n303), .c(new_n293), .d(new_n307), .o1(\s[25] ));
  aoai13aa1n03x5               g213(.a(new_n303), .b(new_n300), .c(new_n214), .d(new_n292), .o1(new_n309));
  nor042aa1d18x5               g214(.a(\b[24] ), .b(\a[25] ), .o1(new_n310));
  inv040aa1n04x5               g215(.a(new_n310), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n306), .c(new_n293), .d(new_n301), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[26] ), .b(\b[25] ), .out0(new_n313));
  norp02aa1n02x5               g218(.a(new_n313), .b(new_n310), .o1(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[26] ));
  nand42aa1n03x5               g220(.a(\b[24] ), .b(\a[25] ), .o1(new_n316));
  xnrc02aa1n12x5               g221(.a(\b[25] ), .b(\a[26] ), .out0(new_n317));
  nano22aa1d15x5               g222(.a(new_n317), .b(new_n311), .c(new_n316), .out0(new_n318));
  nano32aa1n03x7               g223(.a(new_n291), .b(new_n227), .c(new_n318), .d(new_n270), .out0(new_n319));
  aoai13aa1n06x5               g224(.a(new_n319), .b(new_n222), .c(new_n147), .d(new_n205), .o1(new_n320));
  oao003aa1n02x5               g225(.a(\a[26] ), .b(\b[25] ), .c(new_n311), .carry(new_n321));
  inv000aa1d42x5               g226(.a(new_n321), .o1(new_n322));
  tech160nm_fiaoi012aa1n05x5   g227(.a(new_n322), .b(new_n300), .c(new_n318), .o1(new_n323));
  nanp02aa1n03x5               g228(.a(new_n320), .b(new_n323), .o1(new_n324));
  xorc02aa1n12x5               g229(.a(\a[27] ), .b(\b[26] ), .out0(new_n325));
  aoi112aa1n03x4               g230(.a(new_n325), .b(new_n322), .c(new_n300), .d(new_n318), .o1(new_n326));
  aoi022aa1n02x7               g231(.a(new_n324), .b(new_n325), .c(new_n326), .d(new_n320), .o1(\s[27] ));
  inv000aa1d42x5               g232(.a(new_n318), .o1(new_n328));
  aoai13aa1n04x5               g233(.a(new_n321), .b(new_n328), .c(new_n305), .d(new_n299), .o1(new_n329));
  aoai13aa1n03x5               g234(.a(new_n325), .b(new_n329), .c(new_n214), .d(new_n319), .o1(new_n330));
  nor042aa1n03x5               g235(.a(\b[26] ), .b(\a[27] ), .o1(new_n331));
  inv000aa1n03x5               g236(.a(new_n331), .o1(new_n332));
  inv000aa1d42x5               g237(.a(new_n325), .o1(new_n333));
  aoai13aa1n03x5               g238(.a(new_n332), .b(new_n333), .c(new_n320), .d(new_n323), .o1(new_n334));
  xorc02aa1n02x5               g239(.a(\a[28] ), .b(\b[27] ), .out0(new_n335));
  norp02aa1n02x5               g240(.a(new_n335), .b(new_n331), .o1(new_n336));
  aoi022aa1n03x5               g241(.a(new_n334), .b(new_n335), .c(new_n330), .d(new_n336), .o1(\s[28] ));
  and002aa1n02x5               g242(.a(new_n335), .b(new_n325), .o(new_n338));
  aoai13aa1n03x5               g243(.a(new_n338), .b(new_n329), .c(new_n214), .d(new_n319), .o1(new_n339));
  inv000aa1d42x5               g244(.a(new_n338), .o1(new_n340));
  oao003aa1n03x5               g245(.a(\a[28] ), .b(\b[27] ), .c(new_n332), .carry(new_n341));
  aoai13aa1n02x7               g246(.a(new_n341), .b(new_n340), .c(new_n320), .d(new_n323), .o1(new_n342));
  xorc02aa1n02x5               g247(.a(\a[29] ), .b(\b[28] ), .out0(new_n343));
  norb02aa1n02x5               g248(.a(new_n341), .b(new_n343), .out0(new_n344));
  aoi022aa1n02x7               g249(.a(new_n342), .b(new_n343), .c(new_n339), .d(new_n344), .o1(\s[29] ));
  xorb03aa1n02x5               g250(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g251(.a(new_n333), .b(new_n335), .c(new_n343), .out0(new_n347));
  aoai13aa1n03x5               g252(.a(new_n347), .b(new_n329), .c(new_n214), .d(new_n319), .o1(new_n348));
  inv000aa1d42x5               g253(.a(new_n347), .o1(new_n349));
  oao003aa1n02x5               g254(.a(\a[29] ), .b(\b[28] ), .c(new_n341), .carry(new_n350));
  aoai13aa1n03x5               g255(.a(new_n350), .b(new_n349), .c(new_n320), .d(new_n323), .o1(new_n351));
  xorc02aa1n02x5               g256(.a(\a[30] ), .b(\b[29] ), .out0(new_n352));
  norb02aa1n02x5               g257(.a(new_n350), .b(new_n352), .out0(new_n353));
  aoi022aa1n03x5               g258(.a(new_n351), .b(new_n352), .c(new_n348), .d(new_n353), .o1(\s[30] ));
  nano32aa1n03x7               g259(.a(new_n333), .b(new_n352), .c(new_n335), .d(new_n343), .out0(new_n355));
  aoai13aa1n03x5               g260(.a(new_n355), .b(new_n329), .c(new_n214), .d(new_n319), .o1(new_n356));
  xorc02aa1n02x5               g261(.a(\a[31] ), .b(\b[30] ), .out0(new_n357));
  and002aa1n02x5               g262(.a(\b[29] ), .b(\a[30] ), .o(new_n358));
  oabi12aa1n02x5               g263(.a(new_n357), .b(\a[30] ), .c(\b[29] ), .out0(new_n359));
  oab012aa1n02x4               g264(.a(new_n359), .b(new_n350), .c(new_n358), .out0(new_n360));
  inv000aa1d42x5               g265(.a(new_n355), .o1(new_n361));
  oao003aa1n02x5               g266(.a(\a[30] ), .b(\b[29] ), .c(new_n350), .carry(new_n362));
  aoai13aa1n02x7               g267(.a(new_n362), .b(new_n361), .c(new_n320), .d(new_n323), .o1(new_n363));
  aoi022aa1n02x7               g268(.a(new_n363), .b(new_n357), .c(new_n356), .d(new_n360), .o1(\s[31] ));
  xnbna2aa1n03x5               g269(.a(new_n135), .b(new_n100), .c(new_n97), .out0(\s[3] ));
  norb02aa1n02x5               g270(.a(new_n104), .b(new_n105), .out0(new_n366));
  aoi012aa1n02x5               g271(.a(new_n101), .b(new_n134), .c(new_n135), .o1(new_n367));
  oai012aa1n02x5               g272(.a(new_n107), .b(new_n367), .c(new_n366), .o1(\s[4] ));
  xnrc02aa1n02x5               g273(.a(\b[4] ), .b(\a[5] ), .out0(new_n369));
  aoai13aa1n02x5               g274(.a(new_n104), .b(new_n136), .c(new_n134), .d(new_n135), .o1(new_n370));
  and002aa1n02x5               g275(.a(\b[4] ), .b(\a[5] ), .o(new_n371));
  aoi112aa1n02x5               g276(.a(new_n371), .b(new_n109), .c(\a[4] ), .d(\b[3] ), .o1(new_n372));
  aoi022aa1n02x5               g277(.a(new_n370), .b(new_n369), .c(new_n107), .d(new_n372), .o1(\s[5] ));
  aoai13aa1n02x5               g278(.a(new_n372), .b(new_n136), .c(new_n134), .d(new_n135), .o1(new_n374));
  xnbna2aa1n03x5               g279(.a(new_n124), .b(new_n374), .c(new_n118), .out0(\s[6] ));
  nanb02aa1n02x5               g280(.a(new_n143), .b(new_n374), .out0(new_n376));
  nanb02aa1n02x5               g281(.a(new_n108), .b(new_n114), .out0(new_n377));
  aoai13aa1n02x5               g282(.a(new_n113), .b(new_n143), .c(new_n107), .d(new_n372), .o1(new_n378));
  aoi022aa1n02x5               g283(.a(new_n378), .b(new_n377), .c(new_n376), .d(new_n144), .o1(\s[7] ));
  aoi022aa1n02x5               g284(.a(new_n376), .b(new_n144), .c(new_n119), .d(new_n120), .o1(new_n380));
  xnrc02aa1n02x5               g285(.a(new_n380), .b(new_n145), .out0(\s[8] ));
  xorb03aa1n02x5               g286(.a(new_n147), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


