// Benchmark "adder" written by ABC on Wed Jul 17 23:25:45 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n337,
    new_n338, new_n339, new_n340, new_n342, new_n343, new_n345, new_n346,
    new_n347, new_n348, new_n350, new_n352, new_n353, new_n354, new_n356,
    new_n358;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n12x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  norp02aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  orn002aa1n02x7               g003(.a(\a[2] ), .b(\b[1] ), .o(new_n99));
  nand22aa1n06x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  aoi012aa1n12x5               g005(.a(new_n100), .b(\a[2] ), .c(\b[1] ), .o1(new_n101));
  tech160nm_finand02aa1n03p5x5 g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  tech160nm_finand02aa1n03p5x5 g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nor002aa1d32x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanb03aa1n06x5               g009(.a(new_n104), .b(new_n102), .c(new_n103), .out0(new_n105));
  oab012aa1n02x5               g010(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .out0(new_n106));
  aoai13aa1n06x5               g011(.a(new_n106), .b(new_n105), .c(new_n99), .d(new_n101), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\a[7] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[6] ), .o1(new_n109));
  nanp02aa1n02x5               g014(.a(\b[4] ), .b(\a[5] ), .o1(new_n110));
  nand42aa1n02x5               g015(.a(\b[3] ), .b(\a[4] ), .o1(new_n111));
  oai112aa1n02x5               g016(.a(new_n110), .b(new_n111), .c(new_n109), .d(new_n108), .o1(new_n112));
  xnrc02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .out0(new_n113));
  inv000aa1d42x5               g018(.a(\a[6] ), .o1(new_n114));
  inv000aa1d42x5               g019(.a(\b[5] ), .o1(new_n115));
  nor002aa1d32x5               g020(.a(\b[4] ), .b(\a[5] ), .o1(new_n116));
  aoi012aa1d24x5               g021(.a(new_n116), .b(new_n114), .c(new_n115), .o1(new_n117));
  nor042aa1d18x5               g022(.a(\b[6] ), .b(\a[7] ), .o1(new_n118));
  aoi012aa1n02x5               g023(.a(new_n118), .b(\a[6] ), .c(\b[5] ), .o1(new_n119));
  nanp02aa1n02x5               g024(.a(new_n117), .b(new_n119), .o1(new_n120));
  nona32aa1n09x5               g025(.a(new_n107), .b(new_n120), .c(new_n113), .d(new_n112), .out0(new_n121));
  xorc02aa1n12x5               g026(.a(\a[8] ), .b(\b[7] ), .out0(new_n122));
  inv000aa1d42x5               g027(.a(new_n117), .o1(new_n123));
  inv040aa1n02x5               g028(.a(new_n118), .o1(new_n124));
  oaoi03aa1n02x5               g029(.a(\a[8] ), .b(\b[7] ), .c(new_n124), .o1(new_n125));
  and002aa1n03x5               g030(.a(\b[6] ), .b(\a[7] ), .o(new_n126));
  aoi112aa1n03x5               g031(.a(new_n126), .b(new_n118), .c(\a[6] ), .d(\b[5] ), .o1(new_n127));
  aoi013aa1n09x5               g032(.a(new_n125), .b(new_n127), .c(new_n122), .d(new_n123), .o1(new_n128));
  nanp02aa1n03x5               g033(.a(new_n121), .b(new_n128), .o1(new_n129));
  xorc02aa1n12x5               g034(.a(\a[9] ), .b(\b[8] ), .out0(new_n130));
  aoai13aa1n02x5               g035(.a(new_n97), .b(new_n98), .c(new_n129), .d(new_n130), .o1(new_n131));
  norp02aa1n02x5               g036(.a(new_n97), .b(new_n98), .o1(new_n132));
  aob012aa1n03x5               g037(.a(new_n132), .b(new_n129), .c(new_n130), .out0(new_n133));
  nanp02aa1n02x5               g038(.a(new_n131), .b(new_n133), .o1(\s[10] ));
  nor042aa1d18x5               g039(.a(\b[10] ), .b(\a[11] ), .o1(new_n135));
  nand02aa1d12x5               g040(.a(\b[10] ), .b(\a[11] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  aob012aa1n02x5               g042(.a(new_n133), .b(\b[9] ), .c(\a[10] ), .out0(new_n138));
  aoi012aa1n09x5               g043(.a(new_n135), .b(\a[10] ), .c(\b[9] ), .o1(new_n139));
  nand23aa1n03x5               g044(.a(new_n133), .b(new_n136), .c(new_n139), .o1(new_n140));
  aobi12aa1n02x5               g045(.a(new_n140), .b(new_n138), .c(new_n137), .out0(\s[11] ));
  inv000aa1d42x5               g046(.a(\a[11] ), .o1(new_n142));
  oaib12aa1n02x5               g047(.a(new_n140), .b(\b[10] ), .c(new_n142), .out0(new_n143));
  nor002aa1d32x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand02aa1n16x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  norb02aa1n02x5               g050(.a(new_n145), .b(new_n144), .out0(new_n146));
  inv000aa1d42x5               g051(.a(\b[10] ), .o1(new_n147));
  aboi22aa1n03x5               g052(.a(new_n144), .b(new_n145), .c(new_n142), .d(new_n147), .out0(new_n148));
  aoi022aa1n03x5               g053(.a(new_n143), .b(new_n146), .c(new_n140), .d(new_n148), .o1(\s[12] ));
  nona23aa1n09x5               g054(.a(new_n145), .b(new_n136), .c(new_n135), .d(new_n144), .out0(new_n150));
  norb03aa1d15x5               g055(.a(new_n130), .b(new_n150), .c(new_n97), .out0(new_n151));
  nanp02aa1n02x5               g056(.a(new_n129), .b(new_n151), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n151), .o1(new_n153));
  aoai13aa1n12x5               g058(.a(new_n145), .b(new_n144), .c(new_n142), .d(new_n147), .o1(new_n154));
  nanb03aa1n12x5               g059(.a(new_n144), .b(new_n145), .c(new_n136), .out0(new_n155));
  oai022aa1d18x5               g060(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n156));
  nand02aa1n08x5               g061(.a(new_n139), .b(new_n156), .o1(new_n157));
  oai012aa1d24x5               g062(.a(new_n154), .b(new_n157), .c(new_n155), .o1(new_n158));
  inv000aa1d42x5               g063(.a(new_n158), .o1(new_n159));
  aoai13aa1n04x5               g064(.a(new_n159), .b(new_n153), .c(new_n121), .d(new_n128), .o1(new_n160));
  nor002aa1d32x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  nand02aa1n06x5               g066(.a(\b[12] ), .b(\a[13] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  oaib12aa1n02x5               g068(.a(new_n154), .b(new_n161), .c(new_n162), .out0(new_n164));
  oab012aa1n02x4               g069(.a(new_n164), .b(new_n157), .c(new_n155), .out0(new_n165));
  aoi022aa1n02x5               g070(.a(new_n160), .b(new_n163), .c(new_n152), .d(new_n165), .o1(\s[13] ));
  inv000aa1d42x5               g071(.a(new_n161), .o1(new_n167));
  nanp02aa1n02x5               g072(.a(new_n160), .b(new_n163), .o1(new_n168));
  norp02aa1n12x5               g073(.a(\b[13] ), .b(\a[14] ), .o1(new_n169));
  nand42aa1n06x5               g074(.a(\b[13] ), .b(\a[14] ), .o1(new_n170));
  norb02aa1n02x5               g075(.a(new_n170), .b(new_n169), .out0(new_n171));
  xnbna2aa1n03x5               g076(.a(new_n171), .b(new_n168), .c(new_n167), .out0(\s[14] ));
  nona23aa1d18x5               g077(.a(new_n170), .b(new_n162), .c(new_n161), .d(new_n169), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  oaoi03aa1n02x5               g079(.a(\a[14] ), .b(\b[13] ), .c(new_n167), .o1(new_n175));
  nor042aa1n02x5               g080(.a(\b[14] ), .b(\a[15] ), .o1(new_n176));
  nand42aa1n02x5               g081(.a(\b[14] ), .b(\a[15] ), .o1(new_n177));
  norb02aa1n02x7               g082(.a(new_n177), .b(new_n176), .out0(new_n178));
  aoai13aa1n02x5               g083(.a(new_n178), .b(new_n175), .c(new_n160), .d(new_n174), .o1(new_n179));
  aoi112aa1n02x5               g084(.a(new_n178), .b(new_n175), .c(new_n160), .d(new_n174), .o1(new_n180));
  norb02aa1n02x5               g085(.a(new_n179), .b(new_n180), .out0(\s[15] ));
  inv000aa1d42x5               g086(.a(\a[15] ), .o1(new_n182));
  oaib12aa1n02x5               g087(.a(new_n179), .b(\b[14] ), .c(new_n182), .out0(new_n183));
  nor042aa1n04x5               g088(.a(\b[15] ), .b(\a[16] ), .o1(new_n184));
  nand02aa1d04x5               g089(.a(\b[15] ), .b(\a[16] ), .o1(new_n185));
  norb02aa1n03x5               g090(.a(new_n185), .b(new_n184), .out0(new_n186));
  norp02aa1n02x5               g091(.a(new_n186), .b(new_n176), .o1(new_n187));
  aoi022aa1n02x5               g092(.a(new_n183), .b(new_n186), .c(new_n179), .d(new_n187), .o1(\s[16] ));
  nano22aa1n06x5               g093(.a(new_n173), .b(new_n178), .c(new_n186), .out0(new_n189));
  nand02aa1d04x5               g094(.a(new_n151), .b(new_n189), .o1(new_n190));
  aoi012aa1n02x5               g095(.a(new_n190), .b(new_n121), .c(new_n128), .o1(new_n191));
  nanb03aa1n02x5               g096(.a(new_n184), .b(new_n185), .c(new_n177), .out0(new_n192));
  oai122aa1n02x7               g097(.a(new_n170), .b(new_n169), .c(new_n161), .d(\b[14] ), .e(\a[15] ), .o1(new_n193));
  aoi012aa1n02x5               g098(.a(new_n184), .b(new_n176), .c(new_n185), .o1(new_n194));
  oai012aa1n03x5               g099(.a(new_n194), .b(new_n193), .c(new_n192), .o1(new_n195));
  aoi012aa1n06x5               g100(.a(new_n195), .b(new_n158), .c(new_n189), .o1(new_n196));
  aoai13aa1n12x5               g101(.a(new_n196), .b(new_n190), .c(new_n121), .d(new_n128), .o1(new_n197));
  xorc02aa1n06x5               g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  norp02aa1n02x5               g103(.a(new_n193), .b(new_n192), .o1(new_n199));
  nanb02aa1n02x5               g104(.a(new_n198), .b(new_n194), .out0(new_n200));
  aoi112aa1n02x5               g105(.a(new_n200), .b(new_n199), .c(new_n158), .d(new_n189), .o1(new_n201));
  aboi22aa1n03x5               g106(.a(new_n191), .b(new_n201), .c(new_n197), .d(new_n198), .out0(\s[17] ));
  inv000aa1d42x5               g107(.a(\a[17] ), .o1(new_n203));
  nanb02aa1n02x5               g108(.a(\b[16] ), .b(new_n203), .out0(new_n204));
  nanp02aa1n02x5               g109(.a(new_n197), .b(new_n198), .o1(new_n205));
  tech160nm_fixorc02aa1n03p5x5 g110(.a(\a[18] ), .b(\b[17] ), .out0(new_n206));
  xnbna2aa1n03x5               g111(.a(new_n206), .b(new_n205), .c(new_n204), .out0(\s[18] ));
  and002aa1n02x5               g112(.a(new_n206), .b(new_n198), .o(new_n208));
  nand02aa1d04x5               g113(.a(new_n197), .b(new_n208), .o1(new_n209));
  nanp02aa1n02x5               g114(.a(\b[17] ), .b(\a[18] ), .o1(new_n210));
  oai022aa1n06x5               g115(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n211));
  nanp02aa1n02x5               g116(.a(new_n211), .b(new_n210), .o1(new_n212));
  xorc02aa1n02x5               g117(.a(\a[19] ), .b(\b[18] ), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n209), .c(new_n212), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aob012aa1n03x5               g120(.a(new_n213), .b(new_n209), .c(new_n212), .out0(new_n216));
  inv000aa1d42x5               g121(.a(\a[19] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[18] ), .o1(new_n218));
  nand02aa1n02x5               g123(.a(new_n218), .b(new_n217), .o1(new_n219));
  inv000aa1n02x5               g124(.a(new_n213), .o1(new_n220));
  aoai13aa1n02x5               g125(.a(new_n219), .b(new_n220), .c(new_n209), .d(new_n212), .o1(new_n221));
  nor042aa1n06x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nand02aa1n06x5               g127(.a(\b[19] ), .b(\a[20] ), .o1(new_n223));
  norb02aa1n03x5               g128(.a(new_n223), .b(new_n222), .out0(new_n224));
  aboi22aa1n03x5               g129(.a(new_n222), .b(new_n223), .c(new_n217), .d(new_n218), .out0(new_n225));
  aoi022aa1n03x5               g130(.a(new_n221), .b(new_n224), .c(new_n216), .d(new_n225), .o1(\s[20] ));
  nano32aa1n03x7               g131(.a(new_n220), .b(new_n206), .c(new_n198), .d(new_n224), .out0(new_n227));
  nand42aa1n03x5               g132(.a(\b[18] ), .b(\a[19] ), .o1(new_n228));
  nanb03aa1n06x5               g133(.a(new_n222), .b(new_n223), .c(new_n228), .out0(new_n229));
  nand23aa1n03x5               g134(.a(new_n211), .b(new_n219), .c(new_n210), .o1(new_n230));
  aoi013aa1n06x4               g135(.a(new_n222), .b(new_n223), .c(new_n217), .d(new_n218), .o1(new_n231));
  oai012aa1n06x5               g136(.a(new_n231), .b(new_n230), .c(new_n229), .o1(new_n232));
  xorc02aa1n02x5               g137(.a(\a[21] ), .b(\b[20] ), .out0(new_n233));
  aoai13aa1n06x5               g138(.a(new_n233), .b(new_n232), .c(new_n197), .d(new_n227), .o1(new_n234));
  inv000aa1n02x5               g139(.a(new_n233), .o1(new_n235));
  oai112aa1n02x5               g140(.a(new_n235), .b(new_n231), .c(new_n230), .d(new_n229), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n197), .c(new_n227), .o1(new_n237));
  norb02aa1n03x4               g142(.a(new_n234), .b(new_n237), .out0(\s[21] ));
  inv000aa1d42x5               g143(.a(\a[21] ), .o1(new_n239));
  oaib12aa1n06x5               g144(.a(new_n234), .b(\b[20] ), .c(new_n239), .out0(new_n240));
  xorc02aa1n02x5               g145(.a(\a[22] ), .b(\b[21] ), .out0(new_n241));
  norp02aa1n02x5               g146(.a(\b[20] ), .b(\a[21] ), .o1(new_n242));
  norp02aa1n02x5               g147(.a(new_n241), .b(new_n242), .o1(new_n243));
  aoi022aa1n02x7               g148(.a(new_n240), .b(new_n241), .c(new_n234), .d(new_n243), .o1(\s[22] ));
  inv000aa1n02x5               g149(.a(new_n227), .o1(new_n245));
  xnrc02aa1n02x5               g150(.a(\b[21] ), .b(\a[22] ), .out0(new_n246));
  nona32aa1n03x5               g151(.a(new_n197), .b(new_n246), .c(new_n235), .d(new_n245), .out0(new_n247));
  inv000aa1d42x5               g152(.a(\a[22] ), .o1(new_n248));
  xroi22aa1d06x4               g153(.a(new_n239), .b(\b[20] ), .c(new_n248), .d(\b[21] ), .out0(new_n249));
  nand02aa1d06x5               g154(.a(new_n232), .b(new_n249), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\b[21] ), .o1(new_n251));
  oaoi03aa1n02x5               g156(.a(new_n248), .b(new_n251), .c(new_n242), .o1(new_n252));
  nand42aa1n08x5               g157(.a(new_n250), .b(new_n252), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n253), .o1(new_n254));
  tech160nm_fixorc02aa1n03p5x5 g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  aobi12aa1n02x5               g160(.a(new_n255), .b(new_n247), .c(new_n254), .out0(new_n256));
  norb02aa1n02x5               g161(.a(new_n252), .b(new_n255), .out0(new_n257));
  aoi013aa1n02x4               g162(.a(new_n256), .b(new_n250), .c(new_n247), .d(new_n257), .o1(\s[23] ));
  aob012aa1n03x5               g163(.a(new_n255), .b(new_n247), .c(new_n254), .out0(new_n259));
  aoi013aa1n02x4               g164(.a(new_n253), .b(new_n197), .c(new_n227), .d(new_n249), .o1(new_n260));
  oaoi03aa1n02x5               g165(.a(\a[23] ), .b(\b[22] ), .c(new_n260), .o1(new_n261));
  tech160nm_fixorc02aa1n02p5x5 g166(.a(\a[24] ), .b(\b[23] ), .out0(new_n262));
  norp02aa1n02x5               g167(.a(\b[22] ), .b(\a[23] ), .o1(new_n263));
  norp02aa1n02x5               g168(.a(new_n262), .b(new_n263), .o1(new_n264));
  aoi022aa1n03x5               g169(.a(new_n261), .b(new_n262), .c(new_n259), .d(new_n264), .o1(\s[24] ));
  and002aa1n06x5               g170(.a(new_n262), .b(new_n255), .o(new_n266));
  nano22aa1n02x4               g171(.a(new_n245), .b(new_n266), .c(new_n249), .out0(new_n267));
  nand02aa1d04x5               g172(.a(new_n197), .b(new_n267), .o1(new_n268));
  inv000aa1n03x5               g173(.a(new_n263), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[24] ), .b(\b[23] ), .c(new_n269), .carry(new_n270));
  inv000aa1d42x5               g175(.a(new_n270), .o1(new_n271));
  tech160nm_fiaoi012aa1n02p5x5 g176(.a(new_n271), .b(new_n253), .c(new_n266), .o1(new_n272));
  xorc02aa1n12x5               g177(.a(\a[25] ), .b(\b[24] ), .out0(new_n273));
  aob012aa1n03x5               g178(.a(new_n273), .b(new_n268), .c(new_n272), .out0(new_n274));
  aoi112aa1n02x5               g179(.a(new_n273), .b(new_n271), .c(new_n253), .d(new_n266), .o1(new_n275));
  aobi12aa1n02x7               g180(.a(new_n274), .b(new_n275), .c(new_n268), .out0(\s[25] ));
  nor042aa1n03x5               g181(.a(\b[24] ), .b(\a[25] ), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  inv000aa1d42x5               g183(.a(new_n273), .o1(new_n279));
  aoai13aa1n02x5               g184(.a(new_n278), .b(new_n279), .c(new_n268), .d(new_n272), .o1(new_n280));
  xorc02aa1n02x5               g185(.a(\a[26] ), .b(\b[25] ), .out0(new_n281));
  norp02aa1n02x5               g186(.a(new_n281), .b(new_n277), .o1(new_n282));
  aoi022aa1n03x5               g187(.a(new_n280), .b(new_n281), .c(new_n274), .d(new_n282), .o1(\s[26] ));
  and002aa1n02x5               g188(.a(new_n281), .b(new_n273), .o(new_n284));
  aoai13aa1n12x5               g189(.a(new_n284), .b(new_n271), .c(new_n253), .d(new_n266), .o1(new_n285));
  nano32aa1n03x7               g190(.a(new_n245), .b(new_n284), .c(new_n249), .d(new_n266), .out0(new_n286));
  nand22aa1n03x5               g191(.a(new_n197), .b(new_n286), .o1(new_n287));
  oao003aa1n02x5               g192(.a(\a[26] ), .b(\b[25] ), .c(new_n278), .carry(new_n288));
  nand23aa1n03x5               g193(.a(new_n287), .b(new_n285), .c(new_n288), .o1(new_n289));
  nor042aa1n06x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  and002aa1n02x5               g195(.a(\b[26] ), .b(\a[27] ), .o(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n290), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n288), .o1(new_n293));
  aoi112aa1n02x5               g198(.a(new_n292), .b(new_n293), .c(new_n197), .d(new_n286), .o1(new_n294));
  aoi022aa1n02x5               g199(.a(new_n289), .b(new_n292), .c(new_n294), .d(new_n285), .o1(\s[27] ));
  nanp02aa1n03x5               g200(.a(new_n289), .b(new_n292), .o1(new_n296));
  tech160nm_fiaoi012aa1n05x5   g201(.a(new_n293), .b(new_n197), .c(new_n286), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n290), .o1(new_n298));
  aoai13aa1n02x7               g203(.a(new_n298), .b(new_n291), .c(new_n297), .d(new_n285), .o1(new_n299));
  xorc02aa1n02x5               g204(.a(\a[28] ), .b(\b[27] ), .out0(new_n300));
  norp02aa1n02x5               g205(.a(new_n300), .b(new_n290), .o1(new_n301));
  aoi022aa1n03x5               g206(.a(new_n299), .b(new_n300), .c(new_n296), .d(new_n301), .o1(\s[28] ));
  inv000aa1d42x5               g207(.a(\a[27] ), .o1(new_n303));
  inv000aa1d42x5               g208(.a(\a[28] ), .o1(new_n304));
  xroi22aa1d04x5               g209(.a(new_n303), .b(\b[26] ), .c(new_n304), .d(\b[27] ), .out0(new_n305));
  nanp02aa1n03x5               g210(.a(new_n289), .b(new_n305), .o1(new_n306));
  inv000aa1n06x5               g211(.a(new_n305), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n298), .carry(new_n308));
  aoai13aa1n02x7               g213(.a(new_n308), .b(new_n307), .c(new_n297), .d(new_n285), .o1(new_n309));
  xorc02aa1n02x5               g214(.a(\a[29] ), .b(\b[28] ), .out0(new_n310));
  norb02aa1n02x5               g215(.a(new_n308), .b(new_n310), .out0(new_n311));
  aoi022aa1n03x5               g216(.a(new_n309), .b(new_n310), .c(new_n306), .d(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g217(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  and003aa1n02x5               g218(.a(new_n300), .b(new_n310), .c(new_n292), .o(new_n314));
  nanp02aa1n03x5               g219(.a(new_n289), .b(new_n314), .o1(new_n315));
  inv000aa1n02x5               g220(.a(new_n314), .o1(new_n316));
  inv000aa1d42x5               g221(.a(\b[28] ), .o1(new_n317));
  inv000aa1d42x5               g222(.a(\a[29] ), .o1(new_n318));
  oaib12aa1n02x5               g223(.a(new_n308), .b(\b[28] ), .c(new_n318), .out0(new_n319));
  oaib12aa1n02x5               g224(.a(new_n319), .b(new_n317), .c(\a[29] ), .out0(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n316), .c(new_n297), .d(new_n285), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  oaoi13aa1n02x5               g227(.a(new_n322), .b(new_n319), .c(new_n318), .d(new_n317), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n315), .d(new_n323), .o1(\s[30] ));
  nano22aa1n02x4               g229(.a(new_n307), .b(new_n310), .c(new_n322), .out0(new_n325));
  nanp02aa1n03x5               g230(.a(new_n289), .b(new_n325), .o1(new_n326));
  aoi022aa1n02x5               g231(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n327));
  norb02aa1n02x5               g232(.a(\b[30] ), .b(\a[31] ), .out0(new_n328));
  obai22aa1n02x7               g233(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n329));
  aoi112aa1n02x5               g234(.a(new_n329), .b(new_n328), .c(new_n319), .d(new_n327), .o1(new_n330));
  xorc02aa1n02x5               g235(.a(\a[31] ), .b(\b[30] ), .out0(new_n331));
  inv000aa1n02x5               g236(.a(new_n325), .o1(new_n332));
  norp02aa1n02x5               g237(.a(\b[29] ), .b(\a[30] ), .o1(new_n333));
  aoi012aa1n02x5               g238(.a(new_n333), .b(new_n319), .c(new_n327), .o1(new_n334));
  aoai13aa1n02x7               g239(.a(new_n334), .b(new_n332), .c(new_n297), .d(new_n285), .o1(new_n335));
  aoi022aa1n03x5               g240(.a(new_n335), .b(new_n331), .c(new_n326), .d(new_n330), .o1(\s[31] ));
  aoi012aa1n02x5               g241(.a(new_n105), .b(new_n99), .c(new_n101), .o1(new_n337));
  nanp02aa1n02x5               g242(.a(new_n101), .b(new_n99), .o1(new_n338));
  inv000aa1d42x5               g243(.a(new_n104), .o1(new_n339));
  aoi022aa1n02x5               g244(.a(new_n338), .b(new_n102), .c(new_n339), .d(new_n103), .o1(new_n340));
  norp02aa1n02x5               g245(.a(new_n340), .b(new_n337), .o1(\s[3] ));
  inv000aa1n03x5               g246(.a(new_n337), .o1(new_n342));
  xorc02aa1n02x5               g247(.a(\a[4] ), .b(\b[3] ), .out0(new_n343));
  xnbna2aa1n03x5               g248(.a(new_n343), .b(new_n342), .c(new_n339), .out0(\s[4] ));
  nano22aa1n02x4               g249(.a(new_n116), .b(new_n110), .c(new_n111), .out0(new_n345));
  nanp02aa1n02x5               g250(.a(new_n107), .b(new_n345), .o1(new_n346));
  inv000aa1d42x5               g251(.a(new_n116), .o1(new_n347));
  aoi022aa1n02x5               g252(.a(new_n107), .b(new_n111), .c(new_n110), .d(new_n347), .o1(new_n348));
  norb02aa1n02x5               g253(.a(new_n346), .b(new_n348), .out0(\s[5] ));
  xorc02aa1n02x5               g254(.a(\a[6] ), .b(\b[5] ), .out0(new_n350));
  xnbna2aa1n03x5               g255(.a(new_n350), .b(new_n346), .c(new_n347), .out0(\s[6] ));
  nanp02aa1n02x5               g256(.a(new_n115), .b(new_n114), .o1(new_n352));
  aoai13aa1n02x5               g257(.a(new_n350), .b(new_n116), .c(new_n107), .d(new_n345), .o1(new_n353));
  norp02aa1n02x5               g258(.a(new_n126), .b(new_n118), .o1(new_n354));
  xnbna2aa1n03x5               g259(.a(new_n354), .b(new_n353), .c(new_n352), .out0(\s[7] ));
  aob012aa1n02x5               g260(.a(new_n354), .b(new_n353), .c(new_n352), .out0(new_n356));
  xnbna2aa1n03x5               g261(.a(new_n122), .b(new_n356), .c(new_n124), .out0(\s[8] ));
  aoi113aa1n02x5               g262(.a(new_n125), .b(new_n130), .c(new_n127), .d(new_n122), .e(new_n123), .o1(new_n358));
  aoi022aa1n02x5               g263(.a(new_n129), .b(new_n130), .c(new_n121), .d(new_n358), .o1(\s[9] ));
endmodule


