// Benchmark "adder" written by ABC on Wed Jul 17 17:23:22 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n135, new_n136, new_n137, new_n138, new_n139, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n156, new_n157,
    new_n158, new_n159, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n186, new_n187, new_n188,
    new_n189, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n316, new_n319,
    new_n321, new_n322, new_n324;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d32x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  nor002aa1n02x5               g002(.a(\b[3] ), .b(\a[4] ), .o1(new_n98));
  tech160nm_finand02aa1n05x5   g003(.a(\b[3] ), .b(\a[4] ), .o1(new_n99));
  nor042aa1n04x5               g004(.a(\b[2] ), .b(\a[3] ), .o1(new_n100));
  aoi012aa1n02x5               g005(.a(new_n98), .b(new_n100), .c(new_n99), .o1(new_n101));
  inv000aa1d42x5               g006(.a(\a[2] ), .o1(new_n102));
  inv000aa1d42x5               g007(.a(\b[1] ), .o1(new_n103));
  nand22aa1n03x5               g008(.a(\b[0] ), .b(\a[1] ), .o1(new_n104));
  oao003aa1n02x5               g009(.a(new_n102), .b(new_n103), .c(new_n104), .carry(new_n105));
  nand42aa1n03x5               g010(.a(\b[2] ), .b(\a[3] ), .o1(new_n106));
  nano23aa1n02x5               g011(.a(new_n98), .b(new_n100), .c(new_n106), .d(new_n99), .out0(new_n107));
  aobi12aa1n06x5               g012(.a(new_n101), .b(new_n107), .c(new_n105), .out0(new_n108));
  oaih22aa1d12x5               g013(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n109));
  aoi022aa1d24x5               g014(.a(\b[6] ), .b(\a[7] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n110));
  xorc02aa1n03x5               g015(.a(\a[8] ), .b(\b[7] ), .out0(new_n111));
  nand42aa1n08x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  oai122aa1n06x5               g017(.a(new_n112), .b(\a[8] ), .c(\b[7] ), .d(\a[7] ), .e(\b[6] ), .o1(new_n113));
  nona23aa1n09x5               g018(.a(new_n111), .b(new_n110), .c(new_n113), .d(new_n109), .out0(new_n114));
  nanp02aa1n02x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  oai022aa1n02x5               g020(.a(\a[7] ), .b(\b[6] ), .c(\b[7] ), .d(\a[8] ), .o1(new_n116));
  nanp02aa1n02x5               g021(.a(new_n116), .b(new_n115), .o1(new_n117));
  aoi022aa1n02x5               g022(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(new_n109), .b(new_n118), .o1(new_n119));
  oai012aa1n02x5               g024(.a(new_n117), .b(new_n119), .c(new_n113), .o1(new_n120));
  inv000aa1n02x5               g025(.a(new_n120), .o1(new_n121));
  oai012aa1n12x5               g026(.a(new_n121), .b(new_n108), .c(new_n114), .o1(new_n122));
  tech160nm_fixorc02aa1n02p5x5 g027(.a(\a[9] ), .b(\b[8] ), .out0(new_n123));
  tech160nm_fixorc02aa1n04x5   g028(.a(\a[10] ), .b(\b[9] ), .out0(new_n124));
  aoai13aa1n03x5               g029(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n125));
  aoi112aa1n02x5               g030(.a(new_n124), .b(new_n97), .c(new_n122), .d(new_n123), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n125), .b(new_n126), .out0(\s[10] ));
  inv000aa1d42x5               g032(.a(\a[10] ), .o1(new_n128));
  inv040aa1d32x5               g033(.a(\b[9] ), .o1(new_n129));
  oaoi03aa1n12x5               g034(.a(new_n128), .b(new_n129), .c(new_n97), .o1(new_n130));
  nand42aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor002aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  norb02aa1n02x5               g037(.a(new_n131), .b(new_n132), .out0(new_n133));
  xnbna2aa1n03x5               g038(.a(new_n133), .b(new_n125), .c(new_n130), .out0(\s[11] ));
  norp02aa1n04x5               g039(.a(\b[11] ), .b(\a[12] ), .o1(new_n135));
  nanp02aa1n09x5               g040(.a(\b[11] ), .b(\a[12] ), .o1(new_n136));
  nanb02aa1n02x5               g041(.a(new_n135), .b(new_n136), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n130), .o1(new_n138));
  nona22aa1n03x5               g043(.a(new_n125), .b(new_n138), .c(new_n132), .out0(new_n139));
  xnbna2aa1n03x5               g044(.a(new_n137), .b(new_n139), .c(new_n131), .out0(\s[12] ));
  nano23aa1n03x5               g045(.a(new_n135), .b(new_n132), .c(new_n136), .d(new_n131), .out0(new_n141));
  nand03aa1n02x5               g046(.a(new_n141), .b(new_n123), .c(new_n124), .o1(new_n142));
  nanb02aa1n06x5               g047(.a(new_n142), .b(new_n122), .out0(new_n143));
  nona23aa1n12x5               g048(.a(new_n131), .b(new_n136), .c(new_n135), .d(new_n132), .out0(new_n144));
  tech160nm_fioai012aa1n05x5   g049(.a(new_n136), .b(new_n135), .c(new_n132), .o1(new_n145));
  oai012aa1d24x5               g050(.a(new_n145), .b(new_n144), .c(new_n130), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  xorc02aa1n12x5               g052(.a(\a[13] ), .b(\b[12] ), .out0(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n143), .c(new_n147), .out0(\s[13] ));
  nor042aa1d18x5               g054(.a(\b[12] ), .b(\a[13] ), .o1(new_n150));
  inv040aa1n08x5               g055(.a(new_n150), .o1(new_n151));
  nanp02aa1n03x5               g056(.a(new_n143), .b(new_n147), .o1(new_n152));
  nanp02aa1n03x5               g057(.a(new_n152), .b(new_n148), .o1(new_n153));
  xorc02aa1n12x5               g058(.a(\a[14] ), .b(\b[13] ), .out0(new_n154));
  xnbna2aa1n03x5               g059(.a(new_n154), .b(new_n153), .c(new_n151), .out0(\s[14] ));
  nanp02aa1n02x5               g060(.a(new_n154), .b(new_n148), .o1(new_n156));
  oaoi03aa1n12x5               g061(.a(\a[14] ), .b(\b[13] ), .c(new_n151), .o1(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  aoai13aa1n04x5               g063(.a(new_n158), .b(new_n156), .c(new_n143), .d(new_n147), .o1(new_n159));
  xorb03aa1n02x5               g064(.a(new_n159), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n04x5               g065(.a(\b[14] ), .b(\a[15] ), .o1(new_n161));
  nand22aa1n09x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  norb02aa1n02x5               g067(.a(new_n162), .b(new_n161), .out0(new_n163));
  nor042aa1n02x5               g068(.a(\b[15] ), .b(\a[16] ), .o1(new_n164));
  nand22aa1n09x5               g069(.a(\b[15] ), .b(\a[16] ), .o1(new_n165));
  nanb02aa1n02x5               g070(.a(new_n164), .b(new_n165), .out0(new_n166));
  aoai13aa1n02x5               g071(.a(new_n166), .b(new_n161), .c(new_n159), .d(new_n163), .o1(new_n167));
  nanp02aa1n02x5               g072(.a(new_n159), .b(new_n163), .o1(new_n168));
  nona22aa1n02x4               g073(.a(new_n168), .b(new_n166), .c(new_n161), .out0(new_n169));
  nanp02aa1n02x5               g074(.a(new_n169), .b(new_n167), .o1(\s[16] ));
  oaoi03aa1n02x5               g075(.a(new_n102), .b(new_n103), .c(new_n104), .o1(new_n171));
  nona23aa1n02x4               g076(.a(new_n106), .b(new_n99), .c(new_n98), .d(new_n100), .out0(new_n172));
  oai012aa1n02x7               g077(.a(new_n101), .b(new_n172), .c(new_n171), .o1(new_n173));
  oai122aa1n02x7               g078(.a(new_n110), .b(\a[6] ), .c(\b[5] ), .d(\a[5] ), .e(\b[4] ), .o1(new_n174));
  norb03aa1n02x5               g079(.a(new_n111), .b(new_n174), .c(new_n113), .out0(new_n175));
  nano23aa1n06x5               g080(.a(new_n164), .b(new_n161), .c(new_n165), .d(new_n162), .out0(new_n176));
  nand23aa1n03x5               g081(.a(new_n176), .b(new_n148), .c(new_n154), .o1(new_n177));
  nor042aa1n06x5               g082(.a(new_n177), .b(new_n142), .o1(new_n178));
  aoai13aa1n06x5               g083(.a(new_n178), .b(new_n120), .c(new_n173), .d(new_n175), .o1(new_n179));
  norb02aa1n03x5               g084(.a(new_n176), .b(new_n156), .out0(new_n180));
  tech160nm_fiao0012aa1n02p5x5 g085(.a(new_n164), .b(new_n161), .c(new_n165), .o(new_n181));
  aoi012aa1n06x5               g086(.a(new_n181), .b(new_n176), .c(new_n157), .o1(new_n182));
  aobi12aa1n12x5               g087(.a(new_n182), .b(new_n180), .c(new_n146), .out0(new_n183));
  nanp02aa1n06x5               g088(.a(new_n179), .b(new_n183), .o1(new_n184));
  xorb03aa1n02x5               g089(.a(new_n184), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g090(.a(\a[18] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\a[17] ), .o1(new_n187));
  inv000aa1d42x5               g092(.a(\b[16] ), .o1(new_n188));
  oaoi03aa1n02x5               g093(.a(new_n187), .b(new_n188), .c(new_n184), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[17] ), .c(new_n186), .out0(\s[18] ));
  xroi22aa1d04x5               g095(.a(new_n187), .b(\b[16] ), .c(new_n186), .d(\b[17] ), .out0(new_n191));
  nanp02aa1n02x5               g096(.a(\b[17] ), .b(\a[18] ), .o1(new_n192));
  nona22aa1n02x4               g097(.a(new_n192), .b(\b[16] ), .c(\a[17] ), .out0(new_n193));
  oaib12aa1n02x5               g098(.a(new_n193), .b(\b[17] ), .c(new_n186), .out0(new_n194));
  nanp02aa1n03x5               g099(.a(\b[18] ), .b(\a[19] ), .o1(new_n195));
  nor002aa1n12x5               g100(.a(\b[18] ), .b(\a[19] ), .o1(new_n196));
  norb02aa1n02x5               g101(.a(new_n195), .b(new_n196), .out0(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n194), .c(new_n184), .d(new_n191), .o1(new_n198));
  aoi112aa1n02x5               g103(.a(new_n197), .b(new_n194), .c(new_n184), .d(new_n191), .o1(new_n199));
  norb02aa1n02x5               g104(.a(new_n198), .b(new_n199), .out0(\s[19] ));
  xnrc02aa1n02x5               g105(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor022aa1n08x5               g106(.a(\b[19] ), .b(\a[20] ), .o1(new_n202));
  nand02aa1n04x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  nanb02aa1n02x5               g108(.a(new_n202), .b(new_n203), .out0(new_n204));
  tech160nm_fioai012aa1n03p5x5 g109(.a(new_n198), .b(\b[18] ), .c(\a[19] ), .o1(new_n205));
  nanp02aa1n03x5               g110(.a(new_n205), .b(new_n204), .o1(new_n206));
  nona22aa1n02x4               g111(.a(new_n198), .b(new_n204), .c(new_n196), .out0(new_n207));
  nanp02aa1n03x5               g112(.a(new_n206), .b(new_n207), .o1(\s[20] ));
  nano23aa1n02x5               g113(.a(new_n202), .b(new_n196), .c(new_n203), .d(new_n195), .out0(new_n209));
  nand02aa1n02x5               g114(.a(new_n191), .b(new_n209), .o1(new_n210));
  norp02aa1n02x5               g115(.a(\b[17] ), .b(\a[18] ), .o1(new_n211));
  aoi013aa1n06x4               g116(.a(new_n211), .b(new_n192), .c(new_n187), .d(new_n188), .o1(new_n212));
  nona23aa1n06x5               g117(.a(new_n195), .b(new_n203), .c(new_n202), .d(new_n196), .out0(new_n213));
  tech160nm_fioai012aa1n05x5   g118(.a(new_n203), .b(new_n202), .c(new_n196), .o1(new_n214));
  oai012aa1n12x5               g119(.a(new_n214), .b(new_n213), .c(new_n212), .o1(new_n215));
  inv000aa1d42x5               g120(.a(new_n215), .o1(new_n216));
  aoai13aa1n06x5               g121(.a(new_n216), .b(new_n210), .c(new_n179), .d(new_n183), .o1(new_n217));
  xorb03aa1n02x5               g122(.a(new_n217), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g123(.a(\b[20] ), .b(\a[21] ), .o1(new_n219));
  xorc02aa1n02x5               g124(.a(\a[21] ), .b(\b[20] ), .out0(new_n220));
  xorc02aa1n02x5               g125(.a(\a[22] ), .b(\b[21] ), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n02x5               g127(.a(new_n222), .b(new_n219), .c(new_n217), .d(new_n220), .o1(new_n223));
  aoi112aa1n02x7               g128(.a(new_n219), .b(new_n222), .c(new_n217), .d(new_n220), .o1(new_n224));
  nanb02aa1n02x5               g129(.a(new_n224), .b(new_n223), .out0(\s[22] ));
  inv030aa1d32x5               g130(.a(\a[21] ), .o1(new_n226));
  inv040aa1d32x5               g131(.a(\a[22] ), .o1(new_n227));
  xroi22aa1d06x4               g132(.a(new_n226), .b(\b[20] ), .c(new_n227), .d(\b[21] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(\b[21] ), .o1(new_n229));
  oao003aa1n12x5               g134(.a(new_n227), .b(new_n229), .c(new_n219), .carry(new_n230));
  aoi012aa1n02x5               g135(.a(new_n230), .b(new_n215), .c(new_n228), .o1(new_n231));
  inv000aa1d42x5               g136(.a(new_n228), .o1(new_n232));
  nona22aa1n03x5               g137(.a(new_n184), .b(new_n210), .c(new_n232), .out0(new_n233));
  tech160nm_fixnrc02aa1n05x5   g138(.a(\b[22] ), .b(\a[23] ), .out0(new_n234));
  xobna2aa1n03x5               g139(.a(new_n234), .b(new_n233), .c(new_n231), .out0(\s[23] ));
  and002aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o(new_n236));
  xorc02aa1n12x5               g141(.a(\a[24] ), .b(\b[23] ), .out0(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  inv000aa1n02x5               g143(.a(new_n214), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n228), .b(new_n239), .c(new_n209), .d(new_n194), .o1(new_n240));
  nor042aa1d18x5               g145(.a(\b[22] ), .b(\a[23] ), .o1(new_n241));
  nona22aa1n02x4               g146(.a(new_n240), .b(new_n230), .c(new_n241), .out0(new_n242));
  inv000aa1n02x5               g147(.a(new_n242), .o1(new_n243));
  aoai13aa1n03x5               g148(.a(new_n238), .b(new_n236), .c(new_n233), .d(new_n243), .o1(new_n244));
  aoi112aa1n02x7               g149(.a(new_n238), .b(new_n236), .c(new_n233), .d(new_n243), .o1(new_n245));
  norb02aa1n03x4               g150(.a(new_n244), .b(new_n245), .out0(\s[24] ));
  oaib12aa1n09x5               g151(.a(new_n182), .b(new_n177), .c(new_n146), .out0(new_n247));
  norb02aa1n02x5               g152(.a(new_n237), .b(new_n234), .out0(new_n248));
  nano22aa1n03x5               g153(.a(new_n210), .b(new_n248), .c(new_n228), .out0(new_n249));
  aoai13aa1n06x5               g154(.a(new_n249), .b(new_n247), .c(new_n122), .d(new_n178), .o1(new_n250));
  aoai13aa1n06x5               g155(.a(new_n248), .b(new_n230), .c(new_n215), .d(new_n228), .o1(new_n251));
  inv020aa1n04x5               g156(.a(new_n241), .o1(new_n252));
  oaoi03aa1n02x5               g157(.a(\a[24] ), .b(\b[23] ), .c(new_n252), .o1(new_n253));
  inv040aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  nanp03aa1n03x5               g159(.a(new_n250), .b(new_n251), .c(new_n254), .o1(new_n255));
  xorb03aa1n02x5               g160(.a(new_n255), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g161(.a(\b[24] ), .b(\a[25] ), .o1(new_n257));
  xorc02aa1n03x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  nor042aa1n03x5               g163(.a(\b[25] ), .b(\a[26] ), .o1(new_n259));
  nand02aa1d08x5               g164(.a(\b[25] ), .b(\a[26] ), .o1(new_n260));
  norb02aa1n02x5               g165(.a(new_n260), .b(new_n259), .out0(new_n261));
  inv040aa1n03x5               g166(.a(new_n261), .o1(new_n262));
  aoai13aa1n03x5               g167(.a(new_n262), .b(new_n257), .c(new_n255), .d(new_n258), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n230), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n248), .o1(new_n265));
  aoai13aa1n04x5               g170(.a(new_n254), .b(new_n265), .c(new_n240), .d(new_n264), .o1(new_n266));
  aoai13aa1n02x5               g171(.a(new_n258), .b(new_n266), .c(new_n184), .d(new_n249), .o1(new_n267));
  nona22aa1n02x4               g172(.a(new_n267), .b(new_n262), .c(new_n257), .out0(new_n268));
  nanp02aa1n03x5               g173(.a(new_n263), .b(new_n268), .o1(\s[26] ));
  norb02aa1n03x5               g174(.a(new_n258), .b(new_n262), .out0(new_n270));
  inv000aa1n02x5               g175(.a(new_n270), .o1(new_n271));
  nano23aa1n06x5               g176(.a(new_n271), .b(new_n210), .c(new_n248), .d(new_n228), .out0(new_n272));
  aoai13aa1n12x5               g177(.a(new_n272), .b(new_n247), .c(new_n122), .d(new_n178), .o1(new_n273));
  oai012aa1n02x5               g178(.a(new_n260), .b(new_n259), .c(new_n257), .o1(new_n274));
  aobi12aa1n06x5               g179(.a(new_n274), .b(new_n266), .c(new_n270), .out0(new_n275));
  norp02aa1n02x5               g180(.a(\b[26] ), .b(\a[27] ), .o1(new_n276));
  nanp02aa1n02x5               g181(.a(\b[26] ), .b(\a[27] ), .o1(new_n277));
  norb02aa1n02x5               g182(.a(new_n277), .b(new_n276), .out0(new_n278));
  xnbna2aa1n03x5               g183(.a(new_n278), .b(new_n275), .c(new_n273), .out0(\s[27] ));
  norp02aa1n02x5               g184(.a(\b[27] ), .b(\a[28] ), .o1(new_n280));
  nanp02aa1n02x5               g185(.a(\b[27] ), .b(\a[28] ), .o1(new_n281));
  norb02aa1n02x5               g186(.a(new_n281), .b(new_n280), .out0(new_n282));
  oai112aa1n03x5               g187(.a(new_n275), .b(new_n273), .c(\b[26] ), .d(\a[27] ), .o1(new_n283));
  aoi012aa1n03x5               g188(.a(new_n282), .b(new_n283), .c(new_n277), .o1(new_n284));
  aobi12aa1n06x5               g189(.a(new_n272), .b(new_n179), .c(new_n183), .out0(new_n285));
  aoai13aa1n04x5               g190(.a(new_n274), .b(new_n271), .c(new_n251), .d(new_n254), .o1(new_n286));
  norp03aa1n02x5               g191(.a(new_n286), .b(new_n285), .c(new_n276), .o1(new_n287));
  nano22aa1n02x4               g192(.a(new_n287), .b(new_n277), .c(new_n282), .out0(new_n288));
  nor002aa1n02x5               g193(.a(new_n284), .b(new_n288), .o1(\s[28] ));
  nano23aa1n02x4               g194(.a(new_n276), .b(new_n280), .c(new_n281), .d(new_n277), .out0(new_n290));
  oai012aa1n02x5               g195(.a(new_n290), .b(new_n286), .c(new_n285), .o1(new_n291));
  aoi012aa1n02x5               g196(.a(new_n280), .b(new_n276), .c(new_n281), .o1(new_n292));
  xnrc02aa1n02x5               g197(.a(\b[28] ), .b(\a[29] ), .out0(new_n293));
  tech160nm_fiaoi012aa1n02p5x5 g198(.a(new_n293), .b(new_n291), .c(new_n292), .o1(new_n294));
  aobi12aa1n02x7               g199(.a(new_n290), .b(new_n275), .c(new_n273), .out0(new_n295));
  nano22aa1n03x5               g200(.a(new_n295), .b(new_n292), .c(new_n293), .out0(new_n296));
  norp02aa1n03x5               g201(.a(new_n294), .b(new_n296), .o1(\s[29] ));
  xorb03aa1n02x5               g202(.a(new_n104), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g203(.a(new_n293), .b(new_n278), .c(new_n282), .out0(new_n299));
  oai012aa1n02x5               g204(.a(new_n299), .b(new_n286), .c(new_n285), .o1(new_n300));
  oao003aa1n02x5               g205(.a(\a[29] ), .b(\b[28] ), .c(new_n292), .carry(new_n301));
  xnrc02aa1n02x5               g206(.a(\b[29] ), .b(\a[30] ), .out0(new_n302));
  tech160nm_fiaoi012aa1n02p5x5 g207(.a(new_n302), .b(new_n300), .c(new_n301), .o1(new_n303));
  aobi12aa1n02x7               g208(.a(new_n299), .b(new_n275), .c(new_n273), .out0(new_n304));
  nano22aa1n03x5               g209(.a(new_n304), .b(new_n301), .c(new_n302), .out0(new_n305));
  norp02aa1n03x5               g210(.a(new_n303), .b(new_n305), .o1(\s[30] ));
  nano23aa1n02x4               g211(.a(new_n302), .b(new_n293), .c(new_n282), .d(new_n278), .out0(new_n307));
  oai012aa1n02x5               g212(.a(new_n307), .b(new_n286), .c(new_n285), .o1(new_n308));
  oao003aa1n02x5               g213(.a(\a[30] ), .b(\b[29] ), .c(new_n301), .carry(new_n309));
  xnrc02aa1n02x5               g214(.a(\b[30] ), .b(\a[31] ), .out0(new_n310));
  tech160nm_fiaoi012aa1n02p5x5 g215(.a(new_n310), .b(new_n308), .c(new_n309), .o1(new_n311));
  aobi12aa1n02x7               g216(.a(new_n307), .b(new_n275), .c(new_n273), .out0(new_n312));
  nano22aa1n03x5               g217(.a(new_n312), .b(new_n309), .c(new_n310), .out0(new_n313));
  norp02aa1n03x5               g218(.a(new_n311), .b(new_n313), .o1(\s[31] ));
  xnrb03aa1n02x5               g219(.a(new_n171), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g220(.a(\a[3] ), .b(\b[2] ), .c(new_n171), .o1(new_n316));
  xorb03aa1n02x5               g221(.a(new_n316), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g222(.a(new_n173), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g223(.a(\a[5] ), .b(\b[4] ), .c(new_n108), .o1(new_n319));
  xorb03aa1n02x5               g224(.a(new_n319), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  norp02aa1n02x5               g225(.a(\b[5] ), .b(\a[6] ), .o1(new_n321));
  oai012aa1n02x5               g226(.a(new_n112), .b(new_n319), .c(new_n321), .o1(new_n322));
  xnrb03aa1n02x5               g227(.a(new_n322), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g228(.a(\a[7] ), .b(\b[6] ), .c(new_n322), .o1(new_n324));
  xorb03aa1n02x5               g229(.a(new_n324), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g230(.a(new_n122), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


