// Benchmark "adder" written by ABC on Thu Jul 18 03:59:16 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n134, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n332, new_n335, new_n336, new_n338, new_n339, new_n340, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[10] ), .o1(new_n97));
  nor042aa1n02x5               g002(.a(\b[8] ), .b(\a[9] ), .o1(new_n98));
  nor002aa1d32x5               g003(.a(\b[6] ), .b(\a[7] ), .o1(new_n99));
  inv000aa1n02x5               g004(.a(new_n99), .o1(new_n100));
  oaoi03aa1n09x5               g005(.a(\a[8] ), .b(\b[7] ), .c(new_n100), .o1(new_n101));
  nanp02aa1n09x5               g006(.a(\b[7] ), .b(\a[8] ), .o1(new_n102));
  nor042aa1n06x5               g007(.a(\b[7] ), .b(\a[8] ), .o1(new_n103));
  nand42aa1n10x5               g008(.a(\b[6] ), .b(\a[7] ), .o1(new_n104));
  nano23aa1d15x5               g009(.a(new_n99), .b(new_n103), .c(new_n104), .d(new_n102), .out0(new_n105));
  inv040aa1d32x5               g010(.a(\a[5] ), .o1(new_n106));
  inv030aa1d32x5               g011(.a(\b[4] ), .o1(new_n107));
  nand02aa1d04x5               g012(.a(new_n107), .b(new_n106), .o1(new_n108));
  oaoi03aa1n06x5               g013(.a(\a[6] ), .b(\b[5] ), .c(new_n108), .o1(new_n109));
  aoi012aa1d18x5               g014(.a(new_n101), .b(new_n105), .c(new_n109), .o1(new_n110));
  xorc02aa1n02x5               g015(.a(\a[4] ), .b(\b[3] ), .out0(new_n111));
  xorc02aa1n02x5               g016(.a(\a[3] ), .b(\b[2] ), .out0(new_n112));
  nand42aa1n06x5               g017(.a(\b[1] ), .b(\a[2] ), .o1(new_n113));
  nand22aa1n09x5               g018(.a(\b[0] ), .b(\a[1] ), .o1(new_n114));
  nor042aa1n06x5               g019(.a(\b[1] ), .b(\a[2] ), .o1(new_n115));
  oai012aa1n12x5               g020(.a(new_n113), .b(new_n115), .c(new_n114), .o1(new_n116));
  nanb03aa1n03x5               g021(.a(new_n116), .b(new_n111), .c(new_n112), .out0(new_n117));
  inv000aa1d42x5               g022(.a(\a[4] ), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\b[3] ), .o1(new_n119));
  nor042aa1n03x5               g024(.a(\b[2] ), .b(\a[3] ), .o1(new_n120));
  oaoi03aa1n12x5               g025(.a(new_n118), .b(new_n119), .c(new_n120), .o1(new_n121));
  tech160nm_fixnrc02aa1n04x5   g026(.a(\b[5] ), .b(\a[6] ), .out0(new_n122));
  tech160nm_fixnrc02aa1n02p5x5 g027(.a(\b[4] ), .b(\a[5] ), .out0(new_n123));
  nona22aa1n02x4               g028(.a(new_n105), .b(new_n122), .c(new_n123), .out0(new_n124));
  aoai13aa1n06x5               g029(.a(new_n110), .b(new_n124), .c(new_n117), .d(new_n121), .o1(new_n125));
  xorc02aa1n12x5               g030(.a(\a[9] ), .b(\b[8] ), .out0(new_n126));
  aoi012aa1n02x5               g031(.a(new_n98), .b(new_n125), .c(new_n126), .o1(new_n127));
  xorb03aa1n02x5               g032(.a(new_n127), .b(\b[9] ), .c(new_n97), .out0(\s[10] ));
  xorc02aa1n12x5               g033(.a(\a[10] ), .b(\b[9] ), .out0(new_n129));
  inv000aa1d42x5               g034(.a(\b[9] ), .o1(new_n130));
  oao003aa1n02x5               g035(.a(new_n97), .b(new_n130), .c(new_n98), .carry(new_n131));
  aoi013aa1n03x5               g036(.a(new_n131), .b(new_n125), .c(new_n126), .d(new_n129), .o1(new_n132));
  xnrb03aa1n02x5               g037(.a(new_n132), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  oaoi03aa1n02x5               g038(.a(\a[11] ), .b(\b[10] ), .c(new_n132), .o1(new_n134));
  xorb03aa1n02x5               g039(.a(new_n134), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  inv020aa1n03x5               g040(.a(new_n110), .o1(new_n136));
  tech160nm_fixnrc02aa1n02p5x5 g041(.a(\b[3] ), .b(\a[4] ), .out0(new_n137));
  tech160nm_fixnrc02aa1n02p5x5 g042(.a(\b[2] ), .b(\a[3] ), .out0(new_n138));
  oai013aa1n03x5               g043(.a(new_n121), .b(new_n138), .c(new_n137), .d(new_n116), .o1(new_n139));
  norb02aa1n03x5               g044(.a(new_n102), .b(new_n103), .out0(new_n140));
  norb02aa1n06x5               g045(.a(new_n104), .b(new_n99), .out0(new_n141));
  nano23aa1n09x5               g046(.a(new_n123), .b(new_n122), .c(new_n141), .d(new_n140), .out0(new_n142));
  nor042aa1n06x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nand42aa1d28x5               g048(.a(\b[10] ), .b(\a[11] ), .o1(new_n144));
  nor002aa1n12x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nand42aa1n20x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  nano23aa1d15x5               g051(.a(new_n143), .b(new_n145), .c(new_n146), .d(new_n144), .out0(new_n147));
  nand23aa1d12x5               g052(.a(new_n147), .b(new_n126), .c(new_n129), .o1(new_n148));
  inv000aa1d42x5               g053(.a(new_n148), .o1(new_n149));
  aoai13aa1n06x5               g054(.a(new_n149), .b(new_n136), .c(new_n139), .d(new_n142), .o1(new_n150));
  tech160nm_fiaoi012aa1n03p5x5 g055(.a(new_n145), .b(new_n143), .c(new_n146), .o1(new_n151));
  aobi12aa1n06x5               g056(.a(new_n151), .b(new_n147), .c(new_n131), .out0(new_n152));
  nor002aa1d32x5               g057(.a(\b[12] ), .b(\a[13] ), .o1(new_n153));
  nand22aa1n04x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nanb02aa1n02x5               g059(.a(new_n153), .b(new_n154), .out0(new_n155));
  xobna2aa1n03x5               g060(.a(new_n155), .b(new_n150), .c(new_n152), .out0(\s[13] ));
  inv000aa1d42x5               g061(.a(new_n153), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n155), .c(new_n150), .d(new_n152), .o1(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  norp02aa1n24x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nanp02aa1n12x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  nona23aa1n09x5               g066(.a(new_n161), .b(new_n154), .c(new_n153), .d(new_n160), .out0(new_n162));
  oai012aa1d24x5               g067(.a(new_n161), .b(new_n160), .c(new_n153), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n163), .b(new_n162), .c(new_n150), .d(new_n152), .o1(new_n164));
  xorb03aa1n02x5               g069(.a(new_n164), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n03x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  xnrc02aa1n12x5               g071(.a(\b[14] ), .b(\a[15] ), .out0(new_n167));
  inv040aa1n03x5               g072(.a(new_n167), .o1(new_n168));
  xnrc02aa1n12x5               g073(.a(\b[15] ), .b(\a[16] ), .out0(new_n169));
  inv000aa1n02x5               g074(.a(new_n169), .o1(new_n170));
  aoi112aa1n02x5               g075(.a(new_n170), .b(new_n166), .c(new_n164), .d(new_n168), .o1(new_n171));
  nor003aa1n02x5               g076(.a(new_n137), .b(new_n138), .c(new_n116), .o1(new_n172));
  inv000aa1n02x5               g077(.a(new_n121), .o1(new_n173));
  oai012aa1n06x5               g078(.a(new_n142), .b(new_n172), .c(new_n173), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n152), .b(new_n148), .c(new_n174), .d(new_n110), .o1(new_n175));
  nano23aa1n06x5               g080(.a(new_n153), .b(new_n160), .c(new_n161), .d(new_n154), .out0(new_n176));
  inv000aa1d42x5               g081(.a(new_n163), .o1(new_n177));
  aoai13aa1n02x5               g082(.a(new_n168), .b(new_n177), .c(new_n175), .d(new_n176), .o1(new_n178));
  oaoi13aa1n02x5               g083(.a(new_n169), .b(new_n178), .c(\a[15] ), .d(\b[14] ), .o1(new_n179));
  norp02aa1n03x5               g084(.a(new_n179), .b(new_n171), .o1(\s[16] ));
  nano32aa1n03x7               g085(.a(new_n148), .b(new_n170), .c(new_n168), .d(new_n176), .out0(new_n181));
  aoai13aa1n06x5               g086(.a(new_n181), .b(new_n136), .c(new_n139), .d(new_n142), .o1(new_n182));
  oaoi03aa1n02x5               g087(.a(new_n97), .b(new_n130), .c(new_n98), .o1(new_n183));
  nona23aa1n09x5               g088(.a(new_n146), .b(new_n144), .c(new_n143), .d(new_n145), .out0(new_n184));
  tech160nm_fioai012aa1n05x5   g089(.a(new_n151), .b(new_n184), .c(new_n183), .o1(new_n185));
  norp03aa1d12x5               g090(.a(new_n162), .b(new_n169), .c(new_n167), .o1(new_n186));
  inv000aa1n02x5               g091(.a(new_n166), .o1(new_n187));
  oao003aa1n02x5               g092(.a(\a[16] ), .b(\b[15] ), .c(new_n187), .carry(new_n188));
  oai013aa1n09x5               g093(.a(new_n188), .b(new_n169), .c(new_n167), .d(new_n163), .o1(new_n189));
  aoi012aa1d18x5               g094(.a(new_n189), .b(new_n185), .c(new_n186), .o1(new_n190));
  xorc02aa1n02x5               g095(.a(\a[17] ), .b(\b[16] ), .out0(new_n191));
  xnbna2aa1n03x5               g096(.a(new_n191), .b(new_n182), .c(new_n190), .out0(\s[17] ));
  inv040aa1d32x5               g097(.a(\a[17] ), .o1(new_n193));
  inv040aa1d32x5               g098(.a(\b[16] ), .o1(new_n194));
  nanp02aa1n02x5               g099(.a(new_n194), .b(new_n193), .o1(new_n195));
  nona22aa1n02x4               g100(.a(new_n176), .b(new_n169), .c(new_n167), .out0(new_n196));
  oabi12aa1n06x5               g101(.a(new_n189), .b(new_n152), .c(new_n196), .out0(new_n197));
  aoai13aa1n02x5               g102(.a(new_n191), .b(new_n197), .c(new_n125), .d(new_n181), .o1(new_n198));
  nor002aa1d32x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nand42aa1d28x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nanb02aa1n12x5               g105(.a(new_n199), .b(new_n200), .out0(new_n201));
  xobna2aa1n03x5               g106(.a(new_n201), .b(new_n198), .c(new_n195), .out0(\s[18] ));
  nanp02aa1n02x5               g107(.a(\b[16] ), .b(\a[17] ), .o1(new_n203));
  nano22aa1d15x5               g108(.a(new_n201), .b(new_n195), .c(new_n203), .out0(new_n204));
  inv000aa1d42x5               g109(.a(new_n204), .o1(new_n205));
  aoai13aa1n12x5               g110(.a(new_n200), .b(new_n199), .c(new_n193), .d(new_n194), .o1(new_n206));
  aoai13aa1n04x5               g111(.a(new_n206), .b(new_n205), .c(new_n182), .d(new_n190), .o1(new_n207));
  xorb03aa1n02x5               g112(.a(new_n207), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g113(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n24x5               g114(.a(\b[18] ), .b(\a[19] ), .o1(new_n210));
  nanp02aa1n04x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nanb02aa1n09x5               g116(.a(new_n210), .b(new_n211), .out0(new_n212));
  inv000aa1d42x5               g117(.a(new_n212), .o1(new_n213));
  inv000aa1d42x5               g118(.a(\b[19] ), .o1(new_n214));
  nanb02aa1n12x5               g119(.a(\a[20] ), .b(new_n214), .out0(new_n215));
  nanp02aa1n04x5               g120(.a(\b[19] ), .b(\a[20] ), .o1(new_n216));
  nanp02aa1n09x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  inv000aa1d42x5               g122(.a(new_n217), .o1(new_n218));
  aoi112aa1n03x4               g123(.a(new_n210), .b(new_n218), .c(new_n207), .d(new_n213), .o1(new_n219));
  nanb02aa1n12x5               g124(.a(new_n148), .b(new_n186), .out0(new_n220));
  aoai13aa1n12x5               g125(.a(new_n190), .b(new_n220), .c(new_n174), .d(new_n110), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n206), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n213), .b(new_n222), .c(new_n221), .d(new_n204), .o1(new_n223));
  oaoi13aa1n06x5               g128(.a(new_n217), .b(new_n223), .c(\a[19] ), .d(\b[18] ), .o1(new_n224));
  norp02aa1n03x5               g129(.a(new_n224), .b(new_n219), .o1(\s[20] ));
  nona22aa1d18x5               g130(.a(new_n204), .b(new_n212), .c(new_n217), .out0(new_n226));
  nanp02aa1n02x5               g131(.a(new_n210), .b(new_n216), .o1(new_n227));
  nor043aa1n03x5               g132(.a(new_n206), .b(new_n212), .c(new_n217), .o1(new_n228));
  nano22aa1n03x7               g133(.a(new_n228), .b(new_n215), .c(new_n227), .out0(new_n229));
  aoai13aa1n06x5               g134(.a(new_n229), .b(new_n226), .c(new_n182), .d(new_n190), .o1(new_n230));
  xorb03aa1n02x5               g135(.a(new_n230), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g136(.a(\b[20] ), .b(\a[21] ), .o1(new_n232));
  xnrc02aa1n12x5               g137(.a(\b[20] ), .b(\a[21] ), .out0(new_n233));
  inv000aa1d42x5               g138(.a(new_n233), .o1(new_n234));
  xnrc02aa1n12x5               g139(.a(\b[21] ), .b(\a[22] ), .out0(new_n235));
  inv000aa1d42x5               g140(.a(new_n235), .o1(new_n236));
  aoi112aa1n03x4               g141(.a(new_n232), .b(new_n236), .c(new_n230), .d(new_n234), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n226), .o1(new_n238));
  norp02aa1n24x5               g143(.a(\b[19] ), .b(\a[20] ), .o1(new_n239));
  nona23aa1n06x5               g144(.a(new_n216), .b(new_n211), .c(new_n210), .d(new_n239), .out0(new_n240));
  oai112aa1n06x5               g145(.a(new_n227), .b(new_n215), .c(new_n240), .d(new_n206), .o1(new_n241));
  aoai13aa1n06x5               g146(.a(new_n234), .b(new_n241), .c(new_n221), .d(new_n238), .o1(new_n242));
  oaoi13aa1n06x5               g147(.a(new_n235), .b(new_n242), .c(\a[21] ), .d(\b[20] ), .o1(new_n243));
  norp02aa1n03x5               g148(.a(new_n243), .b(new_n237), .o1(\s[22] ));
  nor042aa1n06x5               g149(.a(new_n235), .b(new_n233), .o1(new_n245));
  inv000aa1d42x5               g150(.a(\a[22] ), .o1(new_n246));
  inv000aa1d42x5               g151(.a(\b[21] ), .o1(new_n247));
  oao003aa1n02x5               g152(.a(new_n246), .b(new_n247), .c(new_n232), .carry(new_n248));
  aoi012aa1n02x7               g153(.a(new_n248), .b(new_n241), .c(new_n245), .o1(new_n249));
  inv040aa1n02x5               g154(.a(new_n240), .o1(new_n250));
  nand23aa1d12x5               g155(.a(new_n250), .b(new_n245), .c(new_n204), .o1(new_n251));
  aoai13aa1n06x5               g156(.a(new_n249), .b(new_n251), .c(new_n182), .d(new_n190), .o1(new_n252));
  xorb03aa1n02x5               g157(.a(new_n252), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g158(.a(\b[22] ), .b(\a[23] ), .o1(new_n254));
  xorc02aa1n12x5               g159(.a(\a[23] ), .b(\b[22] ), .out0(new_n255));
  xorc02aa1n12x5               g160(.a(\a[24] ), .b(\b[23] ), .out0(new_n256));
  aoi112aa1n03x4               g161(.a(new_n254), .b(new_n256), .c(new_n252), .d(new_n255), .o1(new_n257));
  inv000aa1d42x5               g162(.a(new_n254), .o1(new_n258));
  inv000aa1n02x5               g163(.a(new_n249), .o1(new_n259));
  inv000aa1d42x5               g164(.a(new_n251), .o1(new_n260));
  aoai13aa1n03x5               g165(.a(new_n255), .b(new_n259), .c(new_n221), .d(new_n260), .o1(new_n261));
  aobi12aa1n06x5               g166(.a(new_n256), .b(new_n261), .c(new_n258), .out0(new_n262));
  nor042aa1n03x5               g167(.a(new_n262), .b(new_n257), .o1(\s[24] ));
  nano32aa1n03x7               g168(.a(new_n226), .b(new_n256), .c(new_n245), .d(new_n255), .out0(new_n264));
  inv020aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  xnrc02aa1n02x5               g170(.a(\b[22] ), .b(\a[23] ), .out0(new_n266));
  norb02aa1n09x5               g171(.a(new_n256), .b(new_n266), .out0(new_n267));
  norp02aa1n02x5               g172(.a(\b[23] ), .b(\a[24] ), .o1(new_n268));
  aoi112aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n269));
  nanp03aa1n02x5               g174(.a(new_n248), .b(new_n255), .c(new_n256), .o1(new_n270));
  nona22aa1n02x4               g175(.a(new_n270), .b(new_n269), .c(new_n268), .out0(new_n271));
  aoi013aa1n03x5               g176(.a(new_n271), .b(new_n241), .c(new_n245), .d(new_n267), .o1(new_n272));
  aoai13aa1n04x5               g177(.a(new_n272), .b(new_n265), .c(new_n182), .d(new_n190), .o1(new_n273));
  xorb03aa1n02x5               g178(.a(new_n273), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g179(.a(\b[24] ), .b(\a[25] ), .o1(new_n275));
  tech160nm_fixorc02aa1n05x5   g180(.a(\a[25] ), .b(\b[24] ), .out0(new_n276));
  tech160nm_fixorc02aa1n04x5   g181(.a(\a[26] ), .b(\b[25] ), .out0(new_n277));
  aoi112aa1n03x4               g182(.a(new_n275), .b(new_n277), .c(new_n273), .d(new_n276), .o1(new_n278));
  inv000aa1n03x5               g183(.a(new_n275), .o1(new_n279));
  inv030aa1n02x5               g184(.a(new_n272), .o1(new_n280));
  aoai13aa1n03x5               g185(.a(new_n276), .b(new_n280), .c(new_n221), .d(new_n264), .o1(new_n281));
  aobi12aa1n03x5               g186(.a(new_n277), .b(new_n281), .c(new_n279), .out0(new_n282));
  nor002aa1n02x5               g187(.a(new_n282), .b(new_n278), .o1(\s[26] ));
  and002aa1n06x5               g188(.a(new_n277), .b(new_n276), .o(new_n284));
  nano22aa1d15x5               g189(.a(new_n251), .b(new_n284), .c(new_n267), .out0(new_n285));
  aoai13aa1n06x5               g190(.a(new_n285), .b(new_n197), .c(new_n125), .d(new_n181), .o1(new_n286));
  nano22aa1n03x7               g191(.a(new_n229), .b(new_n245), .c(new_n267), .out0(new_n287));
  oao003aa1n02x5               g192(.a(\a[26] ), .b(\b[25] ), .c(new_n279), .carry(new_n288));
  inv000aa1n02x5               g193(.a(new_n288), .o1(new_n289));
  oaoi13aa1n09x5               g194(.a(new_n289), .b(new_n284), .c(new_n287), .d(new_n271), .o1(new_n290));
  xorc02aa1n12x5               g195(.a(\a[27] ), .b(\b[26] ), .out0(new_n291));
  xnbna2aa1n03x5               g196(.a(new_n291), .b(new_n290), .c(new_n286), .out0(\s[27] ));
  norp02aa1n02x5               g197(.a(\b[26] ), .b(\a[27] ), .o1(new_n293));
  inv040aa1n03x5               g198(.a(new_n293), .o1(new_n294));
  aobi12aa1n06x5               g199(.a(new_n291), .b(new_n290), .c(new_n286), .out0(new_n295));
  xnrc02aa1n02x5               g200(.a(\b[27] ), .b(\a[28] ), .out0(new_n296));
  nano22aa1n03x7               g201(.a(new_n295), .b(new_n294), .c(new_n296), .out0(new_n297));
  aoi113aa1n02x5               g202(.a(new_n269), .b(new_n268), .c(new_n248), .d(new_n256), .e(new_n255), .o1(new_n298));
  nanp02aa1n02x5               g203(.a(new_n256), .b(new_n255), .o1(new_n299));
  nona32aa1n03x5               g204(.a(new_n241), .b(new_n299), .c(new_n235), .d(new_n233), .out0(new_n300));
  inv000aa1d42x5               g205(.a(new_n284), .o1(new_n301));
  aoai13aa1n06x5               g206(.a(new_n288), .b(new_n301), .c(new_n300), .d(new_n298), .o1(new_n302));
  aoai13aa1n03x5               g207(.a(new_n291), .b(new_n302), .c(new_n221), .d(new_n285), .o1(new_n303));
  aoi012aa1n03x5               g208(.a(new_n296), .b(new_n303), .c(new_n294), .o1(new_n304));
  nor002aa1n02x5               g209(.a(new_n304), .b(new_n297), .o1(\s[28] ));
  norb02aa1n02x5               g210(.a(new_n291), .b(new_n296), .out0(new_n306));
  aoai13aa1n03x5               g211(.a(new_n306), .b(new_n302), .c(new_n221), .d(new_n285), .o1(new_n307));
  oao003aa1n02x5               g212(.a(\a[28] ), .b(\b[27] ), .c(new_n294), .carry(new_n308));
  xnrc02aa1n02x5               g213(.a(\b[28] ), .b(\a[29] ), .out0(new_n309));
  aoi012aa1n02x7               g214(.a(new_n309), .b(new_n307), .c(new_n308), .o1(new_n310));
  aobi12aa1n02x7               g215(.a(new_n306), .b(new_n290), .c(new_n286), .out0(new_n311));
  nano22aa1n02x4               g216(.a(new_n311), .b(new_n308), .c(new_n309), .out0(new_n312));
  nor002aa1n02x5               g217(.a(new_n310), .b(new_n312), .o1(\s[29] ));
  xorb03aa1n02x5               g218(.a(new_n114), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g219(.a(new_n291), .b(new_n309), .c(new_n296), .out0(new_n315));
  aoai13aa1n03x5               g220(.a(new_n315), .b(new_n302), .c(new_n221), .d(new_n285), .o1(new_n316));
  oao003aa1n02x5               g221(.a(\a[29] ), .b(\b[28] ), .c(new_n308), .carry(new_n317));
  xnrc02aa1n02x5               g222(.a(\b[29] ), .b(\a[30] ), .out0(new_n318));
  aoi012aa1n03x5               g223(.a(new_n318), .b(new_n316), .c(new_n317), .o1(new_n319));
  aobi12aa1n02x7               g224(.a(new_n315), .b(new_n290), .c(new_n286), .out0(new_n320));
  nano22aa1n03x5               g225(.a(new_n320), .b(new_n317), .c(new_n318), .out0(new_n321));
  norp02aa1n03x5               g226(.a(new_n319), .b(new_n321), .o1(\s[30] ));
  xnrc02aa1n02x5               g227(.a(\b[30] ), .b(\a[31] ), .out0(new_n323));
  norb02aa1n02x5               g228(.a(new_n315), .b(new_n318), .out0(new_n324));
  aobi12aa1n02x7               g229(.a(new_n324), .b(new_n290), .c(new_n286), .out0(new_n325));
  oao003aa1n02x5               g230(.a(\a[30] ), .b(\b[29] ), .c(new_n317), .carry(new_n326));
  nano22aa1n03x5               g231(.a(new_n325), .b(new_n323), .c(new_n326), .out0(new_n327));
  aoai13aa1n03x5               g232(.a(new_n324), .b(new_n302), .c(new_n221), .d(new_n285), .o1(new_n328));
  aoi012aa1n02x7               g233(.a(new_n323), .b(new_n328), .c(new_n326), .o1(new_n329));
  nor002aa1n02x5               g234(.a(new_n329), .b(new_n327), .o1(\s[31] ));
  xnrb03aa1n02x5               g235(.a(new_n116), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g236(.a(\a[3] ), .b(\b[2] ), .c(new_n116), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g238(.a(new_n139), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  inv000aa1d42x5               g239(.a(\a[6] ), .o1(new_n335));
  tech160nm_fioaoi03aa1n03p5x5 g240(.a(new_n106), .b(new_n107), .c(new_n139), .o1(new_n336));
  xorb03aa1n02x5               g241(.a(new_n336), .b(\b[5] ), .c(new_n335), .out0(\s[6] ));
  inv000aa1d42x5               g242(.a(\b[5] ), .o1(new_n338));
  nanb02aa1n06x5               g243(.a(new_n122), .b(new_n336), .out0(new_n339));
  oai112aa1n03x5               g244(.a(new_n339), .b(new_n141), .c(new_n338), .d(new_n335), .o1(new_n340));
  oaoi13aa1n02x5               g245(.a(new_n141), .b(new_n339), .c(new_n335), .d(new_n338), .o1(new_n341));
  norb02aa1n02x5               g246(.a(new_n340), .b(new_n341), .out0(\s[7] ));
  xnbna2aa1n03x5               g247(.a(new_n140), .b(new_n340), .c(new_n100), .out0(\s[8] ));
  xorb03aa1n02x5               g248(.a(new_n125), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


