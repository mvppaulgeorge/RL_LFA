// Benchmark "adder" written by ABC on Thu Jul 18 07:16:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n154, new_n155, new_n156,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n192, new_n193, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n262, new_n263, new_n264, new_n265, new_n266, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n330, new_n331,
    new_n332, new_n335, new_n336, new_n337, new_n339, new_n341;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor042aa1n12x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\a[2] ), .o1(new_n99));
  inv000aa1d42x5               g004(.a(\b[1] ), .o1(new_n100));
  nand22aa1n12x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  oaoi03aa1n06x5               g006(.a(new_n99), .b(new_n100), .c(new_n101), .o1(new_n102));
  nand02aa1n04x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nor022aa1n16x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand02aa1n06x5               g009(.a(\b[3] ), .b(\a[4] ), .o1(new_n105));
  nor002aa1n20x5               g010(.a(\b[3] ), .b(\a[4] ), .o1(new_n106));
  nona23aa1n09x5               g011(.a(new_n105), .b(new_n103), .c(new_n106), .d(new_n104), .out0(new_n107));
  inv000aa1d42x5               g012(.a(\a[3] ), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\b[2] ), .o1(new_n109));
  aoai13aa1n04x5               g014(.a(new_n105), .b(new_n106), .c(new_n109), .d(new_n108), .o1(new_n110));
  oai012aa1n12x5               g015(.a(new_n110), .b(new_n107), .c(new_n102), .o1(new_n111));
  nor022aa1n04x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nanp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor002aa1d32x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand02aa1d16x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nona23aa1n03x5               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  xnrc02aa1n02x5               g021(.a(\b[6] ), .b(\a[7] ), .out0(new_n117));
  tech160nm_fixnrc02aa1n02p5x5 g022(.a(\b[4] ), .b(\a[5] ), .out0(new_n118));
  nor043aa1n03x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\a[7] ), .o1(new_n120));
  inv000aa1d42x5               g025(.a(\b[6] ), .o1(new_n121));
  nor042aa1d18x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  aoi122aa1n12x5               g027(.a(new_n114), .b(new_n121), .c(new_n120), .d(new_n122), .e(new_n115), .o1(new_n123));
  aoi022aa1n02x5               g028(.a(\b[7] ), .b(\a[8] ), .c(\a[7] ), .d(\b[6] ), .o1(new_n124));
  obai22aa1n09x5               g029(.a(new_n124), .b(new_n123), .c(\a[8] ), .d(\b[7] ), .out0(new_n125));
  nanp02aa1n04x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n97), .out0(new_n127));
  aoai13aa1n06x5               g032(.a(new_n127), .b(new_n125), .c(new_n111), .d(new_n119), .o1(new_n128));
  nor002aa1n12x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand02aa1d20x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g037(.a(new_n129), .o1(new_n133));
  inv000aa1d42x5               g038(.a(new_n130), .o1(new_n134));
  aoai13aa1n06x5               g039(.a(new_n133), .b(new_n134), .c(new_n128), .d(new_n98), .o1(new_n135));
  xorb03aa1n02x5               g040(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor042aa1n04x5               g041(.a(\b[10] ), .b(\a[11] ), .o1(new_n137));
  nand02aa1d08x5               g042(.a(\b[10] ), .b(\a[11] ), .o1(new_n138));
  nor042aa1n04x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  nanp02aa1n12x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  norb02aa1n06x4               g045(.a(new_n140), .b(new_n139), .out0(new_n141));
  aoai13aa1n04x5               g046(.a(new_n141), .b(new_n137), .c(new_n135), .d(new_n138), .o1(new_n142));
  aoi112aa1n02x7               g047(.a(new_n137), .b(new_n141), .c(new_n135), .d(new_n138), .o1(new_n143));
  norb02aa1n03x4               g048(.a(new_n142), .b(new_n143), .out0(\s[12] ));
  nano23aa1n06x5               g049(.a(new_n137), .b(new_n139), .c(new_n140), .d(new_n138), .out0(new_n145));
  nano23aa1n06x5               g050(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n126), .out0(new_n146));
  and002aa1n02x5               g051(.a(new_n146), .b(new_n145), .o(new_n147));
  aoai13aa1n03x5               g052(.a(new_n147), .b(new_n125), .c(new_n111), .d(new_n119), .o1(new_n148));
  aob012aa1n02x5               g053(.a(new_n133), .b(new_n97), .c(new_n130), .out0(new_n149));
  aoi112aa1n02x5               g054(.a(\b[10] ), .b(\a[11] ), .c(\a[12] ), .d(\b[11] ), .o1(new_n150));
  aoi112aa1n02x7               g055(.a(new_n150), .b(new_n139), .c(new_n145), .d(new_n149), .o1(new_n151));
  nanp02aa1n02x5               g056(.a(new_n148), .b(new_n151), .o1(new_n152));
  xorb03aa1n02x5               g057(.a(new_n152), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  nor042aa1d18x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand22aa1n04x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  aoi012aa1n02x5               g060(.a(new_n154), .b(new_n152), .c(new_n155), .o1(new_n156));
  xnrb03aa1n02x5               g061(.a(new_n156), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g062(.a(\b[13] ), .b(\a[14] ), .o1(new_n158));
  nand02aa1d16x5               g063(.a(\b[13] ), .b(\a[14] ), .o1(new_n159));
  nona23aa1n03x5               g064(.a(new_n159), .b(new_n155), .c(new_n154), .d(new_n158), .out0(new_n160));
  ao0012aa1n12x5               g065(.a(new_n158), .b(new_n154), .c(new_n159), .o(new_n161));
  inv000aa1d42x5               g066(.a(new_n161), .o1(new_n162));
  aoai13aa1n03x5               g067(.a(new_n162), .b(new_n160), .c(new_n148), .d(new_n151), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n06x5               g069(.a(\b[14] ), .b(\a[15] ), .o1(new_n165));
  nand42aa1d28x5               g070(.a(\b[14] ), .b(\a[15] ), .o1(new_n166));
  nor042aa1n06x5               g071(.a(\b[15] ), .b(\a[16] ), .o1(new_n167));
  nand42aa1n10x5               g072(.a(\b[15] ), .b(\a[16] ), .o1(new_n168));
  norb02aa1n03x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  aoai13aa1n03x5               g074(.a(new_n169), .b(new_n165), .c(new_n163), .d(new_n166), .o1(new_n170));
  norb02aa1n02x7               g075(.a(new_n166), .b(new_n165), .out0(new_n171));
  aoi112aa1n02x5               g076(.a(new_n165), .b(new_n169), .c(new_n163), .d(new_n171), .o1(new_n172));
  norb02aa1n03x4               g077(.a(new_n170), .b(new_n172), .out0(\s[16] ));
  nano23aa1n06x5               g078(.a(new_n154), .b(new_n158), .c(new_n159), .d(new_n155), .out0(new_n174));
  nano23aa1d15x5               g079(.a(new_n165), .b(new_n167), .c(new_n168), .d(new_n166), .out0(new_n175));
  nand02aa1d04x5               g080(.a(new_n175), .b(new_n174), .o1(new_n176));
  nano22aa1n03x7               g081(.a(new_n176), .b(new_n145), .c(new_n146), .out0(new_n177));
  aoai13aa1n12x5               g082(.a(new_n177), .b(new_n125), .c(new_n111), .d(new_n119), .o1(new_n178));
  aoi112aa1n02x7               g083(.a(\b[8] ), .b(\a[9] ), .c(\a[10] ), .d(\b[9] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n138), .b(new_n137), .out0(new_n180));
  oai112aa1n03x5               g085(.a(new_n180), .b(new_n141), .c(new_n179), .d(new_n129), .o1(new_n181));
  nona22aa1n03x5               g086(.a(new_n181), .b(new_n150), .c(new_n139), .out0(new_n182));
  nano22aa1n03x7               g087(.a(new_n160), .b(new_n171), .c(new_n169), .out0(new_n183));
  aoi112aa1n09x5               g088(.a(\b[14] ), .b(\a[15] ), .c(\a[16] ), .d(\b[15] ), .o1(new_n184));
  nand42aa1n16x5               g089(.a(new_n175), .b(new_n161), .o1(new_n185));
  nona22aa1d18x5               g090(.a(new_n185), .b(new_n184), .c(new_n167), .out0(new_n186));
  aoi012aa1d24x5               g091(.a(new_n186), .b(new_n182), .c(new_n183), .o1(new_n187));
  nor042aa1n09x5               g092(.a(\b[16] ), .b(\a[17] ), .o1(new_n188));
  nand42aa1n20x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  norb02aa1n02x5               g094(.a(new_n189), .b(new_n188), .out0(new_n190));
  xnbna2aa1n03x5               g095(.a(new_n190), .b(new_n178), .c(new_n187), .out0(\s[17] ));
  nanp02aa1n09x5               g096(.a(new_n178), .b(new_n187), .o1(new_n192));
  tech160nm_fiaoi012aa1n05x5   g097(.a(new_n188), .b(new_n192), .c(new_n190), .o1(new_n193));
  xnrb03aa1n03x5               g098(.a(new_n193), .b(\b[17] ), .c(\a[18] ), .out0(\s[18] ));
  nor022aa1n06x5               g099(.a(\b[17] ), .b(\a[18] ), .o1(new_n195));
  nand42aa1n20x5               g100(.a(\b[17] ), .b(\a[18] ), .o1(new_n196));
  nano23aa1d15x5               g101(.a(new_n188), .b(new_n195), .c(new_n196), .d(new_n189), .out0(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  oa0012aa1n02x5               g103(.a(new_n196), .b(new_n195), .c(new_n188), .o(new_n199));
  inv000aa1n02x5               g104(.a(new_n199), .o1(new_n200));
  aoai13aa1n06x5               g105(.a(new_n200), .b(new_n198), .c(new_n178), .d(new_n187), .o1(new_n201));
  xorb03aa1n02x5               g106(.a(new_n201), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g107(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv040aa1d32x5               g108(.a(\a[19] ), .o1(new_n204));
  inv000aa1d42x5               g109(.a(\b[18] ), .o1(new_n205));
  nand22aa1n12x5               g110(.a(new_n205), .b(new_n204), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  nand42aa1n04x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  nor002aa1n16x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nanp02aa1n12x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n02x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  aoai13aa1n03x5               g116(.a(new_n211), .b(new_n207), .c(new_n201), .d(new_n208), .o1(new_n212));
  aoi112aa1n02x5               g117(.a(new_n207), .b(new_n211), .c(new_n201), .d(new_n208), .o1(new_n213));
  norb02aa1n02x7               g118(.a(new_n212), .b(new_n213), .out0(\s[20] ));
  nano22aa1n12x5               g119(.a(new_n209), .b(new_n208), .c(new_n210), .out0(new_n215));
  nand23aa1n02x5               g120(.a(new_n197), .b(new_n206), .c(new_n215), .o1(new_n216));
  nanb03aa1n12x5               g121(.a(new_n209), .b(new_n210), .c(new_n208), .out0(new_n217));
  oaih22aa1n06x5               g122(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n218));
  nand23aa1n03x5               g123(.a(new_n218), .b(new_n206), .c(new_n196), .o1(new_n219));
  aoai13aa1n12x5               g124(.a(new_n210), .b(new_n209), .c(new_n204), .d(new_n205), .o1(new_n220));
  oai012aa1n18x5               g125(.a(new_n220), .b(new_n219), .c(new_n217), .o1(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  aoai13aa1n06x5               g127(.a(new_n222), .b(new_n216), .c(new_n178), .d(new_n187), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor042aa1n03x5               g129(.a(\b[20] ), .b(\a[21] ), .o1(new_n225));
  xnrc02aa1n12x5               g130(.a(\b[20] ), .b(\a[21] ), .out0(new_n226));
  inv000aa1d42x5               g131(.a(new_n226), .o1(new_n227));
  xnrc02aa1n12x5               g132(.a(\b[21] ), .b(\a[22] ), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  aoai13aa1n03x5               g134(.a(new_n229), .b(new_n225), .c(new_n223), .d(new_n227), .o1(new_n230));
  aoi112aa1n02x5               g135(.a(new_n225), .b(new_n229), .c(new_n223), .d(new_n227), .o1(new_n231));
  norb02aa1n02x7               g136(.a(new_n230), .b(new_n231), .out0(\s[22] ));
  nor042aa1d18x5               g137(.a(new_n228), .b(new_n226), .o1(new_n233));
  nona23aa1n09x5               g138(.a(new_n233), .b(new_n197), .c(new_n207), .d(new_n217), .out0(new_n234));
  inv000aa1d42x5               g139(.a(\a[22] ), .o1(new_n235));
  inv000aa1d42x5               g140(.a(\b[21] ), .o1(new_n236));
  oaoi03aa1n12x5               g141(.a(new_n235), .b(new_n236), .c(new_n225), .o1(new_n237));
  inv000aa1n02x5               g142(.a(new_n237), .o1(new_n238));
  aoi012aa1n02x5               g143(.a(new_n238), .b(new_n221), .c(new_n233), .o1(new_n239));
  aoai13aa1n06x5               g144(.a(new_n239), .b(new_n234), .c(new_n178), .d(new_n187), .o1(new_n240));
  xorb03aa1n02x5               g145(.a(new_n240), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g146(.a(\b[22] ), .b(\a[23] ), .o1(new_n242));
  xorc02aa1n12x5               g147(.a(\a[23] ), .b(\b[22] ), .out0(new_n243));
  tech160nm_fixorc02aa1n05x5   g148(.a(\a[24] ), .b(\b[23] ), .out0(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n242), .c(new_n240), .d(new_n243), .o1(new_n245));
  aoi112aa1n02x5               g150(.a(new_n242), .b(new_n244), .c(new_n240), .d(new_n243), .o1(new_n246));
  norb02aa1n03x4               g151(.a(new_n245), .b(new_n246), .out0(\s[24] ));
  inv000aa1d42x5               g152(.a(new_n233), .o1(new_n248));
  nand02aa1d04x5               g153(.a(new_n244), .b(new_n243), .o1(new_n249));
  nor043aa1n02x5               g154(.a(new_n216), .b(new_n248), .c(new_n249), .o1(new_n250));
  oai012aa1n02x5               g155(.a(new_n196), .b(\b[18] ), .c(\a[19] ), .o1(new_n251));
  oab012aa1n06x5               g156(.a(new_n251), .b(new_n188), .c(new_n195), .out0(new_n252));
  inv000aa1n02x5               g157(.a(new_n220), .o1(new_n253));
  aoai13aa1n06x5               g158(.a(new_n233), .b(new_n253), .c(new_n252), .d(new_n215), .o1(new_n254));
  orn002aa1n02x5               g159(.a(\a[23] ), .b(\b[22] ), .o(new_n255));
  oao003aa1n02x5               g160(.a(\a[24] ), .b(\b[23] ), .c(new_n255), .carry(new_n256));
  aoai13aa1n06x5               g161(.a(new_n256), .b(new_n249), .c(new_n254), .d(new_n237), .o1(new_n257));
  xorc02aa1n12x5               g162(.a(\a[25] ), .b(\b[24] ), .out0(new_n258));
  aoai13aa1n06x5               g163(.a(new_n258), .b(new_n257), .c(new_n192), .d(new_n250), .o1(new_n259));
  aoi112aa1n02x5               g164(.a(new_n258), .b(new_n257), .c(new_n192), .d(new_n250), .o1(new_n260));
  norb02aa1n03x4               g165(.a(new_n259), .b(new_n260), .out0(\s[25] ));
  nor042aa1n03x5               g166(.a(\b[24] ), .b(\a[25] ), .o1(new_n262));
  inv000aa1d42x5               g167(.a(new_n262), .o1(new_n263));
  tech160nm_fixorc02aa1n02p5x5 g168(.a(\a[26] ), .b(\b[25] ), .out0(new_n264));
  aobi12aa1n06x5               g169(.a(new_n264), .b(new_n259), .c(new_n263), .out0(new_n265));
  nona22aa1n03x5               g170(.a(new_n259), .b(new_n264), .c(new_n262), .out0(new_n266));
  norb02aa1n03x4               g171(.a(new_n266), .b(new_n265), .out0(\s[26] ));
  oao003aa1n02x5               g172(.a(new_n99), .b(new_n100), .c(new_n101), .carry(new_n268));
  nano23aa1n02x4               g173(.a(new_n106), .b(new_n104), .c(new_n103), .d(new_n105), .out0(new_n269));
  nanp02aa1n02x5               g174(.a(new_n269), .b(new_n268), .o1(new_n270));
  nano23aa1n02x5               g175(.a(new_n112), .b(new_n114), .c(new_n115), .d(new_n113), .out0(new_n271));
  nona22aa1n02x4               g176(.a(new_n271), .b(new_n117), .c(new_n118), .out0(new_n272));
  aoi012aa1n06x5               g177(.a(new_n114), .b(new_n122), .c(new_n115), .o1(new_n273));
  oaib12aa1n02x5               g178(.a(new_n273), .b(\b[6] ), .c(new_n120), .out0(new_n274));
  tech160nm_fiaoi012aa1n02p5x5 g179(.a(new_n112), .b(new_n274), .c(new_n124), .o1(new_n275));
  aoai13aa1n04x5               g180(.a(new_n275), .b(new_n272), .c(new_n270), .d(new_n110), .o1(new_n276));
  inv000aa1n02x5               g181(.a(new_n186), .o1(new_n277));
  oai012aa1n03x5               g182(.a(new_n277), .b(new_n151), .c(new_n176), .o1(new_n278));
  inv000aa1n02x5               g183(.a(new_n249), .o1(new_n279));
  nand42aa1n02x5               g184(.a(new_n264), .b(new_n258), .o1(new_n280));
  inv030aa1n02x5               g185(.a(new_n280), .o1(new_n281));
  nano22aa1n06x5               g186(.a(new_n234), .b(new_n279), .c(new_n281), .out0(new_n282));
  aoai13aa1n06x5               g187(.a(new_n282), .b(new_n278), .c(new_n276), .d(new_n177), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .c(new_n263), .carry(new_n284));
  aobi12aa1n06x5               g189(.a(new_n284), .b(new_n257), .c(new_n281), .out0(new_n285));
  xorc02aa1n12x5               g190(.a(\a[27] ), .b(\b[26] ), .out0(new_n286));
  xnbna2aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n283), .out0(\s[27] ));
  norp02aa1n02x5               g192(.a(\b[26] ), .b(\a[27] ), .o1(new_n288));
  inv040aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  nona23aa1n03x5               g194(.a(new_n281), .b(new_n233), .c(new_n216), .d(new_n249), .out0(new_n290));
  aoi012aa1n06x5               g195(.a(new_n290), .b(new_n178), .c(new_n187), .o1(new_n291));
  aoai13aa1n06x5               g196(.a(new_n279), .b(new_n238), .c(new_n221), .d(new_n233), .o1(new_n292));
  aoai13aa1n06x5               g197(.a(new_n284), .b(new_n280), .c(new_n292), .d(new_n256), .o1(new_n293));
  oaih12aa1n02x5               g198(.a(new_n286), .b(new_n293), .c(new_n291), .o1(new_n294));
  xnrc02aa1n12x5               g199(.a(\b[27] ), .b(\a[28] ), .out0(new_n295));
  aoi012aa1n02x5               g200(.a(new_n295), .b(new_n294), .c(new_n289), .o1(new_n296));
  inv000aa1d42x5               g201(.a(new_n286), .o1(new_n297));
  aoi012aa1n03x5               g202(.a(new_n297), .b(new_n285), .c(new_n283), .o1(new_n298));
  nano22aa1n03x5               g203(.a(new_n298), .b(new_n289), .c(new_n295), .out0(new_n299));
  norp02aa1n03x5               g204(.a(new_n296), .b(new_n299), .o1(\s[28] ));
  norb02aa1d21x5               g205(.a(new_n286), .b(new_n295), .out0(new_n301));
  oaih12aa1n02x5               g206(.a(new_n301), .b(new_n293), .c(new_n291), .o1(new_n302));
  oao003aa1n02x5               g207(.a(\a[28] ), .b(\b[27] ), .c(new_n289), .carry(new_n303));
  xnrc02aa1n02x5               g208(.a(\b[28] ), .b(\a[29] ), .out0(new_n304));
  aoi012aa1n02x5               g209(.a(new_n304), .b(new_n302), .c(new_n303), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n301), .o1(new_n306));
  aoi012aa1n03x5               g211(.a(new_n306), .b(new_n285), .c(new_n283), .o1(new_n307));
  nano22aa1n03x5               g212(.a(new_n307), .b(new_n303), .c(new_n304), .out0(new_n308));
  norp02aa1n03x5               g213(.a(new_n305), .b(new_n308), .o1(\s[29] ));
  xorb03aa1n02x5               g214(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n09x5               g215(.a(new_n286), .b(new_n304), .c(new_n295), .out0(new_n311));
  oaih12aa1n02x5               g216(.a(new_n311), .b(new_n293), .c(new_n291), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .c(new_n303), .carry(new_n313));
  xnrc02aa1n02x5               g218(.a(\b[29] ), .b(\a[30] ), .out0(new_n314));
  aoi012aa1n02x5               g219(.a(new_n314), .b(new_n312), .c(new_n313), .o1(new_n315));
  inv000aa1d42x5               g220(.a(new_n311), .o1(new_n316));
  aoi012aa1n03x5               g221(.a(new_n316), .b(new_n285), .c(new_n283), .o1(new_n317));
  nano22aa1n03x5               g222(.a(new_n317), .b(new_n313), .c(new_n314), .out0(new_n318));
  norp02aa1n03x5               g223(.a(new_n315), .b(new_n318), .o1(\s[30] ));
  norb02aa1n02x5               g224(.a(new_n311), .b(new_n314), .out0(new_n320));
  inv000aa1n02x5               g225(.a(new_n320), .o1(new_n321));
  aoi012aa1n03x5               g226(.a(new_n321), .b(new_n285), .c(new_n283), .o1(new_n322));
  oao003aa1n02x5               g227(.a(\a[30] ), .b(\b[29] ), .c(new_n313), .carry(new_n323));
  xnrc02aa1n02x5               g228(.a(\b[30] ), .b(\a[31] ), .out0(new_n324));
  nano22aa1n03x5               g229(.a(new_n322), .b(new_n323), .c(new_n324), .out0(new_n325));
  oaih12aa1n02x5               g230(.a(new_n320), .b(new_n293), .c(new_n291), .o1(new_n326));
  tech160nm_fiaoi012aa1n02p5x5 g231(.a(new_n324), .b(new_n326), .c(new_n323), .o1(new_n327));
  norp02aa1n03x5               g232(.a(new_n327), .b(new_n325), .o1(\s[31] ));
  xorb03aa1n02x5               g233(.a(new_n102), .b(\b[2] ), .c(new_n108), .out0(\s[3] ));
  norb02aa1n02x5               g234(.a(new_n105), .b(new_n106), .out0(new_n330));
  oaoi03aa1n02x5               g235(.a(new_n108), .b(new_n109), .c(new_n268), .o1(new_n331));
  oabi12aa1n02x5               g236(.a(new_n104), .b(new_n107), .c(new_n102), .out0(new_n332));
  mtn022aa1n02x5               g237(.a(new_n332), .b(new_n331), .sa(new_n330), .o1(\s[4] ));
  xorb03aa1n02x5               g238(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g239(.a(new_n114), .b(new_n115), .out0(new_n335));
  inv000aa1d42x5               g240(.a(new_n122), .o1(new_n336));
  nanb02aa1n02x5               g241(.a(new_n118), .b(new_n111), .out0(new_n337));
  xobna2aa1n03x5               g242(.a(new_n335), .b(new_n337), .c(new_n336), .out0(\s[6] ));
  aoai13aa1n02x5               g243(.a(new_n273), .b(new_n335), .c(new_n337), .d(new_n336), .o1(new_n339));
  xorb03aa1n02x5               g244(.a(new_n339), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g245(.a(new_n120), .b(new_n121), .c(new_n339), .o1(new_n341));
  xnrb03aa1n02x5               g246(.a(new_n341), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g247(.a(new_n276), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


