// Benchmark "adder" written by ABC on Thu Jul 18 12:16:15 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n335, new_n336, new_n337,
    new_n339, new_n340, new_n342, new_n344, new_n345, new_n346, new_n347,
    new_n349, new_n351, new_n352, new_n353, new_n355, new_n356;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[9] ), .o1(new_n97));
  nanb02aa1n02x5               g002(.a(\b[8] ), .b(new_n97), .out0(new_n98));
  and002aa1n12x5               g003(.a(\b[0] ), .b(\a[1] ), .o(new_n99));
  oaoi03aa1n09x5               g004(.a(\a[2] ), .b(\b[1] ), .c(new_n99), .o1(new_n100));
  nor042aa1n02x5               g005(.a(\b[3] ), .b(\a[4] ), .o1(new_n101));
  tech160nm_finand02aa1n03p5x5 g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  norb02aa1n06x4               g007(.a(new_n102), .b(new_n101), .out0(new_n103));
  tech160nm_finor002aa1n05x5   g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n04x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  norb02aa1n06x4               g010(.a(new_n105), .b(new_n104), .out0(new_n106));
  nanp03aa1n06x5               g011(.a(new_n100), .b(new_n103), .c(new_n106), .o1(new_n107));
  tech160nm_fiaoi012aa1n04x5   g012(.a(new_n101), .b(new_n104), .c(new_n102), .o1(new_n108));
  nand42aa1n02x5               g013(.a(new_n107), .b(new_n108), .o1(new_n109));
  oai022aa1d18x5               g014(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n110));
  aoi022aa1n09x5               g015(.a(\b[5] ), .b(\a[6] ), .c(\a[5] ), .d(\b[4] ), .o1(new_n111));
  inv040aa1d32x5               g016(.a(\a[8] ), .o1(new_n112));
  inv040aa1d32x5               g017(.a(\b[7] ), .o1(new_n113));
  oai022aa1d18x5               g018(.a(new_n112), .b(new_n113), .c(\a[7] ), .d(\b[6] ), .o1(new_n114));
  nand02aa1d28x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  oai012aa1d24x5               g020(.a(new_n115), .b(\b[7] ), .c(\a[8] ), .o1(new_n116));
  inv040aa1n04x5               g021(.a(new_n116), .o1(new_n117));
  nona23aa1d18x5               g022(.a(new_n111), .b(new_n117), .c(new_n114), .d(new_n110), .out0(new_n118));
  inv000aa1d42x5               g023(.a(new_n118), .o1(new_n119));
  nand02aa1n03x5               g024(.a(\b[5] ), .b(\a[6] ), .o1(new_n120));
  nano23aa1n06x5               g025(.a(new_n116), .b(new_n114), .c(new_n110), .d(new_n120), .out0(new_n121));
  norp02aa1n04x5               g026(.a(\b[6] ), .b(\a[7] ), .o1(new_n122));
  tech160nm_fioaoi03aa1n02p5x5 g027(.a(new_n112), .b(new_n113), .c(new_n122), .o1(new_n123));
  nanb02aa1n06x5               g028(.a(new_n121), .b(new_n123), .out0(new_n124));
  tech160nm_fixorc02aa1n03p5x5 g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n06x5               g030(.a(new_n125), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n126));
  tech160nm_fixorc02aa1n03p5x5 g031(.a(\a[10] ), .b(\b[9] ), .out0(new_n127));
  xnbna2aa1n03x5               g032(.a(new_n127), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  oa0022aa1n03x5               g033(.a(\b[9] ), .b(\a[10] ), .c(\b[8] ), .d(\a[9] ), .o(new_n129));
  nanp02aa1n02x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n06x5               g035(.a(\b[10] ), .b(\a[11] ), .o1(new_n131));
  nor042aa1n04x5               g036(.a(\b[10] ), .b(\a[11] ), .o1(new_n132));
  nanb03aa1n02x5               g037(.a(new_n132), .b(new_n130), .c(new_n131), .out0(new_n133));
  tech160nm_fiao0012aa1n02p5x5 g038(.a(new_n133), .b(new_n126), .c(new_n129), .o(new_n134));
  norb02aa1n02x5               g039(.a(new_n131), .b(new_n132), .out0(new_n135));
  aoi022aa1n02x5               g040(.a(new_n126), .b(new_n129), .c(\b[9] ), .d(\a[10] ), .o1(new_n136));
  oa0012aa1n02x5               g041(.a(new_n134), .b(new_n135), .c(new_n136), .o(\s[11] ));
  nor042aa1n04x5               g042(.a(\b[11] ), .b(\a[12] ), .o1(new_n138));
  nanp02aa1n12x5               g043(.a(\b[11] ), .b(\a[12] ), .o1(new_n139));
  norb02aa1n02x5               g044(.a(new_n139), .b(new_n138), .out0(new_n140));
  aoib12aa1n02x5               g045(.a(new_n132), .b(new_n139), .c(new_n138), .out0(new_n141));
  tech160nm_fioai012aa1n03p5x5 g046(.a(new_n134), .b(\b[10] ), .c(\a[11] ), .o1(new_n142));
  aoi022aa1n02x5               g047(.a(new_n142), .b(new_n140), .c(new_n134), .d(new_n141), .o1(\s[12] ));
  nano23aa1n03x7               g048(.a(new_n138), .b(new_n132), .c(new_n139), .d(new_n131), .out0(new_n144));
  and003aa1n02x5               g049(.a(new_n144), .b(new_n127), .c(new_n125), .o(new_n145));
  aoai13aa1n06x5               g050(.a(new_n145), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n146));
  nano22aa1n03x5               g051(.a(new_n138), .b(new_n131), .c(new_n139), .out0(new_n147));
  nona23aa1n06x5               g052(.a(new_n147), .b(new_n130), .c(new_n129), .d(new_n132), .out0(new_n148));
  aoi012aa1d24x5               g053(.a(new_n138), .b(new_n132), .c(new_n139), .o1(new_n149));
  nanp02aa1n02x5               g054(.a(new_n148), .b(new_n149), .o1(new_n150));
  nanb02aa1n02x5               g055(.a(new_n150), .b(new_n146), .out0(new_n151));
  xnrc02aa1n12x5               g056(.a(\b[12] ), .b(\a[13] ), .out0(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  and003aa1n02x5               g058(.a(new_n148), .b(new_n152), .c(new_n149), .o(new_n154));
  aoi022aa1n02x5               g059(.a(new_n151), .b(new_n153), .c(new_n146), .d(new_n154), .o1(\s[13] ));
  orn002aa1n02x5               g060(.a(\a[13] ), .b(\b[12] ), .o(new_n156));
  norb02aa1n03x5               g061(.a(new_n123), .b(new_n121), .out0(new_n157));
  aoai13aa1n06x5               g062(.a(new_n157), .b(new_n118), .c(new_n107), .d(new_n108), .o1(new_n158));
  aoai13aa1n02x5               g063(.a(new_n153), .b(new_n150), .c(new_n158), .d(new_n145), .o1(new_n159));
  xorc02aa1n12x5               g064(.a(\a[14] ), .b(\b[13] ), .out0(new_n160));
  xnbna2aa1n03x5               g065(.a(new_n160), .b(new_n159), .c(new_n156), .out0(\s[14] ));
  xnrc02aa1n02x5               g066(.a(\b[13] ), .b(\a[14] ), .out0(new_n162));
  norp02aa1n02x5               g067(.a(new_n162), .b(new_n152), .o1(new_n163));
  aoai13aa1n03x5               g068(.a(new_n163), .b(new_n150), .c(new_n158), .d(new_n145), .o1(new_n164));
  tech160nm_fioaoi03aa1n03p5x5 g069(.a(\a[14] ), .b(\b[13] ), .c(new_n156), .o1(new_n165));
  inv000aa1d42x5               g070(.a(new_n165), .o1(new_n166));
  nor002aa1d32x5               g071(.a(\b[14] ), .b(\a[15] ), .o1(new_n167));
  nand42aa1n02x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(new_n169));
  xnbna2aa1n03x5               g074(.a(new_n169), .b(new_n164), .c(new_n166), .out0(\s[15] ));
  aoai13aa1n02x5               g075(.a(new_n169), .b(new_n165), .c(new_n151), .d(new_n163), .o1(new_n171));
  xorc02aa1n12x5               g076(.a(\a[16] ), .b(\b[15] ), .out0(new_n172));
  inv040aa1d32x5               g077(.a(\a[16] ), .o1(new_n173));
  inv000aa1d42x5               g078(.a(\b[15] ), .o1(new_n174));
  nanp02aa1n02x5               g079(.a(new_n174), .b(new_n173), .o1(new_n175));
  nanp02aa1n02x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  aoi012aa1n02x5               g081(.a(new_n167), .b(new_n175), .c(new_n176), .o1(new_n177));
  inv000aa1d42x5               g082(.a(new_n167), .o1(new_n178));
  nanb02aa1n03x5               g083(.a(new_n167), .b(new_n168), .out0(new_n179));
  aoai13aa1n02x5               g084(.a(new_n178), .b(new_n179), .c(new_n164), .d(new_n166), .o1(new_n180));
  aoi022aa1n02x7               g085(.a(new_n180), .b(new_n172), .c(new_n171), .d(new_n177), .o1(\s[16] ));
  nona23aa1d18x5               g086(.a(new_n172), .b(new_n160), .c(new_n152), .d(new_n179), .out0(new_n182));
  nano32aa1d12x5               g087(.a(new_n182), .b(new_n144), .c(new_n127), .d(new_n125), .out0(new_n183));
  aoai13aa1n06x5               g088(.a(new_n183), .b(new_n124), .c(new_n109), .d(new_n119), .o1(new_n184));
  nanp03aa1n02x5               g089(.a(new_n175), .b(new_n168), .c(new_n176), .o1(new_n185));
  inv000aa1d42x5               g090(.a(\a[14] ), .o1(new_n186));
  inv000aa1d42x5               g091(.a(\b[13] ), .o1(new_n187));
  oai022aa1n02x5               g092(.a(\a[13] ), .b(\b[12] ), .c(\b[13] ), .d(\a[14] ), .o1(new_n188));
  oai122aa1n02x7               g093(.a(new_n188), .b(\a[15] ), .c(\b[14] ), .d(new_n186), .e(new_n187), .o1(new_n189));
  oaoi03aa1n02x5               g094(.a(new_n173), .b(new_n174), .c(new_n167), .o1(new_n190));
  oa0012aa1n06x5               g095(.a(new_n190), .b(new_n189), .c(new_n185), .o(new_n191));
  aoai13aa1n12x5               g096(.a(new_n191), .b(new_n182), .c(new_n148), .d(new_n149), .o1(new_n192));
  inv040aa1n08x5               g097(.a(new_n192), .o1(new_n193));
  nanp02aa1n09x5               g098(.a(new_n184), .b(new_n193), .o1(new_n194));
  xorc02aa1n02x5               g099(.a(\a[17] ), .b(\b[16] ), .out0(new_n195));
  xnrc02aa1n02x5               g100(.a(\b[16] ), .b(\a[17] ), .out0(new_n196));
  oai112aa1n02x5               g101(.a(new_n190), .b(new_n196), .c(new_n189), .d(new_n185), .o1(new_n197));
  aoib12aa1n02x5               g102(.a(new_n197), .b(new_n150), .c(new_n182), .out0(new_n198));
  aoi022aa1n02x5               g103(.a(new_n194), .b(new_n195), .c(new_n184), .d(new_n198), .o1(\s[17] ));
  nor002aa1d32x5               g104(.a(\b[16] ), .b(\a[17] ), .o1(new_n200));
  inv000aa1d42x5               g105(.a(new_n200), .o1(new_n201));
  aoai13aa1n04x5               g106(.a(new_n195), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n202));
  nor042aa1n06x5               g107(.a(\b[17] ), .b(\a[18] ), .o1(new_n203));
  nand42aa1n16x5               g108(.a(\b[17] ), .b(\a[18] ), .o1(new_n204));
  norb02aa1n03x5               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  xnbna2aa1n03x5               g110(.a(new_n205), .b(new_n202), .c(new_n201), .out0(\s[18] ));
  norb02aa1n02x5               g111(.a(new_n205), .b(new_n196), .out0(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n208));
  oaoi03aa1n02x5               g113(.a(\a[18] ), .b(\b[17] ), .c(new_n201), .o1(new_n209));
  inv000aa1d42x5               g114(.a(new_n209), .o1(new_n210));
  nor002aa1d32x5               g115(.a(\b[18] ), .b(\a[19] ), .o1(new_n211));
  nand42aa1n16x5               g116(.a(\b[18] ), .b(\a[19] ), .o1(new_n212));
  norb02aa1n12x5               g117(.a(new_n212), .b(new_n211), .out0(new_n213));
  xnbna2aa1n03x5               g118(.a(new_n213), .b(new_n208), .c(new_n210), .out0(\s[19] ));
  xnrc02aa1n02x5               g119(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  aoai13aa1n03x5               g120(.a(new_n213), .b(new_n209), .c(new_n194), .d(new_n207), .o1(new_n216));
  nor002aa1d32x5               g121(.a(\b[19] ), .b(\a[20] ), .o1(new_n217));
  nand02aa1d28x5               g122(.a(\b[19] ), .b(\a[20] ), .o1(new_n218));
  norb02aa1n02x5               g123(.a(new_n218), .b(new_n217), .out0(new_n219));
  inv000aa1d42x5               g124(.a(\a[19] ), .o1(new_n220));
  inv000aa1d42x5               g125(.a(\b[18] ), .o1(new_n221));
  aboi22aa1n03x5               g126(.a(new_n217), .b(new_n218), .c(new_n220), .d(new_n221), .out0(new_n222));
  inv020aa1n04x5               g127(.a(new_n211), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n213), .o1(new_n224));
  aoai13aa1n02x5               g129(.a(new_n223), .b(new_n224), .c(new_n208), .d(new_n210), .o1(new_n225));
  aoi022aa1n03x5               g130(.a(new_n225), .b(new_n219), .c(new_n216), .d(new_n222), .o1(\s[20] ));
  nano32aa1n03x7               g131(.a(new_n196), .b(new_n219), .c(new_n205), .d(new_n213), .out0(new_n227));
  aoai13aa1n03x5               g132(.a(new_n227), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n228));
  nanb03aa1n06x5               g133(.a(new_n217), .b(new_n218), .c(new_n212), .out0(new_n229));
  oai112aa1n06x5               g134(.a(new_n223), .b(new_n204), .c(new_n203), .d(new_n200), .o1(new_n230));
  aoi012aa1d24x5               g135(.a(new_n217), .b(new_n211), .c(new_n218), .o1(new_n231));
  oaih12aa1n12x5               g136(.a(new_n231), .b(new_n230), .c(new_n229), .o1(new_n232));
  nor002aa1d32x5               g137(.a(\b[20] ), .b(\a[21] ), .o1(new_n233));
  nand02aa1n08x5               g138(.a(\b[20] ), .b(\a[21] ), .o1(new_n234));
  norb02aa1n12x5               g139(.a(new_n234), .b(new_n233), .out0(new_n235));
  aoai13aa1n06x5               g140(.a(new_n235), .b(new_n232), .c(new_n194), .d(new_n227), .o1(new_n236));
  nano22aa1n03x7               g141(.a(new_n217), .b(new_n212), .c(new_n218), .out0(new_n237));
  tech160nm_fioai012aa1n03p5x5 g142(.a(new_n204), .b(\b[18] ), .c(\a[19] ), .o1(new_n238));
  oab012aa1n06x5               g143(.a(new_n238), .b(new_n200), .c(new_n203), .out0(new_n239));
  inv020aa1n03x5               g144(.a(new_n231), .o1(new_n240));
  aoi112aa1n02x5               g145(.a(new_n240), .b(new_n235), .c(new_n239), .d(new_n237), .o1(new_n241));
  aobi12aa1n02x7               g146(.a(new_n236), .b(new_n241), .c(new_n228), .out0(\s[21] ));
  nor042aa1n04x5               g147(.a(\b[21] ), .b(\a[22] ), .o1(new_n243));
  nand42aa1n16x5               g148(.a(\b[21] ), .b(\a[22] ), .o1(new_n244));
  norb02aa1n02x5               g149(.a(new_n244), .b(new_n243), .out0(new_n245));
  aoib12aa1n02x5               g150(.a(new_n233), .b(new_n244), .c(new_n243), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n232), .o1(new_n247));
  inv000aa1d42x5               g152(.a(new_n233), .o1(new_n248));
  inv000aa1d42x5               g153(.a(new_n235), .o1(new_n249));
  aoai13aa1n02x7               g154(.a(new_n248), .b(new_n249), .c(new_n228), .d(new_n247), .o1(new_n250));
  aoi022aa1n03x5               g155(.a(new_n250), .b(new_n245), .c(new_n236), .d(new_n246), .o1(\s[22] ));
  inv000aa1n02x5               g156(.a(new_n227), .o1(new_n252));
  nano22aa1n03x7               g157(.a(new_n252), .b(new_n235), .c(new_n245), .out0(new_n253));
  aoai13aa1n03x5               g158(.a(new_n253), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n254));
  nano23aa1d12x5               g159(.a(new_n233), .b(new_n243), .c(new_n244), .d(new_n234), .out0(new_n255));
  aoi012aa1n12x5               g160(.a(new_n243), .b(new_n233), .c(new_n244), .o1(new_n256));
  inv000aa1n02x5               g161(.a(new_n256), .o1(new_n257));
  aoi012aa1n02x5               g162(.a(new_n257), .b(new_n232), .c(new_n255), .o1(new_n258));
  inv040aa1n03x5               g163(.a(new_n258), .o1(new_n259));
  xorc02aa1n12x5               g164(.a(\a[23] ), .b(\b[22] ), .out0(new_n260));
  aoai13aa1n06x5               g165(.a(new_n260), .b(new_n259), .c(new_n194), .d(new_n253), .o1(new_n261));
  aoi112aa1n02x5               g166(.a(new_n260), .b(new_n257), .c(new_n232), .d(new_n255), .o1(new_n262));
  aobi12aa1n02x7               g167(.a(new_n261), .b(new_n262), .c(new_n254), .out0(\s[23] ));
  tech160nm_fixorc02aa1n02p5x5 g168(.a(\a[24] ), .b(\b[23] ), .out0(new_n264));
  nor042aa1n06x5               g169(.a(\b[22] ), .b(\a[23] ), .o1(new_n265));
  norp02aa1n02x5               g170(.a(new_n264), .b(new_n265), .o1(new_n266));
  inv000aa1d42x5               g171(.a(new_n265), .o1(new_n267));
  inv000aa1d42x5               g172(.a(new_n260), .o1(new_n268));
  aoai13aa1n02x7               g173(.a(new_n267), .b(new_n268), .c(new_n254), .d(new_n258), .o1(new_n269));
  aoi022aa1n02x7               g174(.a(new_n269), .b(new_n264), .c(new_n261), .d(new_n266), .o1(\s[24] ));
  and002aa1n06x5               g175(.a(new_n264), .b(new_n260), .o(new_n271));
  nano22aa1n03x7               g176(.a(new_n252), .b(new_n271), .c(new_n255), .out0(new_n272));
  aoai13aa1n03x5               g177(.a(new_n272), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n273));
  aoai13aa1n04x5               g178(.a(new_n255), .b(new_n240), .c(new_n239), .d(new_n237), .o1(new_n274));
  inv000aa1n06x5               g179(.a(new_n271), .o1(new_n275));
  oao003aa1n02x5               g180(.a(\a[24] ), .b(\b[23] ), .c(new_n267), .carry(new_n276));
  aoai13aa1n12x5               g181(.a(new_n276), .b(new_n275), .c(new_n274), .d(new_n256), .o1(new_n277));
  xorc02aa1n12x5               g182(.a(\a[25] ), .b(\b[24] ), .out0(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n277), .c(new_n194), .d(new_n272), .o1(new_n279));
  aoai13aa1n04x5               g184(.a(new_n271), .b(new_n257), .c(new_n232), .d(new_n255), .o1(new_n280));
  inv000aa1d42x5               g185(.a(new_n278), .o1(new_n281));
  and003aa1n02x5               g186(.a(new_n280), .b(new_n281), .c(new_n276), .o(new_n282));
  aobi12aa1n03x7               g187(.a(new_n279), .b(new_n282), .c(new_n273), .out0(\s[25] ));
  xorc02aa1n02x5               g188(.a(\a[26] ), .b(\b[25] ), .out0(new_n284));
  nor042aa1n03x5               g189(.a(\b[24] ), .b(\a[25] ), .o1(new_n285));
  norp02aa1n02x5               g190(.a(new_n284), .b(new_n285), .o1(new_n286));
  inv000aa1d42x5               g191(.a(new_n277), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n285), .o1(new_n288));
  aoai13aa1n02x7               g193(.a(new_n288), .b(new_n281), .c(new_n273), .d(new_n287), .o1(new_n289));
  aoi022aa1n02x7               g194(.a(new_n289), .b(new_n284), .c(new_n279), .d(new_n286), .o1(\s[26] ));
  and002aa1n02x5               g195(.a(new_n284), .b(new_n278), .o(new_n291));
  nano32aa1n03x7               g196(.a(new_n252), .b(new_n291), .c(new_n255), .d(new_n271), .out0(new_n292));
  aoai13aa1n06x5               g197(.a(new_n292), .b(new_n192), .c(new_n158), .d(new_n183), .o1(new_n293));
  inv000aa1n02x5               g198(.a(new_n291), .o1(new_n294));
  oao003aa1n02x5               g199(.a(\a[26] ), .b(\b[25] ), .c(new_n288), .carry(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n294), .c(new_n280), .d(new_n276), .o1(new_n296));
  xorc02aa1n12x5               g201(.a(\a[27] ), .b(\b[26] ), .out0(new_n297));
  aoai13aa1n06x5               g202(.a(new_n297), .b(new_n296), .c(new_n194), .d(new_n292), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n295), .o1(new_n299));
  aoi112aa1n02x5               g204(.a(new_n297), .b(new_n299), .c(new_n277), .d(new_n291), .o1(new_n300));
  aobi12aa1n02x7               g205(.a(new_n298), .b(new_n300), .c(new_n293), .out0(\s[27] ));
  tech160nm_fixorc02aa1n02p5x5 g206(.a(\a[28] ), .b(\b[27] ), .out0(new_n302));
  norp02aa1n02x5               g207(.a(\b[26] ), .b(\a[27] ), .o1(new_n303));
  norp02aa1n02x5               g208(.a(new_n302), .b(new_n303), .o1(new_n304));
  tech160nm_fiaoi012aa1n05x5   g209(.a(new_n299), .b(new_n277), .c(new_n291), .o1(new_n305));
  inv000aa1n03x5               g210(.a(new_n303), .o1(new_n306));
  inv000aa1d42x5               g211(.a(new_n297), .o1(new_n307));
  aoai13aa1n02x7               g212(.a(new_n306), .b(new_n307), .c(new_n305), .d(new_n293), .o1(new_n308));
  aoi022aa1n02x7               g213(.a(new_n308), .b(new_n302), .c(new_n298), .d(new_n304), .o1(\s[28] ));
  and002aa1n02x5               g214(.a(new_n302), .b(new_n297), .o(new_n310));
  aoai13aa1n03x5               g215(.a(new_n310), .b(new_n296), .c(new_n194), .d(new_n292), .o1(new_n311));
  inv000aa1d42x5               g216(.a(new_n310), .o1(new_n312));
  oao003aa1n02x5               g217(.a(\a[28] ), .b(\b[27] ), .c(new_n306), .carry(new_n313));
  aoai13aa1n02x7               g218(.a(new_n313), .b(new_n312), .c(new_n305), .d(new_n293), .o1(new_n314));
  xorc02aa1n02x5               g219(.a(\a[29] ), .b(\b[28] ), .out0(new_n315));
  norb02aa1n02x5               g220(.a(new_n313), .b(new_n315), .out0(new_n316));
  aoi022aa1n03x5               g221(.a(new_n314), .b(new_n315), .c(new_n311), .d(new_n316), .o1(\s[29] ));
  xnrb03aa1n02x5               g222(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g223(.a(new_n307), .b(new_n302), .c(new_n315), .out0(new_n319));
  aoai13aa1n03x5               g224(.a(new_n319), .b(new_n296), .c(new_n194), .d(new_n292), .o1(new_n320));
  inv000aa1d42x5               g225(.a(new_n319), .o1(new_n321));
  oao003aa1n02x5               g226(.a(\a[29] ), .b(\b[28] ), .c(new_n313), .carry(new_n322));
  aoai13aa1n02x7               g227(.a(new_n322), .b(new_n321), .c(new_n305), .d(new_n293), .o1(new_n323));
  xorc02aa1n02x5               g228(.a(\a[30] ), .b(\b[29] ), .out0(new_n324));
  norb02aa1n02x5               g229(.a(new_n322), .b(new_n324), .out0(new_n325));
  aoi022aa1n03x5               g230(.a(new_n323), .b(new_n324), .c(new_n320), .d(new_n325), .o1(\s[30] ));
  nano32aa1n03x7               g231(.a(new_n307), .b(new_n324), .c(new_n302), .d(new_n315), .out0(new_n327));
  aoai13aa1n03x5               g232(.a(new_n327), .b(new_n296), .c(new_n194), .d(new_n292), .o1(new_n328));
  xorc02aa1n02x5               g233(.a(\a[31] ), .b(\b[30] ), .out0(new_n329));
  oao003aa1n02x5               g234(.a(\a[30] ), .b(\b[29] ), .c(new_n322), .carry(new_n330));
  norb02aa1n02x5               g235(.a(new_n330), .b(new_n329), .out0(new_n331));
  inv000aa1d42x5               g236(.a(new_n327), .o1(new_n332));
  aoai13aa1n02x7               g237(.a(new_n330), .b(new_n332), .c(new_n305), .d(new_n293), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n333), .b(new_n329), .c(new_n328), .d(new_n331), .o1(\s[31] ));
  orn002aa1n02x5               g239(.a(\a[2] ), .b(\b[1] ), .o(new_n335));
  nanp02aa1n02x5               g240(.a(\b[1] ), .b(\a[2] ), .o1(new_n336));
  nanb03aa1n02x5               g241(.a(new_n99), .b(new_n335), .c(new_n336), .out0(new_n337));
  xnbna2aa1n03x5               g242(.a(new_n106), .b(new_n337), .c(new_n335), .out0(\s[3] ));
  aoai13aa1n02x5               g243(.a(new_n103), .b(new_n104), .c(new_n100), .d(new_n105), .o1(new_n339));
  aoi112aa1n02x5               g244(.a(new_n104), .b(new_n103), .c(new_n100), .d(new_n105), .o1(new_n340));
  norb02aa1n02x5               g245(.a(new_n339), .b(new_n340), .out0(\s[4] ));
  xorc02aa1n02x5               g246(.a(\a[5] ), .b(\b[4] ), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n342), .b(new_n107), .c(new_n108), .out0(\s[5] ));
  xorc02aa1n02x5               g248(.a(\a[6] ), .b(\b[5] ), .out0(new_n344));
  nanp02aa1n02x5               g249(.a(new_n109), .b(new_n342), .o1(new_n345));
  oa0012aa1n02x5               g250(.a(new_n345), .b(\b[4] ), .c(\a[5] ), .o(new_n346));
  nanb03aa1n06x5               g251(.a(new_n110), .b(new_n345), .c(new_n120), .out0(new_n347));
  oai012aa1n02x5               g252(.a(new_n347), .b(new_n346), .c(new_n344), .o1(\s[6] ));
  norb02aa1n02x5               g253(.a(new_n115), .b(new_n122), .out0(new_n349));
  xobna2aa1n03x5               g254(.a(new_n349), .b(new_n347), .c(new_n120), .out0(\s[7] ));
  aoi013aa1n02x4               g255(.a(new_n122), .b(new_n347), .c(new_n120), .d(new_n349), .o1(new_n351));
  xorc02aa1n02x5               g256(.a(\a[8] ), .b(\b[7] ), .out0(new_n352));
  aoi113aa1n02x5               g257(.a(new_n352), .b(new_n122), .c(new_n347), .d(new_n349), .e(new_n120), .o1(new_n353));
  aoib12aa1n03x5               g258(.a(new_n353), .b(new_n352), .c(new_n351), .out0(\s[8] ));
  nanp02aa1n02x5               g259(.a(new_n109), .b(new_n119), .o1(new_n355));
  norb03aa1n02x5               g260(.a(new_n123), .b(new_n121), .c(new_n125), .out0(new_n356));
  aoi022aa1n02x5               g261(.a(new_n158), .b(new_n125), .c(new_n355), .d(new_n356), .o1(\s[9] ));
endmodule


