// Benchmark "adder" written by ABC on Wed Jul 17 14:12:10 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n191, new_n192, new_n193, new_n194, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n208, new_n209, new_n210, new_n211, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n291, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n311, new_n312, new_n314, new_n315, new_n316, new_n317,
    new_n320, new_n321, new_n323, new_n324, new_n325;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  norp02aa1n04x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nand42aa1n06x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  norb02aa1n02x5               g003(.a(new_n98), .b(new_n97), .out0(new_n99));
  nand42aa1n06x5               g004(.a(\b[8] ), .b(\a[9] ), .o1(new_n100));
  nor042aa1n06x5               g005(.a(\b[1] ), .b(\a[2] ), .o1(new_n101));
  aoi022aa1n09x5               g006(.a(\b[1] ), .b(\a[2] ), .c(\a[1] ), .d(\b[0] ), .o1(new_n102));
  nor042aa1n03x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nanp02aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  norb02aa1n03x4               g009(.a(new_n104), .b(new_n103), .out0(new_n105));
  oai012aa1n06x5               g010(.a(new_n105), .b(new_n102), .c(new_n101), .o1(new_n106));
  oai022aa1n02x5               g011(.a(\a[3] ), .b(\b[2] ), .c(\b[3] ), .d(\a[4] ), .o1(new_n107));
  nanb02aa1n06x5               g012(.a(new_n107), .b(new_n106), .out0(new_n108));
  xnrc02aa1n02x5               g013(.a(\b[4] ), .b(\a[5] ), .out0(new_n109));
  nor002aa1d32x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n03x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  nand42aa1n04x5               g016(.a(\b[5] ), .b(\a[6] ), .o1(new_n112));
  nanb03aa1n03x5               g017(.a(new_n110), .b(new_n112), .c(new_n111), .out0(new_n113));
  norp02aa1n04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand42aa1n20x5               g019(.a(\b[7] ), .b(\a[8] ), .o1(new_n115));
  nand02aa1d08x5               g020(.a(\b[3] ), .b(\a[4] ), .o1(new_n116));
  norp02aa1n02x5               g021(.a(\b[5] ), .b(\a[6] ), .o1(new_n117));
  nona23aa1n02x4               g022(.a(new_n116), .b(new_n115), .c(new_n117), .d(new_n114), .out0(new_n118));
  nor043aa1n03x5               g023(.a(new_n118), .b(new_n113), .c(new_n109), .o1(new_n119));
  oai022aa1n04x7               g024(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n120));
  nanb03aa1n02x5               g025(.a(new_n114), .b(new_n120), .c(new_n115), .out0(new_n121));
  inv000aa1d42x5               g026(.a(new_n110), .o1(new_n122));
  oaoi03aa1n02x5               g027(.a(\a[8] ), .b(\b[7] ), .c(new_n122), .o1(new_n123));
  oabi12aa1n06x5               g028(.a(new_n123), .b(new_n121), .c(new_n113), .out0(new_n124));
  aoai13aa1n03x5               g029(.a(new_n100), .b(new_n124), .c(new_n119), .d(new_n108), .o1(new_n125));
  nor022aa1n03x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  oaoi13aa1n02x5               g031(.a(new_n107), .b(new_n105), .c(new_n102), .d(new_n101), .o1(new_n127));
  xorc02aa1n02x5               g032(.a(\a[5] ), .b(\b[4] ), .out0(new_n128));
  nano22aa1n03x7               g033(.a(new_n110), .b(new_n111), .c(new_n112), .out0(new_n129));
  inv000aa1d42x5               g034(.a(new_n115), .o1(new_n130));
  oai012aa1n02x5               g035(.a(new_n116), .b(\b[5] ), .c(\a[6] ), .o1(new_n131));
  nor003aa1n02x5               g036(.a(new_n131), .b(new_n130), .c(new_n114), .o1(new_n132));
  nanp03aa1n02x5               g037(.a(new_n132), .b(new_n128), .c(new_n129), .o1(new_n133));
  norb02aa1n02x5               g038(.a(new_n115), .b(new_n114), .out0(new_n134));
  aoi013aa1n03x5               g039(.a(new_n123), .b(new_n129), .c(new_n134), .d(new_n120), .o1(new_n135));
  oai012aa1n02x7               g040(.a(new_n135), .b(new_n133), .c(new_n127), .o1(new_n136));
  aoi012aa1n02x5               g041(.a(new_n126), .b(new_n136), .c(new_n100), .o1(new_n137));
  nona22aa1n02x4               g042(.a(new_n98), .b(new_n126), .c(new_n97), .out0(new_n138));
  obai22aa1n02x7               g043(.a(new_n125), .b(new_n138), .c(new_n137), .d(new_n99), .out0(\s[10] ));
  norb03aa1n03x4               g044(.a(new_n98), .b(new_n97), .c(new_n126), .out0(new_n140));
  aoi022aa1n02x5               g045(.a(new_n125), .b(new_n140), .c(\b[9] ), .d(\a[10] ), .o1(new_n141));
  xorb03aa1n02x5               g046(.a(new_n141), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  nor002aa1n03x5               g047(.a(\b[11] ), .b(\a[12] ), .o1(new_n143));
  nand02aa1n06x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  norb02aa1n06x4               g049(.a(new_n144), .b(new_n143), .out0(new_n145));
  nand42aa1n03x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  nor002aa1n02x5               g051(.a(\b[10] ), .b(\a[11] ), .o1(new_n147));
  aoi012aa1n03x5               g052(.a(new_n147), .b(new_n141), .c(new_n146), .o1(new_n148));
  xnrc02aa1n02x5               g053(.a(new_n148), .b(new_n145), .out0(\s[12] ));
  aoi012aa1n03x5               g054(.a(new_n124), .b(new_n119), .c(new_n108), .o1(new_n150));
  nano22aa1n03x5               g055(.a(new_n147), .b(new_n98), .c(new_n146), .out0(new_n151));
  norb03aa1n02x7               g056(.a(new_n100), .b(new_n97), .c(new_n126), .out0(new_n152));
  nanp03aa1n03x5               g057(.a(new_n151), .b(new_n152), .c(new_n145), .o1(new_n153));
  aoi022aa1n02x5               g058(.a(\b[9] ), .b(\a[10] ), .c(\a[11] ), .d(\b[10] ), .o1(new_n154));
  nona23aa1n02x4               g059(.a(new_n154), .b(new_n144), .c(new_n147), .d(new_n143), .out0(new_n155));
  aoi012aa1n02x5               g060(.a(new_n143), .b(new_n147), .c(new_n144), .o1(new_n156));
  tech160nm_fioai012aa1n05x5   g061(.a(new_n156), .b(new_n155), .c(new_n140), .o1(new_n157));
  oabi12aa1n06x5               g062(.a(new_n157), .b(new_n150), .c(new_n153), .out0(new_n158));
  xorb03aa1n02x5               g063(.a(new_n158), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  norp02aa1n04x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  nand42aa1n02x5               g065(.a(\b[12] ), .b(\a[13] ), .o1(new_n161));
  aoi012aa1n02x5               g066(.a(new_n160), .b(new_n158), .c(new_n161), .o1(new_n162));
  xnrb03aa1n02x5               g067(.a(new_n162), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor002aa1n03x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nanp02aa1n02x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  nano23aa1n06x5               g070(.a(new_n160), .b(new_n164), .c(new_n165), .d(new_n161), .out0(new_n166));
  ao0012aa1n06x5               g071(.a(new_n164), .b(new_n160), .c(new_n165), .o(new_n167));
  nor042aa1n06x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  nand42aa1n02x5               g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  norb02aa1n03x5               g074(.a(new_n169), .b(new_n168), .out0(new_n170));
  aoai13aa1n04x5               g075(.a(new_n170), .b(new_n167), .c(new_n158), .d(new_n166), .o1(new_n171));
  aoi112aa1n02x5               g076(.a(new_n170), .b(new_n167), .c(new_n158), .d(new_n166), .o1(new_n172));
  norb02aa1n02x5               g077(.a(new_n171), .b(new_n172), .out0(\s[15] ));
  inv000aa1d42x5               g078(.a(new_n168), .o1(new_n174));
  norp02aa1n04x5               g079(.a(\b[15] ), .b(\a[16] ), .o1(new_n175));
  nand42aa1n04x5               g080(.a(\b[15] ), .b(\a[16] ), .o1(new_n176));
  norb02aa1n02x5               g081(.a(new_n176), .b(new_n175), .out0(new_n177));
  aobi12aa1n06x5               g082(.a(new_n177), .b(new_n171), .c(new_n174), .out0(new_n178));
  nona22aa1n02x4               g083(.a(new_n171), .b(new_n177), .c(new_n168), .out0(new_n179));
  norb02aa1n03x4               g084(.a(new_n179), .b(new_n178), .out0(\s[16] ));
  nano23aa1n06x5               g085(.a(new_n168), .b(new_n175), .c(new_n176), .d(new_n169), .out0(new_n181));
  nano22aa1n03x7               g086(.a(new_n153), .b(new_n166), .c(new_n181), .out0(new_n182));
  aoai13aa1n06x5               g087(.a(new_n182), .b(new_n124), .c(new_n119), .d(new_n108), .o1(new_n183));
  nona23aa1n02x4               g088(.a(new_n165), .b(new_n161), .c(new_n160), .d(new_n164), .out0(new_n184));
  nano22aa1n03x5               g089(.a(new_n184), .b(new_n170), .c(new_n177), .out0(new_n185));
  aoi012aa1n02x5               g090(.a(new_n175), .b(new_n168), .c(new_n176), .o1(new_n186));
  aob012aa1n03x5               g091(.a(new_n186), .b(new_n181), .c(new_n167), .out0(new_n187));
  aoi012aa1n06x5               g092(.a(new_n187), .b(new_n157), .c(new_n185), .o1(new_n188));
  nand02aa1d08x5               g093(.a(new_n183), .b(new_n188), .o1(new_n189));
  xorb03aa1n02x5               g094(.a(new_n189), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g095(.a(\a[18] ), .o1(new_n191));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  inv000aa1d42x5               g097(.a(\b[16] ), .o1(new_n193));
  oaoi03aa1n02x5               g098(.a(new_n192), .b(new_n193), .c(new_n189), .o1(new_n194));
  xorb03aa1n02x5               g099(.a(new_n194), .b(\b[17] ), .c(new_n191), .out0(\s[18] ));
  xroi22aa1d06x4               g100(.a(new_n192), .b(\b[16] ), .c(new_n191), .d(\b[17] ), .out0(new_n196));
  nor042aa1n03x5               g101(.a(\b[17] ), .b(\a[18] ), .o1(new_n197));
  aoi112aa1n09x5               g102(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n198));
  norp02aa1n02x5               g103(.a(new_n198), .b(new_n197), .o1(new_n199));
  inv000aa1n02x5               g104(.a(new_n199), .o1(new_n200));
  nor042aa1d18x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nand02aa1d06x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  norb02aa1n12x5               g107(.a(new_n202), .b(new_n201), .out0(new_n203));
  aoai13aa1n06x5               g108(.a(new_n203), .b(new_n200), .c(new_n189), .d(new_n196), .o1(new_n204));
  aoi112aa1n02x5               g109(.a(new_n203), .b(new_n200), .c(new_n189), .d(new_n196), .o1(new_n205));
  norb02aa1n02x5               g110(.a(new_n204), .b(new_n205), .out0(\s[19] ));
  xnrc02aa1n02x5               g111(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  inv000aa1d42x5               g112(.a(new_n201), .o1(new_n208));
  nor042aa1n09x5               g113(.a(\b[19] ), .b(\a[20] ), .o1(new_n209));
  nand02aa1d28x5               g114(.a(\b[19] ), .b(\a[20] ), .o1(new_n210));
  norb02aa1n12x5               g115(.a(new_n210), .b(new_n209), .out0(new_n211));
  xnbna2aa1n03x5               g116(.a(new_n211), .b(new_n204), .c(new_n208), .out0(\s[20] ));
  nano23aa1n06x5               g117(.a(new_n201), .b(new_n209), .c(new_n210), .d(new_n202), .out0(new_n213));
  and002aa1n02x5               g118(.a(new_n196), .b(new_n213), .o(new_n214));
  oai112aa1n06x5               g119(.a(new_n203), .b(new_n211), .c(new_n198), .d(new_n197), .o1(new_n215));
  tech160nm_fiaoi012aa1n05x5   g120(.a(new_n209), .b(new_n201), .c(new_n210), .o1(new_n216));
  nanp02aa1n02x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  xorc02aa1n12x5               g122(.a(\a[21] ), .b(\b[20] ), .out0(new_n218));
  aoai13aa1n06x5               g123(.a(new_n218), .b(new_n217), .c(new_n189), .d(new_n214), .o1(new_n219));
  aoi112aa1n02x5               g124(.a(new_n218), .b(new_n217), .c(new_n189), .d(new_n214), .o1(new_n220));
  norb02aa1n02x5               g125(.a(new_n219), .b(new_n220), .out0(\s[21] ));
  nor042aa1n06x5               g126(.a(\b[20] ), .b(\a[21] ), .o1(new_n222));
  inv000aa1d42x5               g127(.a(new_n222), .o1(new_n223));
  nor002aa1d32x5               g128(.a(\b[21] ), .b(\a[22] ), .o1(new_n224));
  nand02aa1n08x5               g129(.a(\b[21] ), .b(\a[22] ), .o1(new_n225));
  nanb02aa1n12x5               g130(.a(new_n224), .b(new_n225), .out0(new_n226));
  xobna2aa1n03x5               g131(.a(new_n226), .b(new_n219), .c(new_n223), .out0(\s[22] ));
  nanb02aa1d24x5               g132(.a(new_n226), .b(new_n218), .out0(new_n228));
  tech160nm_fiaoi012aa1n03p5x5 g133(.a(new_n224), .b(new_n222), .c(new_n225), .o1(new_n229));
  aoai13aa1n12x5               g134(.a(new_n229), .b(new_n228), .c(new_n215), .d(new_n216), .o1(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  inv000aa1n02x5               g136(.a(new_n214), .o1(new_n232));
  nona22aa1n02x4               g137(.a(new_n189), .b(new_n232), .c(new_n228), .out0(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[22] ), .b(\a[23] ), .out0(new_n234));
  xobna2aa1n03x5               g139(.a(new_n234), .b(new_n233), .c(new_n231), .out0(\s[23] ));
  nor042aa1n03x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  inv000aa1d42x5               g141(.a(new_n236), .o1(new_n237));
  aoi112aa1n02x5               g142(.a(new_n228), .b(new_n232), .c(new_n183), .d(new_n188), .o1(new_n238));
  oabi12aa1n02x5               g143(.a(new_n234), .b(new_n238), .c(new_n230), .out0(new_n239));
  xnrc02aa1n02x5               g144(.a(\b[23] ), .b(\a[24] ), .out0(new_n240));
  aoi012aa1n02x7               g145(.a(new_n240), .b(new_n239), .c(new_n237), .o1(new_n241));
  aoi012aa1n03x5               g146(.a(new_n234), .b(new_n233), .c(new_n231), .o1(new_n242));
  nano22aa1n02x4               g147(.a(new_n242), .b(new_n237), .c(new_n240), .out0(new_n243));
  norp02aa1n02x5               g148(.a(new_n241), .b(new_n243), .o1(\s[24] ));
  norp02aa1n02x5               g149(.a(new_n240), .b(new_n234), .o1(new_n245));
  oaoi03aa1n02x5               g150(.a(\a[24] ), .b(\b[23] ), .c(new_n237), .o1(new_n246));
  aoi012aa1n02x7               g151(.a(new_n246), .b(new_n230), .c(new_n245), .o1(new_n247));
  nona32aa1n02x4               g152(.a(new_n218), .b(new_n240), .c(new_n234), .d(new_n226), .out0(new_n248));
  nona22aa1n09x5               g153(.a(new_n189), .b(new_n232), .c(new_n248), .out0(new_n249));
  xnrc02aa1n12x5               g154(.a(\b[24] ), .b(\a[25] ), .out0(new_n250));
  xobna2aa1n03x5               g155(.a(new_n250), .b(new_n249), .c(new_n247), .out0(\s[25] ));
  nor042aa1n03x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  inv000aa1d42x5               g157(.a(new_n252), .o1(new_n253));
  inv000aa1n03x5               g158(.a(new_n247), .o1(new_n254));
  aoi112aa1n02x5               g159(.a(new_n248), .b(new_n232), .c(new_n183), .d(new_n188), .o1(new_n255));
  oabi12aa1n03x5               g160(.a(new_n250), .b(new_n255), .c(new_n254), .out0(new_n256));
  xorc02aa1n06x5               g161(.a(\a[26] ), .b(\b[25] ), .out0(new_n257));
  aobi12aa1n03x5               g162(.a(new_n257), .b(new_n256), .c(new_n253), .out0(new_n258));
  tech160nm_fiaoi012aa1n02p5x5 g163(.a(new_n250), .b(new_n249), .c(new_n247), .o1(new_n259));
  norp03aa1n02x5               g164(.a(new_n259), .b(new_n257), .c(new_n252), .o1(new_n260));
  norp02aa1n03x5               g165(.a(new_n258), .b(new_n260), .o1(\s[26] ));
  nanp03aa1n02x5               g166(.a(new_n138), .b(new_n151), .c(new_n145), .o1(new_n262));
  nanp02aa1n02x5               g167(.a(new_n181), .b(new_n166), .o1(new_n263));
  aobi12aa1n06x5               g168(.a(new_n186), .b(new_n181), .c(new_n167), .out0(new_n264));
  aoai13aa1n02x5               g169(.a(new_n264), .b(new_n263), .c(new_n262), .d(new_n156), .o1(new_n265));
  norb02aa1n02x5               g170(.a(new_n257), .b(new_n250), .out0(new_n266));
  nano32aa1n02x4               g171(.a(new_n248), .b(new_n266), .c(new_n196), .d(new_n213), .out0(new_n267));
  aoai13aa1n04x5               g172(.a(new_n267), .b(new_n265), .c(new_n136), .d(new_n182), .o1(new_n268));
  aoai13aa1n09x5               g173(.a(new_n266), .b(new_n246), .c(new_n230), .d(new_n245), .o1(new_n269));
  oao003aa1n02x5               g174(.a(\a[26] ), .b(\b[25] ), .c(new_n253), .carry(new_n270));
  nand23aa1n06x5               g175(.a(new_n268), .b(new_n269), .c(new_n270), .o1(new_n271));
  xorb03aa1n02x5               g176(.a(new_n271), .b(\b[26] ), .c(\a[27] ), .out0(\s[27] ));
  nor042aa1d18x5               g177(.a(\b[26] ), .b(\a[27] ), .o1(new_n273));
  inv040aa1n08x5               g178(.a(new_n273), .o1(new_n274));
  nanp02aa1n02x5               g179(.a(\b[26] ), .b(\a[27] ), .o1(new_n275));
  nand02aa1n02x5               g180(.a(new_n271), .b(new_n275), .o1(new_n276));
  xorc02aa1n12x5               g181(.a(\a[28] ), .b(\b[27] ), .out0(new_n277));
  inv000aa1d42x5               g182(.a(new_n277), .o1(new_n278));
  tech160nm_fiaoi012aa1n02p5x5 g183(.a(new_n278), .b(new_n276), .c(new_n274), .o1(new_n279));
  aoi112aa1n03x4               g184(.a(new_n273), .b(new_n277), .c(new_n271), .d(new_n275), .o1(new_n280));
  nor002aa1n02x5               g185(.a(new_n279), .b(new_n280), .o1(\s[28] ));
  nano22aa1n02x4               g186(.a(new_n278), .b(new_n274), .c(new_n275), .out0(new_n282));
  nand02aa1n02x5               g187(.a(new_n271), .b(new_n282), .o1(new_n283));
  oao003aa1n12x5               g188(.a(\a[28] ), .b(\b[27] ), .c(new_n274), .carry(new_n284));
  xorc02aa1n12x5               g189(.a(\a[29] ), .b(\b[28] ), .out0(new_n285));
  inv000aa1d42x5               g190(.a(new_n285), .o1(new_n286));
  tech160nm_fiaoi012aa1n02p5x5 g191(.a(new_n286), .b(new_n283), .c(new_n284), .o1(new_n287));
  inv000aa1d42x5               g192(.a(new_n284), .o1(new_n288));
  aoi112aa1n03x4               g193(.a(new_n285), .b(new_n288), .c(new_n271), .d(new_n282), .o1(new_n289));
  nor002aa1n02x5               g194(.a(new_n287), .b(new_n289), .o1(\s[29] ));
  nanp02aa1n02x5               g195(.a(\b[0] ), .b(\a[1] ), .o1(new_n291));
  xorb03aa1n02x5               g196(.a(new_n291), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano32aa1n02x4               g197(.a(new_n286), .b(new_n277), .c(new_n275), .d(new_n274), .out0(new_n293));
  nand02aa1n02x5               g198(.a(new_n271), .b(new_n293), .o1(new_n294));
  oao003aa1n12x5               g199(.a(\a[29] ), .b(\b[28] ), .c(new_n284), .carry(new_n295));
  tech160nm_fixorc02aa1n03p5x5 g200(.a(\a[30] ), .b(\b[29] ), .out0(new_n296));
  inv000aa1d42x5               g201(.a(new_n296), .o1(new_n297));
  aoi012aa1n06x5               g202(.a(new_n297), .b(new_n294), .c(new_n295), .o1(new_n298));
  inv000aa1d42x5               g203(.a(new_n295), .o1(new_n299));
  aoi112aa1n03x4               g204(.a(new_n296), .b(new_n299), .c(new_n271), .d(new_n293), .o1(new_n300));
  nor002aa1n02x5               g205(.a(new_n298), .b(new_n300), .o1(\s[30] ));
  xnrc02aa1n02x5               g206(.a(\b[30] ), .b(\a[31] ), .out0(new_n302));
  and003aa1n02x5               g207(.a(new_n282), .b(new_n296), .c(new_n285), .o(new_n303));
  nanp02aa1n03x5               g208(.a(new_n271), .b(new_n303), .o1(new_n304));
  oaoi03aa1n09x5               g209(.a(\a[30] ), .b(\b[29] ), .c(new_n295), .o1(new_n305));
  inv000aa1d42x5               g210(.a(new_n305), .o1(new_n306));
  aoi012aa1n03x5               g211(.a(new_n302), .b(new_n304), .c(new_n306), .o1(new_n307));
  inv000aa1d42x5               g212(.a(new_n302), .o1(new_n308));
  aoi112aa1n02x5               g213(.a(new_n308), .b(new_n305), .c(new_n271), .d(new_n303), .o1(new_n309));
  nor002aa1n02x5               g214(.a(new_n307), .b(new_n309), .o1(\s[31] ));
  inv000aa1d42x5               g215(.a(new_n101), .o1(new_n311));
  nanb02aa1n02x5               g216(.a(new_n102), .b(new_n311), .out0(new_n312));
  xorb03aa1n02x5               g217(.a(new_n312), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  inv000aa1d42x5               g218(.a(\a[4] ), .o1(new_n314));
  inv000aa1d42x5               g219(.a(\b[3] ), .o1(new_n315));
  nanp02aa1n02x5               g220(.a(new_n315), .b(new_n314), .o1(new_n316));
  aoi122aa1n02x5               g221(.a(new_n103), .b(new_n316), .c(new_n116), .d(new_n312), .e(new_n104), .o1(new_n317));
  aoi013aa1n02x4               g222(.a(new_n317), .b(new_n108), .c(new_n116), .d(new_n316), .o1(\s[4] ));
  xnbna2aa1n03x5               g223(.a(new_n109), .b(new_n108), .c(new_n116), .out0(\s[5] ));
  nanp02aa1n02x5               g224(.a(\b[4] ), .b(\a[5] ), .o1(new_n320));
  aoai13aa1n02x5               g225(.a(new_n320), .b(new_n109), .c(new_n108), .d(new_n116), .o1(new_n321));
  xnrb03aa1n02x5               g226(.a(new_n321), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  nanb03aa1n02x5               g227(.a(new_n117), .b(new_n321), .c(new_n112), .out0(new_n323));
  nanp02aa1n03x5               g228(.a(new_n323), .b(new_n129), .o1(new_n324));
  aoi022aa1n02x5               g229(.a(new_n323), .b(new_n112), .c(new_n122), .d(new_n111), .o1(new_n325));
  norb02aa1n02x5               g230(.a(new_n324), .b(new_n325), .out0(\s[7] ));
  xnbna2aa1n03x5               g231(.a(new_n134), .b(new_n324), .c(new_n122), .out0(\s[8] ));
  xorb03aa1n02x5               g232(.a(new_n136), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


