// Benchmark "adder" written by ABC on Wed Jul 17 22:40:49 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n130, new_n131, new_n133, new_n134,
    new_n135, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n149,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n173, new_n174,
    new_n175, new_n176, new_n178, new_n179, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n293, new_n295, new_n297,
    new_n299, new_n300, new_n302, new_n304;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  nand42aa1n08x5               g003(.a(\b[9] ), .b(\a[10] ), .o1(new_n99));
  and002aa1n02x5               g004(.a(\b[3] ), .b(\a[4] ), .o(new_n100));
  nand22aa1n04x5               g005(.a(\b[0] ), .b(\a[1] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(\b[1] ), .b(\a[2] ), .o1(new_n102));
  nor042aa1n02x5               g007(.a(\b[1] ), .b(\a[2] ), .o1(new_n103));
  nanp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  oai112aa1n06x5               g009(.a(new_n104), .b(new_n102), .c(new_n103), .d(new_n101), .o1(new_n105));
  oa0022aa1n09x5               g010(.a(\a[4] ), .b(\b[3] ), .c(\a[3] ), .d(\b[2] ), .o(new_n106));
  nor042aa1d18x5               g011(.a(\b[6] ), .b(\a[7] ), .o1(new_n107));
  nand22aa1n06x5               g012(.a(\b[6] ), .b(\a[7] ), .o1(new_n108));
  norb02aa1n03x5               g013(.a(new_n108), .b(new_n107), .out0(new_n109));
  aoi022aa1n06x5               g014(.a(\b[7] ), .b(\a[8] ), .c(\a[6] ), .d(\b[5] ), .o1(new_n110));
  nanp02aa1n02x5               g015(.a(\b[4] ), .b(\a[5] ), .o1(new_n111));
  nand03aa1n02x5               g016(.a(new_n109), .b(new_n110), .c(new_n111), .o1(new_n112));
  aoi112aa1n09x5               g017(.a(new_n112), .b(new_n100), .c(new_n105), .d(new_n106), .o1(new_n113));
  oai022aa1n02x5               g018(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n114));
  nanp03aa1n02x5               g019(.a(new_n109), .b(new_n110), .c(new_n114), .o1(new_n115));
  inv030aa1n02x5               g020(.a(new_n107), .o1(new_n116));
  oaoi03aa1n02x5               g021(.a(\a[8] ), .b(\b[7] ), .c(new_n116), .o1(new_n117));
  nanb02aa1n12x5               g022(.a(new_n117), .b(new_n115), .out0(new_n118));
  norp02aa1n02x5               g023(.a(new_n113), .b(new_n118), .o1(new_n119));
  oaoi03aa1n02x5               g024(.a(\a[9] ), .b(\b[8] ), .c(new_n119), .o1(new_n120));
  xobna2aa1n03x5               g025(.a(new_n120), .b(new_n99), .c(new_n98), .out0(\s[10] ));
  inv000aa1d42x5               g026(.a(\b[10] ), .o1(new_n122));
  nanb02aa1n02x5               g027(.a(\a[11] ), .b(new_n122), .out0(new_n123));
  nand42aa1n08x5               g028(.a(\b[10] ), .b(\a[11] ), .o1(new_n124));
  nanp02aa1n02x5               g029(.a(new_n123), .b(new_n124), .o1(new_n125));
  xnrc02aa1n02x5               g030(.a(\b[8] ), .b(\a[9] ), .out0(new_n126));
  oabi12aa1n02x5               g031(.a(new_n126), .b(new_n113), .c(new_n118), .out0(new_n127));
  oai112aa1n02x5               g032(.a(new_n127), .b(new_n98), .c(\b[8] ), .d(\a[9] ), .o1(new_n128));
  xnbna2aa1n03x5               g033(.a(new_n125), .b(new_n128), .c(new_n99), .out0(\s[11] ));
  norp02aa1n04x5               g034(.a(\b[10] ), .b(\a[11] ), .o1(new_n130));
  aoi013aa1n02x4               g035(.a(new_n130), .b(new_n128), .c(new_n124), .d(new_n99), .o1(new_n131));
  xnrb03aa1n02x5               g036(.a(new_n131), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1n09x5               g037(.a(\b[11] ), .b(\a[12] ), .o1(new_n133));
  nand42aa1n06x5               g038(.a(\b[11] ), .b(\a[12] ), .o1(new_n134));
  nano22aa1n09x5               g039(.a(new_n133), .b(new_n124), .c(new_n134), .out0(new_n135));
  norb03aa1n09x5               g040(.a(new_n99), .b(new_n97), .c(new_n130), .out0(new_n136));
  nanb03aa1d18x5               g041(.a(new_n126), .b(new_n136), .c(new_n135), .out0(new_n137));
  inv000aa1d42x5               g042(.a(new_n137), .o1(new_n138));
  nanb03aa1n03x5               g043(.a(new_n133), .b(new_n134), .c(new_n124), .out0(new_n139));
  oai022aa1n02x7               g044(.a(\a[10] ), .b(\b[9] ), .c(\b[8] ), .d(\a[9] ), .o1(new_n140));
  nanp03aa1n02x5               g045(.a(new_n140), .b(new_n123), .c(new_n99), .o1(new_n141));
  tech160nm_fiaoi012aa1n04x5   g046(.a(new_n133), .b(new_n130), .c(new_n134), .o1(new_n142));
  oai012aa1n06x5               g047(.a(new_n142), .b(new_n141), .c(new_n139), .o1(new_n143));
  oaoi13aa1n09x5               g048(.a(new_n143), .b(new_n138), .c(new_n113), .d(new_n118), .o1(new_n144));
  nor002aa1n10x5               g049(.a(\b[12] ), .b(\a[13] ), .o1(new_n145));
  inv000aa1n02x5               g050(.a(new_n145), .o1(new_n146));
  nand42aa1n10x5               g051(.a(\b[12] ), .b(\a[13] ), .o1(new_n147));
  xnbna2aa1n03x5               g052(.a(new_n144), .b(new_n147), .c(new_n146), .out0(\s[13] ));
  oaoi03aa1n02x5               g053(.a(\a[13] ), .b(\b[12] ), .c(new_n144), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n02x5               g055(.a(\b[13] ), .b(\a[14] ), .o1(new_n151));
  nand42aa1n03x5               g056(.a(\b[13] ), .b(\a[14] ), .o1(new_n152));
  nano23aa1d12x5               g057(.a(new_n145), .b(new_n151), .c(new_n152), .d(new_n147), .out0(new_n153));
  inv000aa1d42x5               g058(.a(new_n153), .o1(new_n154));
  oaoi03aa1n02x5               g059(.a(\a[14] ), .b(\b[13] ), .c(new_n146), .o1(new_n155));
  oabi12aa1n06x5               g060(.a(new_n155), .b(new_n144), .c(new_n154), .out0(new_n156));
  xorb03aa1n02x5               g061(.a(new_n156), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n02x5               g062(.a(\b[14] ), .b(\a[15] ), .o1(new_n158));
  nanp02aa1n02x5               g063(.a(\b[14] ), .b(\a[15] ), .o1(new_n159));
  nor042aa1n02x5               g064(.a(\b[15] ), .b(\a[16] ), .o1(new_n160));
  nand42aa1n02x5               g065(.a(\b[15] ), .b(\a[16] ), .o1(new_n161));
  norb02aa1n02x5               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  aoi112aa1n02x5               g067(.a(new_n158), .b(new_n162), .c(new_n156), .d(new_n159), .o1(new_n163));
  aoai13aa1n02x5               g068(.a(new_n162), .b(new_n158), .c(new_n156), .d(new_n159), .o1(new_n164));
  norb02aa1n02x5               g069(.a(new_n164), .b(new_n163), .out0(\s[16] ));
  nano23aa1n06x5               g070(.a(new_n158), .b(new_n160), .c(new_n161), .d(new_n159), .out0(new_n166));
  nano22aa1d15x5               g071(.a(new_n137), .b(new_n153), .c(new_n166), .out0(new_n167));
  oai012aa1d24x5               g072(.a(new_n167), .b(new_n113), .c(new_n118), .o1(new_n168));
  aoai13aa1n12x5               g073(.a(new_n166), .b(new_n155), .c(new_n143), .d(new_n153), .o1(new_n169));
  aoi012aa1n09x5               g074(.a(new_n160), .b(new_n158), .c(new_n161), .o1(new_n170));
  nanp03aa1d24x5               g075(.a(new_n168), .b(new_n169), .c(new_n170), .o1(new_n171));
  xorb03aa1n02x5               g076(.a(new_n171), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g077(.a(\a[18] ), .o1(new_n173));
  inv000aa1d42x5               g078(.a(\a[17] ), .o1(new_n174));
  inv000aa1d42x5               g079(.a(\b[16] ), .o1(new_n175));
  oaoi03aa1n02x5               g080(.a(new_n174), .b(new_n175), .c(new_n171), .o1(new_n176));
  xorb03aa1n02x5               g081(.a(new_n176), .b(\b[17] ), .c(new_n173), .out0(\s[18] ));
  xroi22aa1d04x5               g082(.a(new_n174), .b(\b[16] ), .c(new_n173), .d(\b[17] ), .out0(new_n178));
  nanp02aa1n02x5               g083(.a(new_n175), .b(new_n174), .o1(new_n179));
  oaoi03aa1n02x5               g084(.a(\a[18] ), .b(\b[17] ), .c(new_n179), .o1(new_n180));
  aoi012aa1n09x5               g085(.a(new_n180), .b(new_n171), .c(new_n178), .o1(new_n181));
  nor042aa1n09x5               g086(.a(\b[18] ), .b(\a[19] ), .o1(new_n182));
  inv000aa1d42x5               g087(.a(new_n182), .o1(new_n183));
  nanp02aa1n03x5               g088(.a(\b[18] ), .b(\a[19] ), .o1(new_n184));
  xnbna2aa1n03x5               g089(.a(new_n181), .b(new_n184), .c(new_n183), .out0(\s[19] ));
  xnrc02aa1n02x5               g090(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanb02aa1n02x5               g091(.a(new_n182), .b(new_n184), .out0(new_n187));
  nor042aa1n04x5               g092(.a(new_n181), .b(new_n187), .o1(new_n188));
  norp02aa1n06x5               g093(.a(\b[19] ), .b(\a[20] ), .o1(new_n189));
  nand02aa1d04x5               g094(.a(\b[19] ), .b(\a[20] ), .o1(new_n190));
  nanb02aa1n02x5               g095(.a(new_n189), .b(new_n190), .out0(new_n191));
  nano22aa1n02x5               g096(.a(new_n188), .b(new_n183), .c(new_n191), .out0(new_n192));
  oaoi13aa1n04x5               g097(.a(new_n191), .b(new_n183), .c(new_n181), .d(new_n187), .o1(new_n193));
  norp02aa1n03x5               g098(.a(new_n193), .b(new_n192), .o1(\s[20] ));
  nona23aa1n09x5               g099(.a(new_n190), .b(new_n184), .c(new_n182), .d(new_n189), .out0(new_n195));
  norb02aa1n02x5               g100(.a(new_n178), .b(new_n195), .out0(new_n196));
  oai022aa1n02x5               g101(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n197));
  oaib12aa1n02x5               g102(.a(new_n197), .b(new_n173), .c(\b[17] ), .out0(new_n198));
  aoi012aa1n12x5               g103(.a(new_n189), .b(new_n182), .c(new_n190), .o1(new_n199));
  oai012aa1n12x5               g104(.a(new_n199), .b(new_n195), .c(new_n198), .o1(new_n200));
  aoi012aa1n09x5               g105(.a(new_n200), .b(new_n171), .c(new_n196), .o1(new_n201));
  xnrb03aa1n03x5               g106(.a(new_n201), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g107(.a(\b[20] ), .b(\a[21] ), .o1(new_n203));
  inv040aa1n03x5               g108(.a(new_n203), .o1(new_n204));
  tech160nm_fixnrc02aa1n04x5   g109(.a(\b[20] ), .b(\a[21] ), .out0(new_n205));
  nor042aa1n03x5               g110(.a(new_n201), .b(new_n205), .o1(new_n206));
  tech160nm_fixnrc02aa1n04x5   g111(.a(\b[21] ), .b(\a[22] ), .out0(new_n207));
  nano22aa1n03x7               g112(.a(new_n206), .b(new_n204), .c(new_n207), .out0(new_n208));
  oaoi13aa1n06x5               g113(.a(new_n207), .b(new_n204), .c(new_n201), .d(new_n205), .o1(new_n209));
  norp02aa1n03x5               g114(.a(new_n209), .b(new_n208), .o1(\s[22] ));
  nano23aa1n06x5               g115(.a(new_n182), .b(new_n189), .c(new_n190), .d(new_n184), .out0(new_n211));
  nor022aa1n04x5               g116(.a(new_n207), .b(new_n205), .o1(new_n212));
  and003aa1n06x5               g117(.a(new_n178), .b(new_n212), .c(new_n211), .o(new_n213));
  inv000aa1d42x5               g118(.a(new_n199), .o1(new_n214));
  aoai13aa1n06x5               g119(.a(new_n212), .b(new_n214), .c(new_n211), .d(new_n180), .o1(new_n215));
  oao003aa1n02x5               g120(.a(\a[22] ), .b(\b[21] ), .c(new_n204), .carry(new_n216));
  nanp02aa1n02x5               g121(.a(new_n215), .b(new_n216), .o1(new_n217));
  aoi012aa1n12x5               g122(.a(new_n217), .b(new_n171), .c(new_n213), .o1(new_n218));
  xnrb03aa1n03x5               g123(.a(new_n218), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g124(.a(\b[22] ), .b(\a[23] ), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n220), .o1(new_n221));
  xnrc02aa1n12x5               g126(.a(\b[22] ), .b(\a[23] ), .out0(new_n222));
  nor042aa1n03x5               g127(.a(new_n218), .b(new_n222), .o1(new_n223));
  xnrc02aa1n12x5               g128(.a(\b[23] ), .b(\a[24] ), .out0(new_n224));
  nano22aa1n03x7               g129(.a(new_n223), .b(new_n221), .c(new_n224), .out0(new_n225));
  oaoi13aa1n06x5               g130(.a(new_n224), .b(new_n221), .c(new_n218), .d(new_n222), .o1(new_n226));
  norp02aa1n03x5               g131(.a(new_n226), .b(new_n225), .o1(\s[24] ));
  nor002aa1n03x5               g132(.a(new_n224), .b(new_n222), .o1(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  nano32aa1n02x4               g134(.a(new_n229), .b(new_n178), .c(new_n212), .d(new_n211), .out0(new_n230));
  oao003aa1n02x5               g135(.a(\a[24] ), .b(\b[23] ), .c(new_n221), .carry(new_n231));
  aoai13aa1n06x5               g136(.a(new_n231), .b(new_n229), .c(new_n215), .d(new_n216), .o1(new_n232));
  aoi012aa1n02x5               g137(.a(new_n232), .b(new_n171), .c(new_n230), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[24] ), .b(\a[25] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  xnrc02aa1n03x5               g140(.a(new_n233), .b(new_n235), .out0(\s[25] ));
  nor042aa1n03x5               g141(.a(\b[24] ), .b(\a[25] ), .o1(new_n237));
  inv000aa1d42x5               g142(.a(new_n237), .o1(new_n238));
  aoai13aa1n06x5               g143(.a(new_n235), .b(new_n232), .c(new_n171), .d(new_n230), .o1(new_n239));
  xnrc02aa1n12x5               g144(.a(\b[25] ), .b(\a[26] ), .out0(new_n240));
  nanp03aa1n06x5               g145(.a(new_n239), .b(new_n238), .c(new_n240), .o1(new_n241));
  tech160nm_fiaoi012aa1n02p5x5 g146(.a(new_n240), .b(new_n239), .c(new_n238), .o1(new_n242));
  norb02aa1n03x4               g147(.a(new_n241), .b(new_n242), .out0(\s[26] ));
  nor002aa1n02x5               g148(.a(new_n240), .b(new_n234), .o1(new_n244));
  inv020aa1n02x5               g149(.a(new_n244), .o1(new_n245));
  nona32aa1n03x5               g150(.a(new_n213), .b(new_n245), .c(new_n224), .d(new_n222), .out0(new_n246));
  nanb02aa1n12x5               g151(.a(new_n246), .b(new_n171), .out0(new_n247));
  oao003aa1n02x5               g152(.a(\a[26] ), .b(\b[25] ), .c(new_n238), .carry(new_n248));
  aobi12aa1n06x5               g153(.a(new_n248), .b(new_n232), .c(new_n244), .out0(new_n249));
  xorc02aa1n12x5               g154(.a(\a[27] ), .b(\b[26] ), .out0(new_n250));
  xnbna2aa1n03x5               g155(.a(new_n250), .b(new_n247), .c(new_n249), .out0(\s[27] ));
  norp02aa1n02x5               g156(.a(\b[26] ), .b(\a[27] ), .o1(new_n252));
  inv040aa1n03x5               g157(.a(new_n252), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n250), .o1(new_n254));
  tech160nm_fiaoi012aa1n02p5x5 g159(.a(new_n254), .b(new_n247), .c(new_n249), .o1(new_n255));
  xnrc02aa1n02x5               g160(.a(\b[27] ), .b(\a[28] ), .out0(new_n256));
  nano22aa1n03x5               g161(.a(new_n255), .b(new_n253), .c(new_n256), .out0(new_n257));
  aoi013aa1n06x4               g162(.a(new_n246), .b(new_n168), .c(new_n169), .d(new_n170), .o1(new_n258));
  inv030aa1n02x5               g163(.a(new_n216), .o1(new_n259));
  aoai13aa1n04x5               g164(.a(new_n228), .b(new_n259), .c(new_n200), .d(new_n212), .o1(new_n260));
  aoai13aa1n06x5               g165(.a(new_n248), .b(new_n245), .c(new_n260), .d(new_n231), .o1(new_n261));
  oaih12aa1n02x5               g166(.a(new_n250), .b(new_n261), .c(new_n258), .o1(new_n262));
  tech160nm_fiaoi012aa1n02p5x5 g167(.a(new_n256), .b(new_n262), .c(new_n253), .o1(new_n263));
  norp02aa1n03x5               g168(.a(new_n263), .b(new_n257), .o1(\s[28] ));
  norb02aa1n02x5               g169(.a(new_n250), .b(new_n256), .out0(new_n265));
  oaih12aa1n02x5               g170(.a(new_n265), .b(new_n261), .c(new_n258), .o1(new_n266));
  oao003aa1n02x5               g171(.a(\a[28] ), .b(\b[27] ), .c(new_n253), .carry(new_n267));
  xnrc02aa1n02x5               g172(.a(\b[28] ), .b(\a[29] ), .out0(new_n268));
  tech160nm_fiaoi012aa1n02p5x5 g173(.a(new_n268), .b(new_n266), .c(new_n267), .o1(new_n269));
  inv000aa1n02x5               g174(.a(new_n265), .o1(new_n270));
  tech160nm_fiaoi012aa1n05x5   g175(.a(new_n270), .b(new_n247), .c(new_n249), .o1(new_n271));
  nano22aa1n03x5               g176(.a(new_n271), .b(new_n267), .c(new_n268), .out0(new_n272));
  norp02aa1n03x5               g177(.a(new_n269), .b(new_n272), .o1(\s[29] ));
  xorb03aa1n02x5               g178(.a(new_n101), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n06x5               g179(.a(new_n250), .b(new_n268), .c(new_n256), .out0(new_n275));
  oaih12aa1n02x5               g180(.a(new_n275), .b(new_n261), .c(new_n258), .o1(new_n276));
  oao003aa1n02x5               g181(.a(\a[29] ), .b(\b[28] ), .c(new_n267), .carry(new_n277));
  xnrc02aa1n02x5               g182(.a(\b[29] ), .b(\a[30] ), .out0(new_n278));
  tech160nm_fiaoi012aa1n02p5x5 g183(.a(new_n278), .b(new_n276), .c(new_n277), .o1(new_n279));
  inv000aa1d42x5               g184(.a(new_n275), .o1(new_n280));
  tech160nm_fiaoi012aa1n02p5x5 g185(.a(new_n280), .b(new_n247), .c(new_n249), .o1(new_n281));
  nano22aa1n03x5               g186(.a(new_n281), .b(new_n277), .c(new_n278), .out0(new_n282));
  norp02aa1n03x5               g187(.a(new_n279), .b(new_n282), .o1(\s[30] ));
  norb02aa1n02x5               g188(.a(new_n275), .b(new_n278), .out0(new_n284));
  oaih12aa1n02x5               g189(.a(new_n284), .b(new_n261), .c(new_n258), .o1(new_n285));
  oao003aa1n02x5               g190(.a(\a[30] ), .b(\b[29] ), .c(new_n277), .carry(new_n286));
  xnrc02aa1n02x5               g191(.a(\b[30] ), .b(\a[31] ), .out0(new_n287));
  tech160nm_fiaoi012aa1n02p5x5 g192(.a(new_n287), .b(new_n285), .c(new_n286), .o1(new_n288));
  inv000aa1n02x5               g193(.a(new_n284), .o1(new_n289));
  tech160nm_fiaoi012aa1n02p5x5 g194(.a(new_n289), .b(new_n247), .c(new_n249), .o1(new_n290));
  nano22aa1n03x5               g195(.a(new_n290), .b(new_n286), .c(new_n287), .out0(new_n291));
  norp02aa1n03x5               g196(.a(new_n288), .b(new_n291), .o1(\s[31] ));
  oai012aa1n02x5               g197(.a(new_n102), .b(new_n103), .c(new_n101), .o1(new_n293));
  xnrb03aa1n02x5               g198(.a(new_n293), .b(\b[2] ), .c(\a[3] ), .out0(\s[3] ));
  oaoi03aa1n02x5               g199(.a(\a[3] ), .b(\b[2] ), .c(new_n293), .o1(new_n295));
  xorb03aa1n02x5               g200(.a(new_n295), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  aoi022aa1n02x5               g201(.a(new_n105), .b(new_n106), .c(\b[3] ), .d(\a[4] ), .o1(new_n297));
  xorb03aa1n02x5               g202(.a(new_n297), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  norp02aa1n02x5               g203(.a(\b[4] ), .b(\a[5] ), .o1(new_n299));
  oai012aa1n02x5               g204(.a(new_n111), .b(new_n297), .c(new_n299), .o1(new_n300));
  xnrb03aa1n02x5               g205(.a(new_n300), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oao003aa1n02x5               g206(.a(\a[6] ), .b(\b[5] ), .c(new_n300), .carry(new_n302));
  xnbna2aa1n03x5               g207(.a(new_n302), .b(new_n116), .c(new_n108), .out0(\s[7] ));
  oaoi03aa1n02x5               g208(.a(\a[7] ), .b(\b[6] ), .c(new_n302), .o1(new_n304));
  xorb03aa1n02x5               g209(.a(new_n304), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnrb03aa1n02x5               g210(.a(new_n119), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


