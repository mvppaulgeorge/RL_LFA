// Benchmark "adder" written by ABC on Wed Jul 17 16:44:21 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n326, new_n327, new_n330, new_n332, new_n334, new_n335,
    new_n336;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n16x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\a[2] ), .o1(new_n98));
  inv000aa1d42x5               g003(.a(\b[1] ), .o1(new_n99));
  nand02aa1d12x5               g004(.a(\b[0] ), .b(\a[1] ), .o1(new_n100));
  oao003aa1n03x5               g005(.a(new_n98), .b(new_n99), .c(new_n100), .carry(new_n101));
  norp02aa1n06x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nand42aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  norb02aa1n06x4               g008(.a(new_n103), .b(new_n102), .out0(new_n104));
  tech160nm_fixorc02aa1n05x5   g009(.a(\a[3] ), .b(\b[2] ), .out0(new_n105));
  nanp03aa1n02x5               g010(.a(new_n101), .b(new_n104), .c(new_n105), .o1(new_n106));
  inv000aa1d42x5               g011(.a(\a[3] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[2] ), .o1(new_n108));
  aoai13aa1n04x5               g013(.a(new_n103), .b(new_n102), .c(new_n107), .d(new_n108), .o1(new_n109));
  tech160nm_fixnrc02aa1n05x5   g014(.a(\b[5] ), .b(\a[6] ), .out0(new_n110));
  xorc02aa1n12x5               g015(.a(\a[5] ), .b(\b[4] ), .out0(new_n111));
  xorc02aa1n12x5               g016(.a(\a[8] ), .b(\b[7] ), .out0(new_n112));
  tech160nm_fixnrc02aa1n05x5   g017(.a(\b[6] ), .b(\a[7] ), .out0(new_n113));
  nona23aa1n03x5               g018(.a(new_n112), .b(new_n111), .c(new_n113), .d(new_n110), .out0(new_n114));
  xorc02aa1n12x5               g019(.a(\a[7] ), .b(\b[6] ), .out0(new_n115));
  inv000aa1d42x5               g020(.a(\a[6] ), .o1(new_n116));
  inv000aa1d42x5               g021(.a(\b[5] ), .o1(new_n117));
  nor042aa1n06x5               g022(.a(\b[4] ), .b(\a[5] ), .o1(new_n118));
  oao003aa1n03x5               g023(.a(new_n116), .b(new_n117), .c(new_n118), .carry(new_n119));
  inv000aa1d42x5               g024(.a(\a[7] ), .o1(new_n120));
  nanb02aa1n03x5               g025(.a(\b[6] ), .b(new_n120), .out0(new_n121));
  oaoi03aa1n02x5               g026(.a(\a[8] ), .b(\b[7] ), .c(new_n121), .o1(new_n122));
  aoi013aa1n06x4               g027(.a(new_n122), .b(new_n119), .c(new_n115), .d(new_n112), .o1(new_n123));
  aoai13aa1n12x5               g028(.a(new_n123), .b(new_n114), .c(new_n106), .d(new_n109), .o1(new_n124));
  tech160nm_fixorc02aa1n02p5x5 g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoi012aa1n02x5               g030(.a(new_n97), .b(new_n124), .c(new_n125), .o1(new_n126));
  nor042aa1n06x5               g031(.a(\b[9] ), .b(\a[10] ), .o1(new_n127));
  and002aa1n24x5               g032(.a(\b[9] ), .b(\a[10] ), .o(new_n128));
  nor042aa1n04x5               g033(.a(new_n128), .b(new_n127), .o1(new_n129));
  oaoi03aa1n02x5               g034(.a(new_n98), .b(new_n99), .c(new_n100), .o1(new_n130));
  nand02aa1n02x5               g035(.a(new_n105), .b(new_n104), .o1(new_n131));
  tech160nm_fioai012aa1n05x5   g036(.a(new_n109), .b(new_n131), .c(new_n130), .o1(new_n132));
  nano32aa1n03x7               g037(.a(new_n110), .b(new_n115), .c(new_n111), .d(new_n112), .out0(new_n133));
  nanp03aa1n02x5               g038(.a(new_n119), .b(new_n112), .c(new_n115), .o1(new_n134));
  nanb02aa1n06x5               g039(.a(new_n122), .b(new_n134), .out0(new_n135));
  aoai13aa1n02x5               g040(.a(new_n125), .b(new_n135), .c(new_n132), .d(new_n133), .o1(new_n136));
  nor022aa1n04x5               g041(.a(new_n127), .b(new_n97), .o1(new_n137));
  inv030aa1n02x5               g042(.a(new_n137), .o1(new_n138));
  nona22aa1n02x4               g043(.a(new_n136), .b(new_n128), .c(new_n138), .out0(new_n139));
  oai012aa1n02x5               g044(.a(new_n139), .b(new_n126), .c(new_n129), .o1(\s[10] ));
  nanp02aa1n03x5               g045(.a(new_n136), .b(new_n137), .o1(new_n141));
  nand02aa1d08x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nor002aa1d32x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  inv000aa1n02x5               g048(.a(new_n143), .o1(new_n144));
  nanb03aa1n02x5               g049(.a(new_n128), .b(new_n144), .c(new_n142), .out0(new_n145));
  nanb02aa1n12x5               g050(.a(new_n143), .b(new_n142), .out0(new_n146));
  inv000aa1d42x5               g051(.a(new_n128), .o1(new_n147));
  aoai13aa1n02x5               g052(.a(new_n147), .b(new_n138), .c(new_n124), .d(new_n125), .o1(new_n148));
  aboi22aa1n03x5               g053(.a(new_n145), .b(new_n141), .c(new_n148), .d(new_n146), .out0(\s[11] ));
  xorc02aa1n12x5               g054(.a(\a[12] ), .b(\b[11] ), .out0(new_n150));
  aoi113aa1n02x5               g055(.a(new_n150), .b(new_n143), .c(new_n141), .d(new_n142), .e(new_n147), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n144), .b(new_n145), .c(new_n136), .d(new_n137), .o1(new_n152));
  tech160nm_fiaoi012aa1n02p5x5 g057(.a(new_n151), .b(new_n150), .c(new_n152), .o1(\s[12] ));
  nand22aa1n03x5               g058(.a(new_n125), .b(new_n129), .o1(new_n154));
  nano32aa1n02x5               g059(.a(new_n154), .b(new_n150), .c(new_n144), .d(new_n142), .out0(new_n155));
  aoai13aa1n06x5               g060(.a(new_n155), .b(new_n135), .c(new_n132), .d(new_n133), .o1(new_n156));
  oao003aa1n02x5               g061(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .carry(new_n157));
  nona23aa1n06x5               g062(.a(new_n138), .b(new_n150), .c(new_n146), .d(new_n128), .out0(new_n158));
  nanp02aa1n02x5               g063(.a(new_n158), .b(new_n157), .o1(new_n159));
  nanb02aa1n02x5               g064(.a(new_n159), .b(new_n156), .out0(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  tech160nm_ficinv00aa1n08x5   g066(.clk(\a[13] ), .clkout(new_n162));
  nanb02aa1n12x5               g067(.a(\b[12] ), .b(new_n162), .out0(new_n163));
  xorc02aa1n02x5               g068(.a(\a[13] ), .b(\b[12] ), .out0(new_n164));
  aoai13aa1n03x5               g069(.a(new_n164), .b(new_n159), .c(new_n124), .d(new_n155), .o1(new_n165));
  xorc02aa1n02x5               g070(.a(\a[14] ), .b(\b[13] ), .out0(new_n166));
  xnbna2aa1n03x5               g071(.a(new_n166), .b(new_n165), .c(new_n163), .out0(\s[14] ));
  inv040aa1d32x5               g072(.a(\a[14] ), .o1(new_n168));
  xroi22aa1d06x4               g073(.a(new_n162), .b(\b[12] ), .c(new_n168), .d(\b[13] ), .out0(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n159), .c(new_n124), .d(new_n155), .o1(new_n170));
  oaoi03aa1n12x5               g075(.a(\a[14] ), .b(\b[13] ), .c(new_n163), .o1(new_n171));
  inv000aa1d42x5               g076(.a(new_n171), .o1(new_n172));
  xnrc02aa1n12x5               g077(.a(\b[14] ), .b(\a[15] ), .out0(new_n173));
  inv000aa1d42x5               g078(.a(new_n173), .o1(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n170), .c(new_n172), .out0(\s[15] ));
  aoai13aa1n02x5               g080(.a(new_n174), .b(new_n171), .c(new_n160), .d(new_n169), .o1(new_n176));
  xnrc02aa1n12x5               g081(.a(\b[15] ), .b(\a[16] ), .out0(new_n177));
  inv000aa1d42x5               g082(.a(new_n177), .o1(new_n178));
  nor042aa1n09x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  norb02aa1n02x5               g084(.a(new_n177), .b(new_n179), .out0(new_n180));
  inv000aa1d42x5               g085(.a(new_n179), .o1(new_n181));
  aoai13aa1n02x5               g086(.a(new_n181), .b(new_n173), .c(new_n170), .d(new_n172), .o1(new_n182));
  aoi022aa1n03x5               g087(.a(new_n182), .b(new_n178), .c(new_n176), .d(new_n180), .o1(\s[16] ));
  aoi012aa1n09x5               g088(.a(new_n135), .b(new_n132), .c(new_n133), .o1(new_n184));
  nanb02aa1n02x5               g089(.a(new_n146), .b(new_n150), .out0(new_n185));
  nor042aa1n06x5               g090(.a(new_n177), .b(new_n173), .o1(new_n186));
  nona23aa1n06x5               g091(.a(new_n186), .b(new_n169), .c(new_n185), .d(new_n154), .out0(new_n187));
  nand02aa1d04x5               g092(.a(new_n169), .b(new_n186), .o1(new_n188));
  oaoi03aa1n02x5               g093(.a(\a[16] ), .b(\b[15] ), .c(new_n181), .o1(new_n189));
  aoi012aa1n06x5               g094(.a(new_n189), .b(new_n186), .c(new_n171), .o1(new_n190));
  aoai13aa1n12x5               g095(.a(new_n190), .b(new_n188), .c(new_n158), .d(new_n157), .o1(new_n191));
  oabi12aa1n18x5               g096(.a(new_n191), .b(new_n184), .c(new_n187), .out0(new_n192));
  xorb03aa1n02x5               g097(.a(new_n192), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv040aa1d32x5               g098(.a(\a[17] ), .o1(new_n194));
  inv040aa1d28x5               g099(.a(\b[16] ), .o1(new_n195));
  nanp02aa1n02x5               g100(.a(new_n195), .b(new_n194), .o1(new_n196));
  nor043aa1n06x5               g101(.a(new_n188), .b(new_n154), .c(new_n185), .o1(new_n197));
  tech160nm_fixorc02aa1n05x5   g102(.a(\a[17] ), .b(\b[16] ), .out0(new_n198));
  aoai13aa1n03x5               g103(.a(new_n198), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n199));
  nor042aa1n04x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  nand22aa1n06x5               g105(.a(\b[17] ), .b(\a[18] ), .o1(new_n201));
  norb02aa1n06x5               g106(.a(new_n201), .b(new_n200), .out0(new_n202));
  xnbna2aa1n03x5               g107(.a(new_n202), .b(new_n199), .c(new_n196), .out0(\s[18] ));
  and002aa1n02x5               g108(.a(new_n198), .b(new_n202), .o(new_n204));
  aoai13aa1n03x5               g109(.a(new_n204), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n205));
  aoi013aa1n09x5               g110(.a(new_n200), .b(new_n201), .c(new_n194), .d(new_n195), .o1(new_n206));
  nor002aa1d32x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nanp02aa1n06x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n06x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n205), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  oaoi03aa1n03x5               g116(.a(\a[18] ), .b(\b[17] ), .c(new_n196), .o1(new_n212));
  aoai13aa1n03x5               g117(.a(new_n209), .b(new_n212), .c(new_n192), .d(new_n204), .o1(new_n213));
  nor002aa1d32x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nanp02aa1n06x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  aoib12aa1n02x5               g121(.a(new_n207), .b(new_n215), .c(new_n214), .out0(new_n217));
  inv040aa1n03x5               g122(.a(new_n207), .o1(new_n218));
  inv000aa1d42x5               g123(.a(new_n209), .o1(new_n219));
  aoai13aa1n03x5               g124(.a(new_n218), .b(new_n219), .c(new_n205), .d(new_n206), .o1(new_n220));
  aoi022aa1n03x5               g125(.a(new_n220), .b(new_n216), .c(new_n213), .d(new_n217), .o1(\s[20] ));
  nano23aa1n06x5               g126(.a(new_n207), .b(new_n214), .c(new_n215), .d(new_n208), .out0(new_n222));
  nand23aa1n06x5               g127(.a(new_n222), .b(new_n198), .c(new_n202), .o1(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n06x5               g129(.a(new_n224), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n225));
  nona23aa1n09x5               g130(.a(new_n215), .b(new_n208), .c(new_n207), .d(new_n214), .out0(new_n226));
  oaoi03aa1n09x5               g131(.a(\a[20] ), .b(\b[19] ), .c(new_n218), .o1(new_n227));
  oabi12aa1n18x5               g132(.a(new_n227), .b(new_n226), .c(new_n206), .out0(new_n228));
  inv000aa1d42x5               g133(.a(new_n228), .o1(new_n229));
  xnrc02aa1n12x5               g134(.a(\b[20] ), .b(\a[21] ), .out0(new_n230));
  inv000aa1d42x5               g135(.a(new_n230), .o1(new_n231));
  xnbna2aa1n03x5               g136(.a(new_n231), .b(new_n225), .c(new_n229), .out0(\s[21] ));
  aoai13aa1n06x5               g137(.a(new_n231), .b(new_n228), .c(new_n192), .d(new_n224), .o1(new_n233));
  xnrc02aa1n12x5               g138(.a(\b[21] ), .b(\a[22] ), .out0(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  nor042aa1n04x5               g140(.a(\b[20] ), .b(\a[21] ), .o1(new_n236));
  norb02aa1n02x5               g141(.a(new_n234), .b(new_n236), .out0(new_n237));
  inv040aa1n03x5               g142(.a(new_n236), .o1(new_n238));
  aoai13aa1n03x5               g143(.a(new_n238), .b(new_n230), .c(new_n225), .d(new_n229), .o1(new_n239));
  aoi022aa1n03x5               g144(.a(new_n239), .b(new_n235), .c(new_n233), .d(new_n237), .o1(\s[22] ));
  nor042aa1n06x5               g145(.a(new_n234), .b(new_n230), .o1(new_n241));
  norb02aa1n02x7               g146(.a(new_n241), .b(new_n223), .out0(new_n242));
  aoai13aa1n03x5               g147(.a(new_n242), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n243));
  oaoi03aa1n03x5               g148(.a(\a[22] ), .b(\b[21] ), .c(new_n238), .o1(new_n244));
  aoi012aa1n09x5               g149(.a(new_n244), .b(new_n228), .c(new_n241), .o1(new_n245));
  xnrc02aa1n12x5               g150(.a(\b[22] ), .b(\a[23] ), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n246), .o1(new_n247));
  xnbna2aa1n03x5               g152(.a(new_n247), .b(new_n243), .c(new_n245), .out0(\s[23] ));
  inv000aa1d42x5               g153(.a(new_n245), .o1(new_n249));
  aoai13aa1n03x5               g154(.a(new_n247), .b(new_n249), .c(new_n192), .d(new_n242), .o1(new_n250));
  xorc02aa1n12x5               g155(.a(\a[24] ), .b(\b[23] ), .out0(new_n251));
  nor042aa1n09x5               g156(.a(\b[22] ), .b(\a[23] ), .o1(new_n252));
  norp02aa1n02x5               g157(.a(new_n251), .b(new_n252), .o1(new_n253));
  inv000aa1d42x5               g158(.a(new_n252), .o1(new_n254));
  aoai13aa1n03x5               g159(.a(new_n254), .b(new_n246), .c(new_n243), .d(new_n245), .o1(new_n255));
  aoi022aa1n03x5               g160(.a(new_n255), .b(new_n251), .c(new_n250), .d(new_n253), .o1(\s[24] ));
  nano32aa1n02x5               g161(.a(new_n223), .b(new_n251), .c(new_n241), .d(new_n247), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n258));
  aoai13aa1n06x5               g163(.a(new_n241), .b(new_n227), .c(new_n222), .d(new_n212), .o1(new_n259));
  inv000aa1n02x5               g164(.a(new_n244), .o1(new_n260));
  norb02aa1n02x7               g165(.a(new_n251), .b(new_n246), .out0(new_n261));
  inv000aa1n02x5               g166(.a(new_n261), .o1(new_n262));
  oao003aa1n02x5               g167(.a(\a[24] ), .b(\b[23] ), .c(new_n254), .carry(new_n263));
  aoai13aa1n12x5               g168(.a(new_n263), .b(new_n262), .c(new_n259), .d(new_n260), .o1(new_n264));
  inv000aa1n02x5               g169(.a(new_n264), .o1(new_n265));
  xorc02aa1n12x5               g170(.a(\a[25] ), .b(\b[24] ), .out0(new_n266));
  xnbna2aa1n03x5               g171(.a(new_n266), .b(new_n258), .c(new_n265), .out0(\s[25] ));
  aoai13aa1n03x5               g172(.a(new_n266), .b(new_n264), .c(new_n192), .d(new_n257), .o1(new_n268));
  tech160nm_fixorc02aa1n02p5x5 g173(.a(\a[26] ), .b(\b[25] ), .out0(new_n269));
  norp02aa1n02x5               g174(.a(\b[24] ), .b(\a[25] ), .o1(new_n270));
  norp02aa1n02x5               g175(.a(new_n269), .b(new_n270), .o1(new_n271));
  inv000aa1d42x5               g176(.a(new_n270), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n266), .o1(new_n273));
  aoai13aa1n02x5               g178(.a(new_n272), .b(new_n273), .c(new_n258), .d(new_n265), .o1(new_n274));
  aoi022aa1n03x5               g179(.a(new_n274), .b(new_n269), .c(new_n268), .d(new_n271), .o1(\s[26] ));
  and002aa1n12x5               g180(.a(new_n269), .b(new_n266), .o(new_n276));
  nano32aa1n03x7               g181(.a(new_n223), .b(new_n276), .c(new_n241), .d(new_n261), .out0(new_n277));
  aoai13aa1n06x5               g182(.a(new_n277), .b(new_n191), .c(new_n124), .d(new_n197), .o1(new_n278));
  nanp02aa1n02x5               g183(.a(\b[25] ), .b(\a[26] ), .o1(new_n279));
  oai022aa1n02x5               g184(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n280));
  aoi022aa1n09x5               g185(.a(new_n264), .b(new_n276), .c(new_n279), .d(new_n280), .o1(new_n281));
  xorc02aa1n12x5               g186(.a(\a[27] ), .b(\b[26] ), .out0(new_n282));
  xnbna2aa1n03x5               g187(.a(new_n282), .b(new_n281), .c(new_n278), .out0(\s[27] ));
  aoai13aa1n03x5               g188(.a(new_n261), .b(new_n244), .c(new_n228), .d(new_n241), .o1(new_n284));
  inv000aa1n02x5               g189(.a(new_n276), .o1(new_n285));
  nanp02aa1n02x5               g190(.a(new_n280), .b(new_n279), .o1(new_n286));
  aoai13aa1n03x5               g191(.a(new_n286), .b(new_n285), .c(new_n284), .d(new_n263), .o1(new_n287));
  aoai13aa1n02x7               g192(.a(new_n282), .b(new_n287), .c(new_n192), .d(new_n277), .o1(new_n288));
  tech160nm_fixorc02aa1n02p5x5 g193(.a(\a[28] ), .b(\b[27] ), .out0(new_n289));
  nor042aa1n03x5               g194(.a(\b[26] ), .b(\a[27] ), .o1(new_n290));
  norp02aa1n02x5               g195(.a(new_n289), .b(new_n290), .o1(new_n291));
  inv000aa1n06x5               g196(.a(new_n290), .o1(new_n292));
  inv000aa1d42x5               g197(.a(new_n282), .o1(new_n293));
  aoai13aa1n03x5               g198(.a(new_n292), .b(new_n293), .c(new_n281), .d(new_n278), .o1(new_n294));
  aoi022aa1n03x5               g199(.a(new_n294), .b(new_n289), .c(new_n288), .d(new_n291), .o1(\s[28] ));
  and002aa1n02x5               g200(.a(new_n289), .b(new_n282), .o(new_n296));
  aoai13aa1n02x7               g201(.a(new_n296), .b(new_n287), .c(new_n192), .d(new_n277), .o1(new_n297));
  inv000aa1d42x5               g202(.a(new_n296), .o1(new_n298));
  oaoi03aa1n12x5               g203(.a(\a[28] ), .b(\b[27] ), .c(new_n292), .o1(new_n299));
  inv000aa1d42x5               g204(.a(new_n299), .o1(new_n300));
  aoai13aa1n03x5               g205(.a(new_n300), .b(new_n298), .c(new_n281), .d(new_n278), .o1(new_n301));
  tech160nm_fixorc02aa1n04x5   g206(.a(\a[29] ), .b(\b[28] ), .out0(new_n302));
  norp02aa1n02x5               g207(.a(new_n299), .b(new_n302), .o1(new_n303));
  aoi022aa1n03x5               g208(.a(new_n301), .b(new_n302), .c(new_n297), .d(new_n303), .o1(\s[29] ));
  xorb03aa1n02x5               g209(.a(new_n100), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x5               g210(.a(new_n293), .b(new_n289), .c(new_n302), .out0(new_n306));
  aoai13aa1n02x7               g211(.a(new_n306), .b(new_n287), .c(new_n192), .d(new_n277), .o1(new_n307));
  inv000aa1n02x5               g212(.a(new_n306), .o1(new_n308));
  inv000aa1d42x5               g213(.a(\a[29] ), .o1(new_n309));
  inv000aa1d42x5               g214(.a(\b[28] ), .o1(new_n310));
  tech160nm_fioaoi03aa1n03p5x5 g215(.a(new_n309), .b(new_n310), .c(new_n299), .o1(new_n311));
  aoai13aa1n03x5               g216(.a(new_n311), .b(new_n308), .c(new_n281), .d(new_n278), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[30] ), .b(\b[29] ), .out0(new_n313));
  oabi12aa1n02x5               g218(.a(new_n313), .b(\a[29] ), .c(\b[28] ), .out0(new_n314));
  oaoi13aa1n02x5               g219(.a(new_n314), .b(new_n299), .c(new_n309), .d(new_n310), .o1(new_n315));
  aoi022aa1n03x5               g220(.a(new_n312), .b(new_n313), .c(new_n307), .d(new_n315), .o1(\s[30] ));
  nano32aa1d12x5               g221(.a(new_n293), .b(new_n313), .c(new_n289), .d(new_n302), .out0(new_n317));
  aoai13aa1n02x7               g222(.a(new_n317), .b(new_n287), .c(new_n192), .d(new_n277), .o1(new_n318));
  xorc02aa1n02x5               g223(.a(\a[31] ), .b(\b[30] ), .out0(new_n319));
  oao003aa1n02x5               g224(.a(\a[30] ), .b(\b[29] ), .c(new_n311), .carry(new_n320));
  norb02aa1n02x5               g225(.a(new_n320), .b(new_n319), .out0(new_n321));
  inv000aa1d42x5               g226(.a(new_n317), .o1(new_n322));
  aoai13aa1n03x5               g227(.a(new_n320), .b(new_n322), .c(new_n281), .d(new_n278), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n323), .b(new_n319), .c(new_n318), .d(new_n321), .o1(\s[31] ));
  xorb03aa1n02x5               g229(.a(new_n130), .b(\b[2] ), .c(new_n107), .out0(\s[3] ));
  obai22aa1n02x7               g230(.a(new_n103), .b(new_n102), .c(\a[3] ), .d(\b[2] ), .out0(new_n326));
  aoi012aa1n02x5               g231(.a(new_n326), .b(new_n101), .c(new_n105), .o1(new_n327));
  oaoi13aa1n02x5               g232(.a(new_n327), .b(new_n132), .c(\a[4] ), .d(\b[3] ), .o1(\s[4] ));
  xnbna2aa1n03x5               g233(.a(new_n111), .b(new_n106), .c(new_n109), .out0(\s[5] ));
  tech160nm_fiao0012aa1n02p5x5 g234(.a(new_n118), .b(new_n132), .c(new_n111), .o(new_n330));
  xorb03aa1n02x5               g235(.a(new_n330), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  oaoi03aa1n03x5               g236(.a(new_n116), .b(new_n117), .c(new_n330), .o1(new_n332));
  xorb03aa1n02x5               g237(.a(new_n332), .b(\b[6] ), .c(new_n120), .out0(\s[7] ));
  nanb02aa1n02x5               g238(.a(new_n332), .b(new_n115), .out0(new_n334));
  oaoi03aa1n02x5               g239(.a(\a[7] ), .b(\b[6] ), .c(new_n332), .o1(new_n335));
  norb02aa1n02x5               g240(.a(new_n121), .b(new_n112), .out0(new_n336));
  aoi022aa1n02x5               g241(.a(new_n334), .b(new_n336), .c(new_n335), .d(new_n112), .o1(\s[8] ));
  xorb03aa1n02x5               g242(.a(new_n124), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


