// Benchmark "adder" written by ABC on Thu Jul 18 04:29:58 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n152, new_n153, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n178, new_n179, new_n180, new_n181,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n299, new_n302, new_n304, new_n305, new_n307;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  xnrc02aa1n03x5               g001(.a(\b[9] ), .b(\a[10] ), .out0(new_n97));
  orn002aa1n03x5               g002(.a(\a[9] ), .b(\b[8] ), .o(new_n98));
  and002aa1n02x5               g003(.a(\b[3] ), .b(\a[4] ), .o(new_n99));
  inv040aa1d32x5               g004(.a(\a[3] ), .o1(new_n100));
  inv030aa1d32x5               g005(.a(\b[2] ), .o1(new_n101));
  nand42aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  nanp02aa1n02x5               g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand02aa1n03x5               g008(.a(new_n102), .b(new_n103), .o1(new_n104));
  nor002aa1n03x5               g009(.a(\b[1] ), .b(\a[2] ), .o1(new_n105));
  nand02aa1d06x5               g010(.a(\b[0] ), .b(\a[1] ), .o1(new_n106));
  nand02aa1d06x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  aoi012aa1d18x5               g012(.a(new_n105), .b(new_n106), .c(new_n107), .o1(new_n108));
  inv000aa1d42x5               g013(.a(\a[4] ), .o1(new_n109));
  aboi22aa1n09x5               g014(.a(\b[3] ), .b(new_n109), .c(new_n100), .d(new_n101), .out0(new_n110));
  oaoi13aa1n12x5               g015(.a(new_n99), .b(new_n110), .c(new_n108), .d(new_n104), .o1(new_n111));
  norp02aa1n06x5               g016(.a(\b[7] ), .b(\a[8] ), .o1(new_n112));
  nand22aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nor022aa1n08x5               g018(.a(\b[6] ), .b(\a[7] ), .o1(new_n114));
  nand42aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nona23aa1n09x5               g020(.a(new_n115), .b(new_n113), .c(new_n112), .d(new_n114), .out0(new_n116));
  xorc02aa1n02x5               g021(.a(\a[6] ), .b(\b[5] ), .out0(new_n117));
  xorc02aa1n02x5               g022(.a(\a[5] ), .b(\b[4] ), .out0(new_n118));
  nano22aa1n03x7               g023(.a(new_n116), .b(new_n117), .c(new_n118), .out0(new_n119));
  inv000aa1d42x5               g024(.a(\b[5] ), .o1(new_n120));
  oai022aa1n02x5               g025(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n121));
  oaib12aa1n02x5               g026(.a(new_n121), .b(new_n120), .c(\a[6] ), .out0(new_n122));
  aoi012aa1n02x5               g027(.a(new_n112), .b(new_n114), .c(new_n113), .o1(new_n123));
  tech160nm_fioai012aa1n04x5   g028(.a(new_n123), .b(new_n116), .c(new_n122), .o1(new_n124));
  xorc02aa1n02x5               g029(.a(\a[9] ), .b(\b[8] ), .out0(new_n125));
  aoai13aa1n02x5               g030(.a(new_n125), .b(new_n124), .c(new_n119), .d(new_n111), .o1(new_n126));
  xobna2aa1n03x5               g031(.a(new_n97), .b(new_n126), .c(new_n98), .out0(\s[10] ));
  tech160nm_fioai012aa1n04x5   g032(.a(new_n110), .b(new_n108), .c(new_n104), .o1(new_n128));
  oaib12aa1n06x5               g033(.a(new_n128), .b(new_n109), .c(\b[3] ), .out0(new_n129));
  nanb03aa1n02x5               g034(.a(new_n116), .b(new_n118), .c(new_n117), .out0(new_n130));
  oabi12aa1n12x5               g035(.a(new_n124), .b(new_n129), .c(new_n130), .out0(new_n131));
  oaoi03aa1n12x5               g036(.a(\a[10] ), .b(\b[9] ), .c(new_n98), .o1(new_n132));
  nanp02aa1n02x5               g037(.a(\b[8] ), .b(\a[9] ), .o1(new_n133));
  nano22aa1n03x7               g038(.a(new_n97), .b(new_n98), .c(new_n133), .out0(new_n134));
  aoi012aa1n02x5               g039(.a(new_n132), .b(new_n131), .c(new_n134), .o1(new_n135));
  xnrb03aa1n02x5               g040(.a(new_n135), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  oaoi03aa1n02x5               g041(.a(\a[11] ), .b(\b[10] ), .c(new_n135), .o1(new_n137));
  xorb03aa1n02x5               g042(.a(new_n137), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  nor042aa1d18x5               g043(.a(\b[12] ), .b(\a[13] ), .o1(new_n139));
  nand42aa1d28x5               g044(.a(\b[12] ), .b(\a[13] ), .o1(new_n140));
  nanb02aa1n02x5               g045(.a(new_n139), .b(new_n140), .out0(new_n141));
  nor042aa1n02x5               g046(.a(\b[10] ), .b(\a[11] ), .o1(new_n142));
  nand42aa1n03x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  nor042aa1n02x5               g048(.a(\b[11] ), .b(\a[12] ), .o1(new_n144));
  nand42aa1n03x5               g049(.a(\b[11] ), .b(\a[12] ), .o1(new_n145));
  nano23aa1n03x7               g050(.a(new_n142), .b(new_n144), .c(new_n145), .d(new_n143), .out0(new_n146));
  nano22aa1n02x4               g051(.a(new_n97), .b(new_n146), .c(new_n125), .out0(new_n147));
  aoai13aa1n02x5               g052(.a(new_n147), .b(new_n124), .c(new_n119), .d(new_n111), .o1(new_n148));
  ao0012aa1n03x5               g053(.a(new_n144), .b(new_n142), .c(new_n145), .o(new_n149));
  aoi012aa1n06x5               g054(.a(new_n149), .b(new_n146), .c(new_n132), .o1(new_n150));
  xobna2aa1n03x5               g055(.a(new_n141), .b(new_n148), .c(new_n150), .out0(\s[13] ));
  inv000aa1d42x5               g056(.a(new_n139), .o1(new_n152));
  aoai13aa1n02x5               g057(.a(new_n152), .b(new_n141), .c(new_n148), .d(new_n150), .o1(new_n153));
  xorb03aa1n02x5               g058(.a(new_n153), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  nor042aa1n06x5               g059(.a(\b[13] ), .b(\a[14] ), .o1(new_n155));
  nand42aa1n16x5               g060(.a(\b[13] ), .b(\a[14] ), .o1(new_n156));
  nano23aa1d15x5               g061(.a(new_n139), .b(new_n155), .c(new_n156), .d(new_n140), .out0(new_n157));
  inv000aa1d42x5               g062(.a(new_n157), .o1(new_n158));
  oai012aa1n02x5               g063(.a(new_n156), .b(new_n155), .c(new_n139), .o1(new_n159));
  aoai13aa1n03x5               g064(.a(new_n159), .b(new_n158), .c(new_n148), .d(new_n150), .o1(new_n160));
  xorb03aa1n02x5               g065(.a(new_n160), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g066(.a(\b[14] ), .b(\a[15] ), .o1(new_n162));
  xorc02aa1n12x5               g067(.a(\a[15] ), .b(\b[14] ), .out0(new_n163));
  xorc02aa1n12x5               g068(.a(\a[16] ), .b(\b[15] ), .out0(new_n164));
  aoi112aa1n02x5               g069(.a(new_n164), .b(new_n162), .c(new_n160), .d(new_n163), .o1(new_n165));
  aoai13aa1n02x5               g070(.a(new_n164), .b(new_n162), .c(new_n160), .d(new_n163), .o1(new_n166));
  norb02aa1n02x5               g071(.a(new_n166), .b(new_n165), .out0(\s[16] ));
  nand23aa1d12x5               g072(.a(new_n157), .b(new_n163), .c(new_n164), .o1(new_n168));
  nano22aa1n12x5               g073(.a(new_n168), .b(new_n134), .c(new_n146), .out0(new_n169));
  aoai13aa1n06x5               g074(.a(new_n169), .b(new_n124), .c(new_n111), .d(new_n119), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(new_n164), .b(new_n163), .o1(new_n171));
  orn002aa1n02x5               g076(.a(\a[15] ), .b(\b[14] ), .o(new_n172));
  oao003aa1n02x5               g077(.a(\a[16] ), .b(\b[15] ), .c(new_n172), .carry(new_n173));
  oai012aa1n02x5               g078(.a(new_n173), .b(new_n171), .c(new_n159), .o1(new_n174));
  oab012aa1n09x5               g079(.a(new_n174), .b(new_n150), .c(new_n168), .out0(new_n175));
  nand02aa1d08x5               g080(.a(new_n170), .b(new_n175), .o1(new_n176));
  xorb03aa1n02x5               g081(.a(new_n176), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  inv000aa1d42x5               g082(.a(\a[18] ), .o1(new_n178));
  inv000aa1d42x5               g083(.a(\a[17] ), .o1(new_n179));
  inv000aa1d42x5               g084(.a(\b[16] ), .o1(new_n180));
  oaoi03aa1n02x5               g085(.a(new_n179), .b(new_n180), .c(new_n176), .o1(new_n181));
  xorb03aa1n02x5               g086(.a(new_n181), .b(\b[17] ), .c(new_n178), .out0(\s[18] ));
  xroi22aa1d04x5               g087(.a(new_n179), .b(\b[16] ), .c(new_n178), .d(\b[17] ), .out0(new_n183));
  nanp02aa1n02x5               g088(.a(new_n180), .b(new_n179), .o1(new_n184));
  oaoi03aa1n02x5               g089(.a(\a[18] ), .b(\b[17] ), .c(new_n184), .o1(new_n185));
  nor042aa1n04x5               g090(.a(\b[18] ), .b(\a[19] ), .o1(new_n186));
  nand02aa1n03x5               g091(.a(\b[18] ), .b(\a[19] ), .o1(new_n187));
  norb02aa1n02x5               g092(.a(new_n187), .b(new_n186), .out0(new_n188));
  aoai13aa1n06x5               g093(.a(new_n188), .b(new_n185), .c(new_n176), .d(new_n183), .o1(new_n189));
  aoi112aa1n02x5               g094(.a(new_n188), .b(new_n185), .c(new_n176), .d(new_n183), .o1(new_n190));
  norb02aa1n02x5               g095(.a(new_n189), .b(new_n190), .out0(\s[19] ));
  xnrc02aa1n02x5               g096(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor002aa1n04x5               g097(.a(\b[19] ), .b(\a[20] ), .o1(new_n193));
  nand02aa1d04x5               g098(.a(\b[19] ), .b(\a[20] ), .o1(new_n194));
  norb02aa1n02x5               g099(.a(new_n194), .b(new_n193), .out0(new_n195));
  nona22aa1n02x5               g100(.a(new_n189), .b(new_n195), .c(new_n186), .out0(new_n196));
  inv000aa1d42x5               g101(.a(new_n195), .o1(new_n197));
  oaoi13aa1n06x5               g102(.a(new_n197), .b(new_n189), .c(\a[19] ), .d(\b[18] ), .o1(new_n198));
  norb02aa1n03x4               g103(.a(new_n196), .b(new_n198), .out0(\s[20] ));
  nano23aa1n06x5               g104(.a(new_n186), .b(new_n193), .c(new_n194), .d(new_n187), .out0(new_n200));
  nanp02aa1n02x5               g105(.a(new_n183), .b(new_n200), .o1(new_n201));
  oai022aa1n02x5               g106(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n202));
  oaib12aa1n09x5               g107(.a(new_n202), .b(new_n178), .c(\b[17] ), .out0(new_n203));
  nona23aa1n09x5               g108(.a(new_n194), .b(new_n187), .c(new_n186), .d(new_n193), .out0(new_n204));
  aoi012aa1n12x5               g109(.a(new_n193), .b(new_n186), .c(new_n194), .o1(new_n205));
  oai012aa1n18x5               g110(.a(new_n205), .b(new_n204), .c(new_n203), .o1(new_n206));
  inv000aa1d42x5               g111(.a(new_n206), .o1(new_n207));
  aoai13aa1n06x5               g112(.a(new_n207), .b(new_n201), .c(new_n170), .d(new_n175), .o1(new_n208));
  xorb03aa1n02x5               g113(.a(new_n208), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  nor002aa1n02x5               g114(.a(\b[20] ), .b(\a[21] ), .o1(new_n210));
  xorc02aa1n02x5               g115(.a(\a[21] ), .b(\b[20] ), .out0(new_n211));
  xorc02aa1n02x5               g116(.a(\a[22] ), .b(\b[21] ), .out0(new_n212));
  aoi112aa1n02x5               g117(.a(new_n210), .b(new_n212), .c(new_n208), .d(new_n211), .o1(new_n213));
  aoai13aa1n03x5               g118(.a(new_n212), .b(new_n210), .c(new_n208), .d(new_n211), .o1(new_n214));
  norb02aa1n02x5               g119(.a(new_n214), .b(new_n213), .out0(\s[22] ));
  inv000aa1d42x5               g120(.a(\a[21] ), .o1(new_n216));
  inv000aa1d42x5               g121(.a(\a[22] ), .o1(new_n217));
  xroi22aa1d04x5               g122(.a(new_n216), .b(\b[20] ), .c(new_n217), .d(\b[21] ), .out0(new_n218));
  inv000aa1d42x5               g123(.a(\b[21] ), .o1(new_n219));
  oao003aa1n06x5               g124(.a(new_n217), .b(new_n219), .c(new_n210), .carry(new_n220));
  tech160nm_fiaoi012aa1n02p5x5 g125(.a(new_n220), .b(new_n206), .c(new_n218), .o1(new_n221));
  nand03aa1n02x5               g126(.a(new_n218), .b(new_n183), .c(new_n200), .o1(new_n222));
  aoai13aa1n04x5               g127(.a(new_n221), .b(new_n222), .c(new_n170), .d(new_n175), .o1(new_n223));
  xorb03aa1n02x5               g128(.a(new_n223), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g129(.a(\b[22] ), .b(\a[23] ), .o1(new_n225));
  xorc02aa1n03x5               g130(.a(\a[23] ), .b(\b[22] ), .out0(new_n226));
  xorc02aa1n02x5               g131(.a(\a[24] ), .b(\b[23] ), .out0(new_n227));
  aoi112aa1n03x5               g132(.a(new_n225), .b(new_n227), .c(new_n223), .d(new_n226), .o1(new_n228));
  aoai13aa1n03x5               g133(.a(new_n227), .b(new_n225), .c(new_n223), .d(new_n226), .o1(new_n229));
  norb02aa1n03x4               g134(.a(new_n229), .b(new_n228), .out0(\s[24] ));
  and002aa1n06x5               g135(.a(new_n227), .b(new_n226), .o(new_n231));
  inv040aa1n02x5               g136(.a(new_n231), .o1(new_n232));
  nano32aa1n02x4               g137(.a(new_n232), .b(new_n218), .c(new_n183), .d(new_n200), .out0(new_n233));
  inv020aa1n03x5               g138(.a(new_n205), .o1(new_n234));
  aoai13aa1n03x5               g139(.a(new_n218), .b(new_n234), .c(new_n200), .d(new_n185), .o1(new_n235));
  inv000aa1n02x5               g140(.a(new_n220), .o1(new_n236));
  aoi112aa1n02x5               g141(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n237));
  oab012aa1n02x4               g142(.a(new_n237), .b(\a[24] ), .c(\b[23] ), .out0(new_n238));
  aoai13aa1n06x5               g143(.a(new_n238), .b(new_n232), .c(new_n235), .d(new_n236), .o1(new_n239));
  xorc02aa1n02x5               g144(.a(\a[25] ), .b(\b[24] ), .out0(new_n240));
  aoai13aa1n06x5               g145(.a(new_n240), .b(new_n239), .c(new_n176), .d(new_n233), .o1(new_n241));
  aoi112aa1n02x5               g146(.a(new_n240), .b(new_n239), .c(new_n176), .d(new_n233), .o1(new_n242));
  norb02aa1n02x5               g147(.a(new_n241), .b(new_n242), .out0(\s[25] ));
  nor042aa1n03x5               g148(.a(\b[24] ), .b(\a[25] ), .o1(new_n244));
  xorc02aa1n02x5               g149(.a(\a[26] ), .b(\b[25] ), .out0(new_n245));
  nona22aa1n02x5               g150(.a(new_n241), .b(new_n245), .c(new_n244), .out0(new_n246));
  inv000aa1d42x5               g151(.a(new_n244), .o1(new_n247));
  aobi12aa1n06x5               g152(.a(new_n245), .b(new_n241), .c(new_n247), .out0(new_n248));
  norb02aa1n03x4               g153(.a(new_n246), .b(new_n248), .out0(\s[26] ));
  oai122aa1n02x7               g154(.a(new_n173), .b(new_n150), .c(new_n168), .d(new_n171), .e(new_n159), .o1(new_n250));
  inv000aa1d42x5               g155(.a(\a[25] ), .o1(new_n251));
  inv020aa1n04x5               g156(.a(\a[26] ), .o1(new_n252));
  xroi22aa1d06x4               g157(.a(new_n251), .b(\b[24] ), .c(new_n252), .d(\b[25] ), .out0(new_n253));
  nano22aa1n03x7               g158(.a(new_n222), .b(new_n231), .c(new_n253), .out0(new_n254));
  aoai13aa1n06x5               g159(.a(new_n254), .b(new_n250), .c(new_n131), .d(new_n169), .o1(new_n255));
  oao003aa1n02x5               g160(.a(\a[26] ), .b(\b[25] ), .c(new_n247), .carry(new_n256));
  aobi12aa1n06x5               g161(.a(new_n256), .b(new_n239), .c(new_n253), .out0(new_n257));
  norp02aa1n02x5               g162(.a(\b[26] ), .b(\a[27] ), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(\b[26] ), .b(\a[27] ), .o1(new_n259));
  norb02aa1n02x5               g164(.a(new_n259), .b(new_n258), .out0(new_n260));
  xnbna2aa1n03x5               g165(.a(new_n260), .b(new_n257), .c(new_n255), .out0(\s[27] ));
  inv000aa1n06x5               g166(.a(new_n258), .o1(new_n262));
  xnrc02aa1n02x5               g167(.a(\b[27] ), .b(\a[28] ), .out0(new_n263));
  aobi12aa1n06x5               g168(.a(new_n254), .b(new_n170), .c(new_n175), .out0(new_n264));
  aoai13aa1n06x5               g169(.a(new_n231), .b(new_n220), .c(new_n206), .d(new_n218), .o1(new_n265));
  inv000aa1d42x5               g170(.a(new_n253), .o1(new_n266));
  aoai13aa1n06x5               g171(.a(new_n256), .b(new_n266), .c(new_n265), .d(new_n238), .o1(new_n267));
  oaih12aa1n02x5               g172(.a(new_n259), .b(new_n267), .c(new_n264), .o1(new_n268));
  aoi012aa1n03x5               g173(.a(new_n263), .b(new_n268), .c(new_n262), .o1(new_n269));
  aoi022aa1n03x5               g174(.a(new_n257), .b(new_n255), .c(\a[27] ), .d(\b[26] ), .o1(new_n270));
  nano22aa1n03x5               g175(.a(new_n270), .b(new_n262), .c(new_n263), .out0(new_n271));
  norp02aa1n03x5               g176(.a(new_n269), .b(new_n271), .o1(\s[28] ));
  nano22aa1n02x4               g177(.a(new_n263), .b(new_n262), .c(new_n259), .out0(new_n273));
  oaih12aa1n02x5               g178(.a(new_n273), .b(new_n267), .c(new_n264), .o1(new_n274));
  oao003aa1n02x5               g179(.a(\a[28] ), .b(\b[27] ), .c(new_n262), .carry(new_n275));
  xnrc02aa1n02x5               g180(.a(\b[28] ), .b(\a[29] ), .out0(new_n276));
  aoi012aa1n03x5               g181(.a(new_n276), .b(new_n274), .c(new_n275), .o1(new_n277));
  aobi12aa1n02x7               g182(.a(new_n273), .b(new_n257), .c(new_n255), .out0(new_n278));
  nano22aa1n02x4               g183(.a(new_n278), .b(new_n275), .c(new_n276), .out0(new_n279));
  norp02aa1n03x5               g184(.a(new_n277), .b(new_n279), .o1(\s[29] ));
  xorb03aa1n02x5               g185(.a(new_n106), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g186(.a(new_n260), .b(new_n276), .c(new_n263), .out0(new_n282));
  oaih12aa1n02x5               g187(.a(new_n282), .b(new_n267), .c(new_n264), .o1(new_n283));
  oao003aa1n02x5               g188(.a(\a[29] ), .b(\b[28] ), .c(new_n275), .carry(new_n284));
  xnrc02aa1n02x5               g189(.a(\b[29] ), .b(\a[30] ), .out0(new_n285));
  aoi012aa1n03x5               g190(.a(new_n285), .b(new_n283), .c(new_n284), .o1(new_n286));
  aobi12aa1n06x5               g191(.a(new_n282), .b(new_n257), .c(new_n255), .out0(new_n287));
  nano22aa1n03x5               g192(.a(new_n287), .b(new_n284), .c(new_n285), .out0(new_n288));
  norp02aa1n03x5               g193(.a(new_n286), .b(new_n288), .o1(\s[30] ));
  xnrc02aa1n02x5               g194(.a(\b[30] ), .b(\a[31] ), .out0(new_n290));
  norb03aa1n02x5               g195(.a(new_n273), .b(new_n285), .c(new_n276), .out0(new_n291));
  aobi12aa1n06x5               g196(.a(new_n291), .b(new_n257), .c(new_n255), .out0(new_n292));
  oao003aa1n02x5               g197(.a(\a[30] ), .b(\b[29] ), .c(new_n284), .carry(new_n293));
  nano22aa1n03x5               g198(.a(new_n292), .b(new_n290), .c(new_n293), .out0(new_n294));
  oaih12aa1n02x5               g199(.a(new_n291), .b(new_n267), .c(new_n264), .o1(new_n295));
  aoi012aa1n03x5               g200(.a(new_n290), .b(new_n295), .c(new_n293), .o1(new_n296));
  norp02aa1n03x5               g201(.a(new_n296), .b(new_n294), .o1(\s[31] ));
  xnbna2aa1n03x5               g202(.a(new_n108), .b(new_n102), .c(new_n103), .out0(\s[3] ));
  oaoi03aa1n02x5               g203(.a(\a[3] ), .b(\b[2] ), .c(new_n108), .o1(new_n299));
  xorb03aa1n02x5               g204(.a(new_n299), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xorb03aa1n02x5               g205(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  oaoi03aa1n02x5               g206(.a(\a[5] ), .b(\b[4] ), .c(new_n129), .o1(new_n302));
  xorb03aa1n02x5               g207(.a(new_n302), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g208(.a(\a[6] ), .o1(new_n304));
  oaoi03aa1n02x5               g209(.a(new_n304), .b(new_n120), .c(new_n302), .o1(new_n305));
  xnrb03aa1n02x5               g210(.a(new_n305), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g211(.a(\a[7] ), .b(\b[6] ), .c(new_n305), .o1(new_n307));
  xorb03aa1n02x5               g212(.a(new_n307), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g213(.a(new_n131), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


