// Benchmark "adder" written by ABC on Thu Jul 18 07:48:39 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n181, new_n182, new_n183, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n336, new_n339, new_n340,
    new_n342, new_n343, new_n345, new_n346, new_n347, new_n348;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  inv000aa1d42x5               g001(.a(\a[1] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(\b[0] ), .o1(new_n98));
  norp02aa1n02x5               g003(.a(\b[1] ), .b(\a[2] ), .o1(new_n99));
  nanp02aa1n02x5               g004(.a(\b[1] ), .b(\a[2] ), .o1(new_n100));
  oaoi13aa1n06x5               g005(.a(new_n99), .b(new_n100), .c(new_n97), .d(new_n98), .o1(new_n101));
  nand02aa1n03x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  nor022aa1n08x5               g007(.a(\b[3] ), .b(\a[4] ), .o1(new_n103));
  nor042aa1n04x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nand42aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nona23aa1n03x5               g010(.a(new_n102), .b(new_n105), .c(new_n104), .d(new_n103), .out0(new_n106));
  inv000aa1d42x5               g011(.a(\a[3] ), .o1(new_n107));
  inv000aa1d42x5               g012(.a(\b[2] ), .o1(new_n108));
  aoai13aa1n04x5               g013(.a(new_n102), .b(new_n103), .c(new_n108), .d(new_n107), .o1(new_n109));
  oaih12aa1n06x5               g014(.a(new_n109), .b(new_n106), .c(new_n101), .o1(new_n110));
  xnrc02aa1n12x5               g015(.a(\b[5] ), .b(\a[6] ), .out0(new_n111));
  xnrc02aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .out0(new_n112));
  norp02aa1n04x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nand02aa1d04x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  nand42aa1n03x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  norp02aa1n12x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n09x5               g021(.a(new_n115), .b(new_n114), .c(new_n116), .d(new_n113), .out0(new_n117));
  nor043aa1n03x5               g022(.a(new_n117), .b(new_n112), .c(new_n111), .o1(new_n118));
  inv000aa1d42x5               g023(.a(\a[6] ), .o1(new_n119));
  inv000aa1d42x5               g024(.a(\b[5] ), .o1(new_n120));
  norp02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  oaoi03aa1n02x5               g026(.a(new_n119), .b(new_n120), .c(new_n121), .o1(new_n122));
  tech160nm_fiao0012aa1n02p5x5 g027(.a(new_n113), .b(new_n116), .c(new_n114), .o(new_n123));
  oabi12aa1n06x5               g028(.a(new_n123), .b(new_n117), .c(new_n122), .out0(new_n124));
  nor042aa1n06x5               g029(.a(\b[8] ), .b(\a[9] ), .o1(new_n125));
  nanp02aa1n04x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n125), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n128));
  oai012aa1n02x5               g033(.a(new_n128), .b(\b[8] ), .c(\a[9] ), .o1(new_n129));
  xorb03aa1n02x5               g034(.a(new_n129), .b(\b[9] ), .c(\a[10] ), .out0(\s[10] ));
  nor002aa1n20x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  inv000aa1d42x5               g036(.a(new_n131), .o1(new_n132));
  nand42aa1n16x5               g037(.a(\b[9] ), .b(\a[10] ), .o1(new_n133));
  and002aa1n02x5               g038(.a(\b[0] ), .b(\a[1] ), .o(new_n134));
  oaoi03aa1n02x5               g039(.a(\a[2] ), .b(\b[1] ), .c(new_n134), .o1(new_n135));
  norb02aa1n02x5               g040(.a(new_n102), .b(new_n103), .out0(new_n136));
  norb02aa1n02x5               g041(.a(new_n105), .b(new_n104), .out0(new_n137));
  nanp03aa1n03x5               g042(.a(new_n135), .b(new_n136), .c(new_n137), .o1(new_n138));
  nano23aa1n03x5               g043(.a(new_n116), .b(new_n113), .c(new_n114), .d(new_n115), .out0(new_n139));
  nona22aa1n02x4               g044(.a(new_n139), .b(new_n112), .c(new_n111), .out0(new_n140));
  oao003aa1n02x5               g045(.a(new_n119), .b(new_n120), .c(new_n121), .carry(new_n141));
  aoi012aa1n02x5               g046(.a(new_n123), .b(new_n139), .c(new_n141), .o1(new_n142));
  aoai13aa1n06x5               g047(.a(new_n142), .b(new_n140), .c(new_n138), .d(new_n109), .o1(new_n143));
  aoai13aa1n02x5               g048(.a(new_n133), .b(new_n125), .c(new_n143), .d(new_n127), .o1(new_n144));
  nand42aa1n08x5               g049(.a(\b[10] ), .b(\a[11] ), .o1(new_n145));
  nor042aa1n06x5               g050(.a(\b[10] ), .b(\a[11] ), .o1(new_n146));
  nanb02aa1n02x5               g051(.a(new_n146), .b(new_n145), .out0(new_n147));
  inv000aa1d42x5               g052(.a(new_n147), .o1(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n144), .c(new_n132), .out0(\s[11] ));
  aoai13aa1n02x5               g054(.a(new_n148), .b(new_n131), .c(new_n129), .d(new_n133), .o1(new_n150));
  nor042aa1n06x5               g055(.a(\b[11] ), .b(\a[12] ), .o1(new_n151));
  nanp02aa1n12x5               g056(.a(\b[11] ), .b(\a[12] ), .o1(new_n152));
  norb02aa1n02x5               g057(.a(new_n152), .b(new_n151), .out0(new_n153));
  inv000aa1d42x5               g058(.a(\a[11] ), .o1(new_n154));
  inv000aa1d42x5               g059(.a(\b[10] ), .o1(new_n155));
  aboi22aa1n06x5               g060(.a(new_n151), .b(new_n152), .c(new_n154), .d(new_n155), .out0(new_n156));
  inv000aa1n03x5               g061(.a(new_n146), .o1(new_n157));
  aoai13aa1n02x5               g062(.a(new_n157), .b(new_n147), .c(new_n144), .d(new_n132), .o1(new_n158));
  aoi022aa1n02x5               g063(.a(new_n158), .b(new_n153), .c(new_n150), .d(new_n156), .o1(\s[12] ));
  oaib12aa1n09x5               g064(.a(new_n157), .b(new_n151), .c(new_n152), .out0(new_n160));
  norb03aa1n09x5               g065(.a(new_n126), .b(new_n131), .c(new_n125), .out0(new_n161));
  nano22aa1n09x5               g066(.a(new_n146), .b(new_n133), .c(new_n145), .out0(new_n162));
  nand23aa1d12x5               g067(.a(new_n160), .b(new_n162), .c(new_n161), .o1(new_n163));
  inv000aa1d42x5               g068(.a(new_n163), .o1(new_n164));
  aoai13aa1n06x5               g069(.a(new_n164), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n165));
  nanb03aa1n12x5               g070(.a(new_n146), .b(new_n133), .c(new_n145), .out0(new_n166));
  norb03aa1n06x5               g071(.a(new_n133), .b(new_n131), .c(new_n125), .out0(new_n167));
  aoi012aa1n02x7               g072(.a(new_n151), .b(new_n146), .c(new_n152), .o1(new_n168));
  oai013aa1d12x5               g073(.a(new_n168), .b(new_n156), .c(new_n167), .d(new_n166), .o1(new_n169));
  inv000aa1d42x5               g074(.a(new_n169), .o1(new_n170));
  nand42aa1n03x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  nor042aa1n03x5               g076(.a(\b[12] ), .b(\a[13] ), .o1(new_n172));
  norb02aa1n03x5               g077(.a(new_n171), .b(new_n172), .out0(new_n173));
  xnbna2aa1n03x5               g078(.a(new_n173), .b(new_n165), .c(new_n170), .out0(\s[13] ));
  orn002aa1n02x5               g079(.a(\a[13] ), .b(\b[12] ), .o(new_n175));
  aoai13aa1n02x5               g080(.a(new_n173), .b(new_n169), .c(new_n143), .d(new_n164), .o1(new_n176));
  nor002aa1n04x5               g081(.a(\b[13] ), .b(\a[14] ), .o1(new_n177));
  nanp02aa1n09x5               g082(.a(\b[13] ), .b(\a[14] ), .o1(new_n178));
  norb02aa1n03x5               g083(.a(new_n178), .b(new_n177), .out0(new_n179));
  xnbna2aa1n03x5               g084(.a(new_n179), .b(new_n176), .c(new_n175), .out0(\s[14] ));
  nona23aa1n02x4               g085(.a(new_n171), .b(new_n178), .c(new_n177), .d(new_n172), .out0(new_n181));
  tech160nm_fiaoi012aa1n05x5   g086(.a(new_n177), .b(new_n172), .c(new_n178), .o1(new_n182));
  aoai13aa1n06x5               g087(.a(new_n182), .b(new_n181), .c(new_n165), .d(new_n170), .o1(new_n183));
  xorb03aa1n02x5               g088(.a(new_n183), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor042aa1n03x5               g089(.a(\b[14] ), .b(\a[15] ), .o1(new_n185));
  nand22aa1n03x5               g090(.a(\b[14] ), .b(\a[15] ), .o1(new_n186));
  norb02aa1n02x7               g091(.a(new_n186), .b(new_n185), .out0(new_n187));
  nor042aa1n02x5               g092(.a(\b[15] ), .b(\a[16] ), .o1(new_n188));
  nand02aa1n03x5               g093(.a(\b[15] ), .b(\a[16] ), .o1(new_n189));
  nanb02aa1n02x5               g094(.a(new_n188), .b(new_n189), .out0(new_n190));
  aoai13aa1n02x5               g095(.a(new_n190), .b(new_n185), .c(new_n183), .d(new_n187), .o1(new_n191));
  nand22aa1n02x5               g096(.a(new_n183), .b(new_n187), .o1(new_n192));
  nona22aa1n02x4               g097(.a(new_n192), .b(new_n190), .c(new_n185), .out0(new_n193));
  nanp02aa1n03x5               g098(.a(new_n193), .b(new_n191), .o1(\s[16] ));
  nano23aa1n06x5               g099(.a(new_n188), .b(new_n185), .c(new_n189), .d(new_n186), .out0(new_n195));
  nano32aa1d12x5               g100(.a(new_n163), .b(new_n195), .c(new_n173), .d(new_n179), .out0(new_n196));
  aoai13aa1n12x5               g101(.a(new_n196), .b(new_n124), .c(new_n110), .d(new_n118), .o1(new_n197));
  nano32aa1n03x7               g102(.a(new_n190), .b(new_n187), .c(new_n179), .d(new_n173), .out0(new_n198));
  inv000aa1n02x5               g103(.a(new_n182), .o1(new_n199));
  oa0012aa1n02x5               g104(.a(new_n189), .b(new_n188), .c(new_n185), .o(new_n200));
  aoi012aa1n02x7               g105(.a(new_n200), .b(new_n195), .c(new_n199), .o1(new_n201));
  aobi12aa1d24x5               g106(.a(new_n201), .b(new_n169), .c(new_n198), .out0(new_n202));
  xorc02aa1n02x5               g107(.a(\a[17] ), .b(\b[16] ), .out0(new_n203));
  xnbna2aa1n03x5               g108(.a(new_n203), .b(new_n197), .c(new_n202), .out0(\s[17] ));
  inv040aa1d32x5               g109(.a(\a[18] ), .o1(new_n205));
  inv040aa1d30x5               g110(.a(\a[17] ), .o1(new_n206));
  inv000aa1d42x5               g111(.a(\b[16] ), .o1(new_n207));
  nanp02aa1n06x5               g112(.a(new_n197), .b(new_n202), .o1(new_n208));
  oaoi03aa1n03x5               g113(.a(new_n206), .b(new_n207), .c(new_n208), .o1(new_n209));
  xorb03aa1n02x5               g114(.a(new_n209), .b(\b[17] ), .c(new_n205), .out0(\s[18] ));
  xroi22aa1d06x4               g115(.a(new_n206), .b(\b[16] ), .c(new_n205), .d(\b[17] ), .out0(new_n211));
  inv000aa1d42x5               g116(.a(new_n211), .o1(new_n212));
  nor002aa1n02x5               g117(.a(\b[17] ), .b(\a[18] ), .o1(new_n213));
  aoi112aa1n09x5               g118(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n214));
  norp02aa1n02x5               g119(.a(new_n214), .b(new_n213), .o1(new_n215));
  aoai13aa1n04x5               g120(.a(new_n215), .b(new_n212), .c(new_n197), .d(new_n202), .o1(new_n216));
  xorb03aa1n02x5               g121(.a(new_n216), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g122(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  tech160nm_finand02aa1n03p5x5 g123(.a(\b[18] ), .b(\a[19] ), .o1(new_n219));
  nor042aa1n04x5               g124(.a(\b[18] ), .b(\a[19] ), .o1(new_n220));
  nor002aa1n06x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nand42aa1n06x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  norb02aa1n12x5               g127(.a(new_n222), .b(new_n221), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoai13aa1n03x5               g129(.a(new_n224), .b(new_n220), .c(new_n216), .d(new_n219), .o1(new_n225));
  norb02aa1n02x7               g130(.a(new_n219), .b(new_n220), .out0(new_n226));
  nand02aa1n02x5               g131(.a(new_n216), .b(new_n226), .o1(new_n227));
  nona22aa1n02x4               g132(.a(new_n227), .b(new_n224), .c(new_n220), .out0(new_n228));
  nanp02aa1n03x5               g133(.a(new_n228), .b(new_n225), .o1(\s[20] ));
  nano23aa1n02x4               g134(.a(new_n221), .b(new_n220), .c(new_n222), .d(new_n219), .out0(new_n230));
  nand02aa1n02x5               g135(.a(new_n211), .b(new_n230), .o1(new_n231));
  oai112aa1n06x5               g136(.a(new_n226), .b(new_n223), .c(new_n214), .d(new_n213), .o1(new_n232));
  oaih12aa1n02x5               g137(.a(new_n222), .b(new_n221), .c(new_n220), .o1(new_n233));
  nand22aa1n09x5               g138(.a(new_n232), .b(new_n233), .o1(new_n234));
  inv000aa1d42x5               g139(.a(new_n234), .o1(new_n235));
  aoai13aa1n04x5               g140(.a(new_n235), .b(new_n231), .c(new_n197), .d(new_n202), .o1(new_n236));
  xorb03aa1n02x5               g141(.a(new_n236), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n04x5               g142(.a(\b[20] ), .b(\a[21] ), .o1(new_n238));
  nand42aa1n03x5               g143(.a(\b[20] ), .b(\a[21] ), .o1(new_n239));
  norb02aa1n02x5               g144(.a(new_n239), .b(new_n238), .out0(new_n240));
  nor022aa1n08x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  nand42aa1n03x5               g146(.a(\b[21] ), .b(\a[22] ), .o1(new_n242));
  norb02aa1n06x5               g147(.a(new_n242), .b(new_n241), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n243), .o1(new_n244));
  aoai13aa1n03x5               g149(.a(new_n244), .b(new_n238), .c(new_n236), .d(new_n240), .o1(new_n245));
  nand02aa1n02x5               g150(.a(new_n236), .b(new_n240), .o1(new_n246));
  nona22aa1n02x4               g151(.a(new_n246), .b(new_n244), .c(new_n238), .out0(new_n247));
  nanp02aa1n03x5               g152(.a(new_n247), .b(new_n245), .o1(\s[22] ));
  nano23aa1n03x5               g153(.a(new_n241), .b(new_n238), .c(new_n242), .d(new_n239), .out0(new_n249));
  nand23aa1n03x5               g154(.a(new_n211), .b(new_n230), .c(new_n249), .o1(new_n250));
  tech160nm_fiao0012aa1n02p5x5 g155(.a(new_n241), .b(new_n238), .c(new_n242), .o(new_n251));
  aoi012aa1n02x5               g156(.a(new_n251), .b(new_n234), .c(new_n249), .o1(new_n252));
  aoai13aa1n04x5               g157(.a(new_n252), .b(new_n250), .c(new_n197), .d(new_n202), .o1(new_n253));
  xorb03aa1n02x5               g158(.a(new_n253), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n02x5               g159(.a(\b[22] ), .b(\a[23] ), .o1(new_n255));
  nand42aa1n03x5               g160(.a(\b[22] ), .b(\a[23] ), .o1(new_n256));
  norb02aa1n02x5               g161(.a(new_n256), .b(new_n255), .out0(new_n257));
  nor002aa1n03x5               g162(.a(\b[23] ), .b(\a[24] ), .o1(new_n258));
  nanp02aa1n02x5               g163(.a(\b[23] ), .b(\a[24] ), .o1(new_n259));
  nanb02aa1n02x5               g164(.a(new_n258), .b(new_n259), .out0(new_n260));
  aoai13aa1n03x5               g165(.a(new_n260), .b(new_n255), .c(new_n253), .d(new_n257), .o1(new_n261));
  nand02aa1n02x5               g166(.a(new_n253), .b(new_n257), .o1(new_n262));
  nona22aa1n02x4               g167(.a(new_n262), .b(new_n260), .c(new_n255), .out0(new_n263));
  nanp02aa1n03x5               g168(.a(new_n263), .b(new_n261), .o1(\s[24] ));
  nano23aa1n03x5               g169(.a(new_n255), .b(new_n258), .c(new_n259), .d(new_n256), .out0(new_n265));
  nanb03aa1n03x5               g170(.a(new_n231), .b(new_n265), .c(new_n249), .out0(new_n266));
  aoi012aa1n02x5               g171(.a(new_n266), .b(new_n197), .c(new_n202), .o1(new_n267));
  nano32aa1n02x4               g172(.a(new_n260), .b(new_n257), .c(new_n243), .d(new_n240), .out0(new_n268));
  aoi112aa1n02x5               g173(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n269));
  nanp02aa1n03x5               g174(.a(new_n265), .b(new_n251), .o1(new_n270));
  nona22aa1n03x5               g175(.a(new_n270), .b(new_n269), .c(new_n258), .out0(new_n271));
  tech160nm_fiaoi012aa1n04x5   g176(.a(new_n271), .b(new_n234), .c(new_n268), .o1(new_n272));
  aoai13aa1n04x5               g177(.a(new_n272), .b(new_n266), .c(new_n197), .d(new_n202), .o1(new_n273));
  xorc02aa1n12x5               g178(.a(\a[25] ), .b(\b[24] ), .out0(new_n274));
  nand02aa1n02x5               g179(.a(new_n265), .b(new_n249), .o1(new_n275));
  aoi012aa1n03x5               g180(.a(new_n275), .b(new_n232), .c(new_n233), .o1(new_n276));
  norp03aa1n02x5               g181(.a(new_n276), .b(new_n271), .c(new_n274), .o1(new_n277));
  aboi22aa1n03x5               g182(.a(new_n267), .b(new_n277), .c(new_n273), .d(new_n274), .out0(\s[25] ));
  norp02aa1n02x5               g183(.a(\b[24] ), .b(\a[25] ), .o1(new_n279));
  tech160nm_fixnrc02aa1n05x5   g184(.a(\b[25] ), .b(\a[26] ), .out0(new_n280));
  aoai13aa1n03x5               g185(.a(new_n280), .b(new_n279), .c(new_n273), .d(new_n274), .o1(new_n281));
  nand02aa1n02x5               g186(.a(new_n273), .b(new_n274), .o1(new_n282));
  nona22aa1n02x4               g187(.a(new_n282), .b(new_n280), .c(new_n279), .out0(new_n283));
  nanp02aa1n03x5               g188(.a(new_n283), .b(new_n281), .o1(\s[26] ));
  nanb03aa1n02x5               g189(.a(new_n167), .b(new_n160), .c(new_n162), .out0(new_n285));
  nanp03aa1n02x5               g190(.a(new_n195), .b(new_n173), .c(new_n179), .o1(new_n286));
  aoai13aa1n02x5               g191(.a(new_n201), .b(new_n286), .c(new_n285), .d(new_n168), .o1(new_n287));
  norb02aa1n06x5               g192(.a(new_n274), .b(new_n280), .out0(new_n288));
  nano22aa1n03x7               g193(.a(new_n250), .b(new_n265), .c(new_n288), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n287), .c(new_n143), .d(new_n196), .o1(new_n290));
  orn002aa1n02x5               g195(.a(\a[25] ), .b(\b[24] ), .o(new_n291));
  oaoi03aa1n02x5               g196(.a(\a[26] ), .b(\b[25] ), .c(new_n291), .o1(new_n292));
  oaoi13aa1n06x5               g197(.a(new_n292), .b(new_n288), .c(new_n276), .d(new_n271), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  xnbna2aa1n03x5               g199(.a(new_n294), .b(new_n290), .c(new_n293), .out0(\s[27] ));
  inv020aa1n03x5               g200(.a(new_n289), .o1(new_n296));
  aoai13aa1n04x5               g201(.a(new_n293), .b(new_n296), .c(new_n197), .d(new_n202), .o1(new_n297));
  nor042aa1n09x5               g202(.a(\b[26] ), .b(\a[27] ), .o1(new_n298));
  nor042aa1n02x5               g203(.a(\b[27] ), .b(\a[28] ), .o1(new_n299));
  nand02aa1d08x5               g204(.a(\b[27] ), .b(\a[28] ), .o1(new_n300));
  nanb02aa1n06x5               g205(.a(new_n299), .b(new_n300), .out0(new_n301));
  aoai13aa1n03x5               g206(.a(new_n301), .b(new_n298), .c(new_n297), .d(new_n294), .o1(new_n302));
  inv000aa1d42x5               g207(.a(new_n288), .o1(new_n303));
  oabi12aa1n02x7               g208(.a(new_n292), .b(new_n272), .c(new_n303), .out0(new_n304));
  aoai13aa1n02x7               g209(.a(new_n294), .b(new_n304), .c(new_n208), .d(new_n289), .o1(new_n305));
  nona22aa1n02x5               g210(.a(new_n305), .b(new_n301), .c(new_n298), .out0(new_n306));
  nanp02aa1n03x5               g211(.a(new_n302), .b(new_n306), .o1(\s[28] ));
  norb02aa1d27x5               g212(.a(new_n294), .b(new_n301), .out0(new_n308));
  aoai13aa1n03x5               g213(.a(new_n308), .b(new_n304), .c(new_n208), .d(new_n289), .o1(new_n309));
  inv000aa1d42x5               g214(.a(new_n308), .o1(new_n310));
  aoi012aa1n06x5               g215(.a(new_n299), .b(new_n298), .c(new_n300), .o1(new_n311));
  aoai13aa1n02x7               g216(.a(new_n311), .b(new_n310), .c(new_n290), .d(new_n293), .o1(new_n312));
  xorc02aa1n02x5               g217(.a(\a[29] ), .b(\b[28] ), .out0(new_n313));
  norb02aa1n02x5               g218(.a(new_n311), .b(new_n313), .out0(new_n314));
  aoi022aa1n03x5               g219(.a(new_n312), .b(new_n313), .c(new_n309), .d(new_n314), .o1(\s[29] ));
  xnrb03aa1n02x5               g220(.a(new_n134), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nanb03aa1n02x5               g221(.a(new_n301), .b(new_n313), .c(new_n294), .out0(new_n317));
  nanb02aa1n03x5               g222(.a(new_n317), .b(new_n297), .out0(new_n318));
  tech160nm_fioaoi03aa1n02p5x5 g223(.a(\a[29] ), .b(\b[28] ), .c(new_n311), .o1(new_n319));
  inv000aa1d42x5               g224(.a(new_n319), .o1(new_n320));
  aoai13aa1n02x7               g225(.a(new_n320), .b(new_n317), .c(new_n290), .d(new_n293), .o1(new_n321));
  xorc02aa1n02x5               g226(.a(\a[30] ), .b(\b[29] ), .out0(new_n322));
  norp02aa1n02x5               g227(.a(new_n319), .b(new_n322), .o1(new_n323));
  aoi022aa1n03x5               g228(.a(new_n321), .b(new_n322), .c(new_n318), .d(new_n323), .o1(\s[30] ));
  nanp03aa1n02x5               g229(.a(new_n308), .b(new_n313), .c(new_n322), .o1(new_n325));
  nanb02aa1n03x5               g230(.a(new_n325), .b(new_n297), .out0(new_n326));
  xorc02aa1n02x5               g231(.a(\a[31] ), .b(\b[30] ), .out0(new_n327));
  inv000aa1d42x5               g232(.a(\a[30] ), .o1(new_n328));
  inv000aa1d42x5               g233(.a(\b[29] ), .o1(new_n329));
  oabi12aa1n02x5               g234(.a(new_n327), .b(\a[30] ), .c(\b[29] ), .out0(new_n330));
  oaoi13aa1n02x5               g235(.a(new_n330), .b(new_n319), .c(new_n328), .d(new_n329), .o1(new_n331));
  oaoi03aa1n02x5               g236(.a(new_n328), .b(new_n329), .c(new_n319), .o1(new_n332));
  aoai13aa1n02x7               g237(.a(new_n332), .b(new_n325), .c(new_n290), .d(new_n293), .o1(new_n333));
  aoi022aa1n03x5               g238(.a(new_n333), .b(new_n327), .c(new_n326), .d(new_n331), .o1(\s[31] ));
  xorb03aa1n02x5               g239(.a(new_n101), .b(\b[2] ), .c(new_n107), .out0(\s[3] ));
  aoi112aa1n02x5               g240(.a(new_n104), .b(new_n136), .c(new_n135), .d(new_n105), .o1(new_n336));
  aoib12aa1n02x5               g241(.a(new_n336), .b(new_n110), .c(new_n103), .out0(\s[4] ));
  xorb03aa1n02x5               g242(.a(new_n110), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  orn002aa1n02x5               g243(.a(\a[5] ), .b(\b[4] ), .o(new_n339));
  aoai13aa1n02x5               g244(.a(new_n339), .b(new_n112), .c(new_n138), .d(new_n109), .o1(new_n340));
  xorb03aa1n02x5               g245(.a(new_n340), .b(\b[5] ), .c(\a[6] ), .out0(\s[6] ));
  inv000aa1d42x5               g246(.a(new_n111), .o1(new_n342));
  aob012aa1n02x5               g247(.a(new_n122), .b(new_n340), .c(new_n342), .out0(new_n343));
  xorb03aa1n02x5               g248(.a(new_n343), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  nanb02aa1n02x5               g249(.a(new_n116), .b(new_n115), .out0(new_n345));
  inv000aa1d42x5               g250(.a(new_n345), .o1(new_n346));
  aoai13aa1n03x5               g251(.a(new_n346), .b(new_n141), .c(new_n340), .d(new_n342), .o1(new_n347));
  oai012aa1n02x5               g252(.a(new_n347), .b(\b[6] ), .c(\a[7] ), .o1(new_n348));
  xorb03aa1n02x5               g253(.a(new_n348), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xorb03aa1n02x5               g254(.a(new_n143), .b(\b[8] ), .c(\a[9] ), .out0(\s[9] ));
endmodule


