// Benchmark "adder" written by ABC on Thu Jul 11 11:45:12 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n149, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n165, new_n166, new_n167, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n346, new_n349, new_n351, new_n353;
  160nm_ficinv00aa1n08x5       g000(.clk(\a[0] ), .clkout(\s[0] ));
  norp02aa1n02x5               g001(.a(\b[9] ), .b(\a[10] ), .o1(new_n97));
  nanp02aa1n02x5               g002(.a(\b[9] ), .b(\a[10] ), .o1(new_n98));
  nanb02aa1n02x5               g003(.a(new_n97), .b(new_n98), .out0(new_n99));
  160nm_ficinv00aa1n08x5       g004(.clk(\a[9] ), .clkout(new_n100));
  160nm_ficinv00aa1n08x5       g005(.clk(\b[8] ), .clkout(new_n101));
  nanp02aa1n02x5               g006(.a(new_n101), .b(new_n100), .o1(new_n102));
  and002aa1n02x5               g007(.a(\b[3] ), .b(\a[4] ), .o(new_n103));
  norp02aa1n02x5               g008(.a(\b[2] ), .b(\a[3] ), .o1(new_n104));
  nanp02aa1n02x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb02aa1n02x5               g010(.a(new_n104), .b(new_n105), .out0(new_n106));
  norp02aa1n02x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nanp02aa1n02x5               g012(.a(\b[0] ), .b(\a[1] ), .o1(new_n108));
  nanp02aa1n02x5               g013(.a(\b[1] ), .b(\a[2] ), .o1(new_n109));
  aoi012aa1n02x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  oab012aa1n02x4               g015(.a(new_n104), .b(\a[4] ), .c(\b[3] ), .out0(new_n111));
  oaoi13aa1n02x5               g016(.a(new_n103), .b(new_n111), .c(new_n110), .d(new_n106), .o1(new_n112));
  norp02aa1n02x5               g017(.a(\b[7] ), .b(\a[8] ), .o1(new_n113));
  nanp02aa1n02x5               g018(.a(\b[7] ), .b(\a[8] ), .o1(new_n114));
  norp02aa1n02x5               g019(.a(\b[6] ), .b(\a[7] ), .o1(new_n115));
  nanp02aa1n02x5               g020(.a(\b[6] ), .b(\a[7] ), .o1(new_n116));
  nona23aa1n02x4               g021(.a(new_n116), .b(new_n114), .c(new_n113), .d(new_n115), .out0(new_n117));
  norp02aa1n02x5               g022(.a(\b[5] ), .b(\a[6] ), .o1(new_n118));
  nanp02aa1n02x5               g023(.a(\b[5] ), .b(\a[6] ), .o1(new_n119));
  norb02aa1n02x5               g024(.a(new_n119), .b(new_n118), .out0(new_n120));
  norp02aa1n02x5               g025(.a(\b[4] ), .b(\a[5] ), .o1(new_n121));
  nanp02aa1n02x5               g026(.a(\b[4] ), .b(\a[5] ), .o1(new_n122));
  norb02aa1n02x5               g027(.a(new_n122), .b(new_n121), .out0(new_n123));
  nano22aa1n02x4               g028(.a(new_n117), .b(new_n120), .c(new_n123), .out0(new_n124));
  oai012aa1n02x5               g029(.a(new_n119), .b(new_n121), .c(new_n118), .o1(new_n125));
  160nm_fiao0012aa1n02p5x5     g030(.a(new_n113), .b(new_n115), .c(new_n114), .o(new_n126));
  oabi12aa1n02x5               g031(.a(new_n126), .b(new_n117), .c(new_n125), .out0(new_n127));
  xorc02aa1n02x5               g032(.a(\a[9] ), .b(\b[8] ), .out0(new_n128));
  aoai13aa1n02x5               g033(.a(new_n128), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n129));
  xobna2aa1n03x5               g034(.a(new_n99), .b(new_n129), .c(new_n102), .out0(\s[10] ));
  160nm_ficinv00aa1n08x5       g035(.clk(new_n103), .clkout(new_n131));
  norb02aa1n02x5               g036(.a(new_n105), .b(new_n104), .out0(new_n132));
  160nm_ficinv00aa1n08x5       g037(.clk(new_n107), .clkout(new_n133));
  nanp02aa1n02x5               g038(.a(new_n109), .b(new_n108), .o1(new_n134));
  nanp02aa1n02x5               g039(.a(new_n134), .b(new_n133), .o1(new_n135));
  160nm_ficinv00aa1n08x5       g040(.clk(new_n111), .clkout(new_n136));
  aoai13aa1n02x5               g041(.a(new_n131), .b(new_n136), .c(new_n135), .d(new_n132), .o1(new_n137));
  nano23aa1n02x4               g042(.a(new_n113), .b(new_n115), .c(new_n116), .d(new_n114), .out0(new_n138));
  nano23aa1n02x4               g043(.a(new_n118), .b(new_n121), .c(new_n122), .d(new_n119), .out0(new_n139));
  nanp02aa1n02x5               g044(.a(new_n139), .b(new_n138), .o1(new_n140));
  aoib12aa1n02x5               g045(.a(new_n126), .b(new_n138), .c(new_n125), .out0(new_n141));
  oai012aa1n02x5               g046(.a(new_n141), .b(new_n137), .c(new_n140), .o1(new_n142));
  aoai13aa1n02x5               g047(.a(new_n98), .b(new_n97), .c(new_n100), .d(new_n101), .o1(new_n143));
  160nm_ficinv00aa1n08x5       g048(.clk(new_n143), .clkout(new_n144));
  nanp02aa1n02x5               g049(.a(\b[8] ), .b(\a[9] ), .o1(new_n145));
  nano22aa1n02x4               g050(.a(new_n99), .b(new_n102), .c(new_n145), .out0(new_n146));
  aoi012aa1n02x5               g051(.a(new_n144), .b(new_n142), .c(new_n146), .o1(new_n147));
  xnrb03aa1n02x5               g052(.a(new_n147), .b(\b[10] ), .c(\a[11] ), .out0(\s[11] ));
  oaoi03aa1n02x5               g053(.a(\a[11] ), .b(\b[10] ), .c(new_n147), .o1(new_n149));
  xorb03aa1n02x5               g054(.a(new_n149), .b(\b[11] ), .c(\a[12] ), .out0(\s[12] ));
  aoai13aa1n02x5               g055(.a(new_n111), .b(new_n106), .c(new_n134), .d(new_n133), .o1(new_n151));
  nona23aa1n02x4               g056(.a(new_n151), .b(new_n139), .c(new_n117), .d(new_n103), .out0(new_n152));
  norp02aa1n02x5               g057(.a(\b[10] ), .b(\a[11] ), .o1(new_n153));
  nanp02aa1n02x5               g058(.a(\b[10] ), .b(\a[11] ), .o1(new_n154));
  norp02aa1n02x5               g059(.a(\b[11] ), .b(\a[12] ), .o1(new_n155));
  nanp02aa1n02x5               g060(.a(\b[11] ), .b(\a[12] ), .o1(new_n156));
  nona23aa1n02x4               g061(.a(new_n156), .b(new_n154), .c(new_n153), .d(new_n155), .out0(new_n157));
  norb03aa1n02x5               g062(.a(new_n128), .b(new_n157), .c(new_n99), .out0(new_n158));
  160nm_ficinv00aa1n08x5       g063(.clk(new_n158), .clkout(new_n159));
  nano23aa1n02x4               g064(.a(new_n153), .b(new_n155), .c(new_n156), .d(new_n154), .out0(new_n160));
  aoi012aa1n02x5               g065(.a(new_n155), .b(new_n153), .c(new_n156), .o1(new_n161));
  aobi12aa1n02x5               g066(.a(new_n161), .b(new_n160), .c(new_n144), .out0(new_n162));
  aoai13aa1n02x5               g067(.a(new_n162), .b(new_n159), .c(new_n152), .d(new_n141), .o1(new_n163));
  xorb03aa1n02x5               g068(.a(new_n163), .b(\b[12] ), .c(\a[13] ), .out0(\s[13] ));
  160nm_ficinv00aa1n08x5       g069(.clk(\a[13] ), .clkout(new_n165));
  160nm_ficinv00aa1n08x5       g070(.clk(\b[12] ), .clkout(new_n166));
  oaoi03aa1n02x5               g071(.a(new_n165), .b(new_n166), .c(new_n163), .o1(new_n167));
  xnrb03aa1n02x5               g072(.a(new_n167), .b(\b[13] ), .c(\a[14] ), .out0(\s[14] ));
  aoai13aa1n02x5               g073(.a(new_n158), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n169));
  norp02aa1n02x5               g074(.a(\b[12] ), .b(\a[13] ), .o1(new_n170));
  nanp02aa1n02x5               g075(.a(\b[12] ), .b(\a[13] ), .o1(new_n171));
  norp02aa1n02x5               g076(.a(\b[13] ), .b(\a[14] ), .o1(new_n172));
  nanp02aa1n02x5               g077(.a(\b[13] ), .b(\a[14] ), .o1(new_n173));
  nona23aa1n02x4               g078(.a(new_n173), .b(new_n171), .c(new_n170), .d(new_n172), .out0(new_n174));
  aoai13aa1n02x5               g079(.a(new_n173), .b(new_n172), .c(new_n165), .d(new_n166), .o1(new_n175));
  aoai13aa1n02x5               g080(.a(new_n175), .b(new_n174), .c(new_n169), .d(new_n162), .o1(new_n176));
  xorb03aa1n02x5               g081(.a(new_n176), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  norp02aa1n02x5               g082(.a(\b[14] ), .b(\a[15] ), .o1(new_n178));
  nanp02aa1n02x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  nanb02aa1n02x5               g084(.a(new_n178), .b(new_n179), .out0(new_n180));
  160nm_ficinv00aa1n08x5       g085(.clk(new_n180), .clkout(new_n181));
  norp02aa1n02x5               g086(.a(\b[15] ), .b(\a[16] ), .o1(new_n182));
  nanp02aa1n02x5               g087(.a(\b[15] ), .b(\a[16] ), .o1(new_n183));
  nanb02aa1n02x5               g088(.a(new_n182), .b(new_n183), .out0(new_n184));
  160nm_ficinv00aa1n08x5       g089(.clk(new_n184), .clkout(new_n185));
  aoi112aa1n02x5               g090(.a(new_n185), .b(new_n178), .c(new_n176), .d(new_n181), .o1(new_n186));
  160nm_ficinv00aa1n08x5       g091(.clk(new_n178), .clkout(new_n187));
  nano23aa1n02x4               g092(.a(new_n170), .b(new_n172), .c(new_n173), .d(new_n171), .out0(new_n188));
  160nm_ficinv00aa1n08x5       g093(.clk(new_n175), .clkout(new_n189));
  aoai13aa1n02x5               g094(.a(new_n181), .b(new_n189), .c(new_n163), .d(new_n188), .o1(new_n190));
  aoi012aa1n02x5               g095(.a(new_n184), .b(new_n190), .c(new_n187), .o1(new_n191));
  norp02aa1n02x5               g096(.a(new_n191), .b(new_n186), .o1(\s[16] ));
  nona23aa1n02x4               g097(.a(new_n183), .b(new_n179), .c(new_n178), .d(new_n182), .out0(new_n193));
  nona23aa1n02x4               g098(.a(new_n188), .b(new_n146), .c(new_n193), .d(new_n157), .out0(new_n194));
  oai012aa1n02x5               g099(.a(new_n161), .b(new_n157), .c(new_n143), .o1(new_n195));
  norp02aa1n02x5               g100(.a(new_n193), .b(new_n174), .o1(new_n196));
  aoi012aa1n02x5               g101(.a(new_n182), .b(new_n178), .c(new_n183), .o1(new_n197));
  oai012aa1n02x5               g102(.a(new_n197), .b(new_n193), .c(new_n175), .o1(new_n198));
  aoi012aa1n02x5               g103(.a(new_n198), .b(new_n195), .c(new_n196), .o1(new_n199));
  aoai13aa1n02x5               g104(.a(new_n199), .b(new_n194), .c(new_n152), .d(new_n141), .o1(new_n200));
  xorb03aa1n02x5               g105(.a(new_n200), .b(\b[16] ), .c(\a[17] ), .out0(\s[17] ));
  160nm_ficinv00aa1n08x5       g106(.clk(\a[18] ), .clkout(new_n202));
  160nm_ficinv00aa1n08x5       g107(.clk(\a[17] ), .clkout(new_n203));
  160nm_ficinv00aa1n08x5       g108(.clk(\b[16] ), .clkout(new_n204));
  oaoi03aa1n02x5               g109(.a(new_n203), .b(new_n204), .c(new_n200), .o1(new_n205));
  xorb03aa1n02x5               g110(.a(new_n205), .b(\b[17] ), .c(new_n202), .out0(\s[18] ));
  nona22aa1n02x4               g111(.a(new_n188), .b(new_n184), .c(new_n180), .out0(new_n207));
  nano22aa1n02x4               g112(.a(new_n207), .b(new_n146), .c(new_n160), .out0(new_n208));
  aoai13aa1n02x5               g113(.a(new_n208), .b(new_n127), .c(new_n112), .d(new_n124), .o1(new_n209));
  xroi22aa1d04x5               g114(.a(new_n203), .b(\b[16] ), .c(new_n202), .d(\b[17] ), .out0(new_n210));
  160nm_ficinv00aa1n08x5       g115(.clk(new_n210), .clkout(new_n211));
  oai022aa1n02x5               g116(.a(\a[17] ), .b(\b[16] ), .c(\b[17] ), .d(\a[18] ), .o1(new_n212));
  oaib12aa1n02x5               g117(.a(new_n212), .b(new_n202), .c(\b[17] ), .out0(new_n213));
  aoai13aa1n02x5               g118(.a(new_n213), .b(new_n211), .c(new_n209), .d(new_n199), .o1(new_n214));
  xorb03aa1n02x5               g119(.a(new_n214), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g120(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  norp02aa1n02x5               g121(.a(\b[18] ), .b(\a[19] ), .o1(new_n217));
  nanp02aa1n02x5               g122(.a(\b[18] ), .b(\a[19] ), .o1(new_n218));
  nanb02aa1n02x5               g123(.a(new_n217), .b(new_n218), .out0(new_n219));
  160nm_ficinv00aa1n08x5       g124(.clk(new_n219), .clkout(new_n220));
  norp02aa1n02x5               g125(.a(\b[19] ), .b(\a[20] ), .o1(new_n221));
  nanp02aa1n02x5               g126(.a(\b[19] ), .b(\a[20] ), .o1(new_n222));
  nanb02aa1n02x5               g127(.a(new_n221), .b(new_n222), .out0(new_n223));
  160nm_ficinv00aa1n08x5       g128(.clk(new_n223), .clkout(new_n224));
  aoi112aa1n02x5               g129(.a(new_n217), .b(new_n224), .c(new_n214), .d(new_n220), .o1(new_n225));
  160nm_ficinv00aa1n08x5       g130(.clk(new_n217), .clkout(new_n226));
  nanp02aa1n02x5               g131(.a(new_n204), .b(new_n203), .o1(new_n227));
  oaoi03aa1n02x5               g132(.a(\a[18] ), .b(\b[17] ), .c(new_n227), .o1(new_n228));
  aoai13aa1n02x5               g133(.a(new_n220), .b(new_n228), .c(new_n200), .d(new_n210), .o1(new_n229));
  aoi012aa1n02x5               g134(.a(new_n223), .b(new_n229), .c(new_n226), .o1(new_n230));
  norp02aa1n02x5               g135(.a(new_n230), .b(new_n225), .o1(\s[20] ));
  nona23aa1n02x4               g136(.a(new_n222), .b(new_n218), .c(new_n217), .d(new_n221), .out0(new_n232));
  norb02aa1n02x5               g137(.a(new_n210), .b(new_n232), .out0(new_n233));
  160nm_ficinv00aa1n08x5       g138(.clk(new_n233), .clkout(new_n234));
  nano23aa1n02x4               g139(.a(new_n217), .b(new_n221), .c(new_n222), .d(new_n218), .out0(new_n235));
  oaoi03aa1n02x5               g140(.a(\a[20] ), .b(\b[19] ), .c(new_n226), .o1(new_n236));
  aoi012aa1n02x5               g141(.a(new_n236), .b(new_n235), .c(new_n228), .o1(new_n237));
  aoai13aa1n02x5               g142(.a(new_n237), .b(new_n234), .c(new_n209), .d(new_n199), .o1(new_n238));
  xorb03aa1n02x5               g143(.a(new_n238), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g144(.a(\b[20] ), .b(\a[21] ), .o1(new_n240));
  xnrc02aa1n02x5               g145(.a(\b[20] ), .b(\a[21] ), .out0(new_n241));
  160nm_ficinv00aa1n08x5       g146(.clk(new_n241), .clkout(new_n242));
  norp02aa1n02x5               g147(.a(\b[21] ), .b(\a[22] ), .o1(new_n243));
  nanp02aa1n02x5               g148(.a(\b[21] ), .b(\a[22] ), .o1(new_n244));
  nanb02aa1n02x5               g149(.a(new_n243), .b(new_n244), .out0(new_n245));
  160nm_ficinv00aa1n08x5       g150(.clk(new_n245), .clkout(new_n246));
  aoi112aa1n02x5               g151(.a(new_n240), .b(new_n246), .c(new_n238), .d(new_n242), .o1(new_n247));
  160nm_ficinv00aa1n08x5       g152(.clk(new_n240), .clkout(new_n248));
  oabi12aa1n02x5               g153(.a(new_n236), .b(new_n232), .c(new_n213), .out0(new_n249));
  aoai13aa1n02x5               g154(.a(new_n242), .b(new_n249), .c(new_n200), .d(new_n233), .o1(new_n250));
  aoi012aa1n02x5               g155(.a(new_n245), .b(new_n250), .c(new_n248), .o1(new_n251));
  norp02aa1n02x5               g156(.a(new_n251), .b(new_n247), .o1(\s[22] ));
  norp02aa1n02x5               g157(.a(new_n241), .b(new_n245), .o1(new_n253));
  nanp03aa1n02x5               g158(.a(new_n210), .b(new_n253), .c(new_n235), .o1(new_n254));
  oai012aa1n02x5               g159(.a(new_n244), .b(new_n243), .c(new_n240), .o1(new_n255));
  aobi12aa1n02x5               g160(.a(new_n255), .b(new_n249), .c(new_n253), .out0(new_n256));
  aoai13aa1n02x5               g161(.a(new_n256), .b(new_n254), .c(new_n209), .d(new_n199), .o1(new_n257));
  xorb03aa1n02x5               g162(.a(new_n257), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  norp02aa1n02x5               g163(.a(\b[22] ), .b(\a[23] ), .o1(new_n259));
  nanp02aa1n02x5               g164(.a(\b[22] ), .b(\a[23] ), .o1(new_n260));
  nanb02aa1n02x5               g165(.a(new_n259), .b(new_n260), .out0(new_n261));
  160nm_ficinv00aa1n08x5       g166(.clk(new_n261), .clkout(new_n262));
  norp02aa1n02x5               g167(.a(\b[23] ), .b(\a[24] ), .o1(new_n263));
  nanp02aa1n02x5               g168(.a(\b[23] ), .b(\a[24] ), .o1(new_n264));
  nanb02aa1n02x5               g169(.a(new_n263), .b(new_n264), .out0(new_n265));
  160nm_ficinv00aa1n08x5       g170(.clk(new_n265), .clkout(new_n266));
  aoi112aa1n02x5               g171(.a(new_n259), .b(new_n266), .c(new_n257), .d(new_n262), .o1(new_n267));
  160nm_ficinv00aa1n08x5       g172(.clk(new_n259), .clkout(new_n268));
  160nm_ficinv00aa1n08x5       g173(.clk(new_n254), .clkout(new_n269));
  160nm_ficinv00aa1n08x5       g174(.clk(new_n256), .clkout(new_n270));
  aoai13aa1n02x5               g175(.a(new_n262), .b(new_n270), .c(new_n200), .d(new_n269), .o1(new_n271));
  aoi012aa1n02x5               g176(.a(new_n265), .b(new_n271), .c(new_n268), .o1(new_n272));
  norp02aa1n02x5               g177(.a(new_n272), .b(new_n267), .o1(\s[24] ));
  nona23aa1n02x4               g178(.a(new_n264), .b(new_n260), .c(new_n259), .d(new_n263), .out0(new_n274));
  160nm_ficinv00aa1n08x5       g179(.clk(new_n274), .clkout(new_n275));
  nano32aa1n02x4               g180(.a(new_n211), .b(new_n275), .c(new_n235), .d(new_n253), .out0(new_n276));
  160nm_ficinv00aa1n08x5       g181(.clk(new_n276), .clkout(new_n277));
  oaoi03aa1n02x5               g182(.a(\a[24] ), .b(\b[23] ), .c(new_n268), .o1(new_n278));
  oabi12aa1n02x5               g183(.a(new_n278), .b(new_n274), .c(new_n255), .out0(new_n279));
  aoi013aa1n02x4               g184(.a(new_n279), .b(new_n249), .c(new_n253), .d(new_n275), .o1(new_n280));
  aoai13aa1n02x5               g185(.a(new_n280), .b(new_n277), .c(new_n209), .d(new_n199), .o1(new_n281));
  xorb03aa1n02x5               g186(.a(new_n281), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g187(.a(\b[24] ), .b(\a[25] ), .o1(new_n283));
  xorc02aa1n02x5               g188(.a(\a[25] ), .b(\b[24] ), .out0(new_n284));
  xorc02aa1n02x5               g189(.a(\a[26] ), .b(\b[25] ), .out0(new_n285));
  aoi112aa1n02x5               g190(.a(new_n283), .b(new_n285), .c(new_n281), .d(new_n284), .o1(new_n286));
  160nm_ficinv00aa1n08x5       g191(.clk(new_n283), .clkout(new_n287));
  160nm_ficinv00aa1n08x5       g192(.clk(new_n280), .clkout(new_n288));
  aoai13aa1n02x5               g193(.a(new_n284), .b(new_n288), .c(new_n200), .d(new_n276), .o1(new_n289));
  160nm_ficinv00aa1n08x5       g194(.clk(new_n285), .clkout(new_n290));
  aoi012aa1n02x5               g195(.a(new_n290), .b(new_n289), .c(new_n287), .o1(new_n291));
  norp02aa1n02x5               g196(.a(new_n291), .b(new_n286), .o1(\s[26] ));
  oabi12aa1n02x5               g197(.a(new_n198), .b(new_n162), .c(new_n207), .out0(new_n293));
  and002aa1n02x5               g198(.a(new_n285), .b(new_n284), .o(new_n294));
  nano22aa1n02x4               g199(.a(new_n254), .b(new_n294), .c(new_n275), .out0(new_n295));
  aoai13aa1n02x5               g200(.a(new_n295), .b(new_n293), .c(new_n142), .d(new_n208), .o1(new_n296));
  nano22aa1n02x4               g201(.a(new_n237), .b(new_n253), .c(new_n275), .out0(new_n297));
  oao003aa1n02x5               g202(.a(\a[26] ), .b(\b[25] ), .c(new_n287), .carry(new_n298));
  160nm_ficinv00aa1n08x5       g203(.clk(new_n298), .clkout(new_n299));
  oaoi13aa1n02x5               g204(.a(new_n299), .b(new_n294), .c(new_n297), .d(new_n279), .o1(new_n300));
  norp02aa1n02x5               g205(.a(\b[26] ), .b(\a[27] ), .o1(new_n301));
  and002aa1n02x5               g206(.a(\b[26] ), .b(\a[27] ), .o(new_n302));
  norp02aa1n02x5               g207(.a(new_n302), .b(new_n301), .o1(new_n303));
  xnbna2aa1n03x5               g208(.a(new_n303), .b(new_n296), .c(new_n300), .out0(\s[27] ));
  160nm_ficinv00aa1n08x5       g209(.clk(new_n301), .clkout(new_n305));
  xnrc02aa1n02x5               g210(.a(\b[27] ), .b(\a[28] ), .out0(new_n306));
  nona32aa1n02x4               g211(.a(new_n249), .b(new_n274), .c(new_n245), .d(new_n241), .out0(new_n307));
  160nm_ficinv00aa1n08x5       g212(.clk(new_n279), .clkout(new_n308));
  160nm_ficinv00aa1n08x5       g213(.clk(new_n294), .clkout(new_n309));
  aoai13aa1n02x5               g214(.a(new_n298), .b(new_n309), .c(new_n307), .d(new_n308), .o1(new_n310));
  160nm_ficinv00aa1n08x5       g215(.clk(new_n302), .clkout(new_n311));
  aoai13aa1n02x5               g216(.a(new_n311), .b(new_n310), .c(new_n200), .d(new_n295), .o1(new_n312));
  aoi012aa1n02x5               g217(.a(new_n306), .b(new_n312), .c(new_n305), .o1(new_n313));
  aoi012aa1n02x5               g218(.a(new_n302), .b(new_n296), .c(new_n300), .o1(new_n314));
  nano22aa1n02x4               g219(.a(new_n314), .b(new_n305), .c(new_n306), .out0(new_n315));
  norp02aa1n02x5               g220(.a(new_n313), .b(new_n315), .o1(\s[28] ));
  nano22aa1n02x4               g221(.a(new_n306), .b(new_n311), .c(new_n305), .out0(new_n317));
  aoai13aa1n02x5               g222(.a(new_n317), .b(new_n310), .c(new_n200), .d(new_n295), .o1(new_n318));
  oao003aa1n02x5               g223(.a(\a[28] ), .b(\b[27] ), .c(new_n305), .carry(new_n319));
  xnrc02aa1n02x5               g224(.a(\b[28] ), .b(\a[29] ), .out0(new_n320));
  aoi012aa1n02x5               g225(.a(new_n320), .b(new_n318), .c(new_n319), .o1(new_n321));
  160nm_ficinv00aa1n08x5       g226(.clk(new_n317), .clkout(new_n322));
  aoi012aa1n02x5               g227(.a(new_n322), .b(new_n296), .c(new_n300), .o1(new_n323));
  nano22aa1n02x4               g228(.a(new_n323), .b(new_n319), .c(new_n320), .out0(new_n324));
  norp02aa1n02x5               g229(.a(new_n321), .b(new_n324), .o1(\s[29] ));
  xorb03aa1n02x5               g230(.a(new_n108), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  norb03aa1n02x5               g231(.a(new_n303), .b(new_n320), .c(new_n306), .out0(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n310), .c(new_n200), .d(new_n295), .o1(new_n328));
  oao003aa1n02x5               g233(.a(\a[29] ), .b(\b[28] ), .c(new_n319), .carry(new_n329));
  xnrc02aa1n02x5               g234(.a(\b[29] ), .b(\a[30] ), .out0(new_n330));
  aoi012aa1n02x5               g235(.a(new_n330), .b(new_n328), .c(new_n329), .o1(new_n331));
  160nm_ficinv00aa1n08x5       g236(.clk(new_n327), .clkout(new_n332));
  aoi012aa1n02x5               g237(.a(new_n332), .b(new_n296), .c(new_n300), .o1(new_n333));
  nano22aa1n02x4               g238(.a(new_n333), .b(new_n329), .c(new_n330), .out0(new_n334));
  norp02aa1n02x5               g239(.a(new_n331), .b(new_n334), .o1(\s[30] ));
  xnrc02aa1n02x5               g240(.a(\b[30] ), .b(\a[31] ), .out0(new_n336));
  norb03aa1n02x5               g241(.a(new_n317), .b(new_n330), .c(new_n320), .out0(new_n337));
  160nm_ficinv00aa1n08x5       g242(.clk(new_n337), .clkout(new_n338));
  aoi012aa1n02x5               g243(.a(new_n338), .b(new_n296), .c(new_n300), .o1(new_n339));
  oao003aa1n02x5               g244(.a(\a[30] ), .b(\b[29] ), .c(new_n329), .carry(new_n340));
  nano22aa1n02x4               g245(.a(new_n339), .b(new_n336), .c(new_n340), .out0(new_n341));
  aoai13aa1n02x5               g246(.a(new_n337), .b(new_n310), .c(new_n200), .d(new_n295), .o1(new_n342));
  aoi012aa1n02x5               g247(.a(new_n336), .b(new_n342), .c(new_n340), .o1(new_n343));
  norp02aa1n02x5               g248(.a(new_n343), .b(new_n341), .o1(\s[31] ));
  xnbna2aa1n03x5               g249(.a(new_n132), .b(new_n134), .c(new_n133), .out0(\s[3] ));
  oaoi03aa1n02x5               g250(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n346));
  xorb03aa1n02x5               g251(.a(new_n346), .b(\b[3] ), .c(\a[4] ), .out0(\s[4] ));
  xobna2aa1n03x5               g252(.a(new_n123), .b(new_n151), .c(new_n131), .out0(\s[5] ));
  aoai13aa1n02x5               g253(.a(new_n122), .b(new_n121), .c(new_n151), .d(new_n131), .o1(new_n349));
  xnrc02aa1n02x5               g254(.a(new_n349), .b(new_n120), .out0(\s[6] ));
  aobi12aa1n02x5               g255(.a(new_n125), .b(new_n112), .c(new_n139), .out0(new_n351));
  xnrb03aa1n02x5               g256(.a(new_n351), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  oaoi03aa1n02x5               g257(.a(\a[7] ), .b(\b[6] ), .c(new_n351), .o1(new_n353));
  xorb03aa1n02x5               g258(.a(new_n353), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  xnbna2aa1n03x5               g259(.a(new_n128), .b(new_n152), .c(new_n141), .out0(\s[9] ));
endmodule


