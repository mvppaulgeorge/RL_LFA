// Benchmark "adder" written by ABC on Wed Jul 17 19:41:10 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n133, new_n134, new_n135, new_n136, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n158, new_n159, new_n160, new_n161, new_n162, new_n164,
    new_n165, new_n166, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n187, new_n188,
    new_n189, new_n190, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n305, new_n306, new_n307, new_n310, new_n311, new_n312,
    new_n313, new_n315, new_n317, new_n319;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1d24x5               g001(.a(\b[8] ), .b(\a[9] ), .o1(new_n97));
  inv000aa1d42x5               g002(.a(new_n97), .o1(new_n98));
  and002aa1n12x5               g003(.a(\b[3] ), .b(\a[4] ), .o(new_n99));
  inv040aa1d32x5               g004(.a(\a[3] ), .o1(new_n100));
  inv040aa1d28x5               g005(.a(\b[2] ), .o1(new_n101));
  nor042aa1n02x5               g006(.a(\b[3] ), .b(\a[4] ), .o1(new_n102));
  aoi112aa1n06x5               g007(.a(new_n99), .b(new_n102), .c(new_n100), .d(new_n101), .o1(new_n103));
  tech160nm_finand02aa1n03p5x5 g008(.a(new_n101), .b(new_n100), .o1(new_n104));
  tech160nm_finand02aa1n03p5x5 g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nand22aa1n03x5               g010(.a(new_n104), .b(new_n105), .o1(new_n106));
  nand42aa1n03x5               g011(.a(\b[1] ), .b(\a[2] ), .o1(new_n107));
  nor042aa1d18x5               g012(.a(\b[1] ), .b(\a[2] ), .o1(new_n108));
  nand02aa1n16x5               g013(.a(\b[0] ), .b(\a[1] ), .o1(new_n109));
  oai012aa1n12x5               g014(.a(new_n107), .b(new_n108), .c(new_n109), .o1(new_n110));
  oaoi13aa1n12x5               g015(.a(new_n99), .b(new_n103), .c(new_n110), .d(new_n106), .o1(new_n111));
  nanp02aa1n02x5               g016(.a(\b[4] ), .b(\a[5] ), .o1(new_n112));
  nor042aa1n04x5               g017(.a(\b[4] ), .b(\a[5] ), .o1(new_n113));
  nor002aa1n03x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand42aa1n08x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  norb03aa1n03x5               g020(.a(new_n115), .b(new_n113), .c(new_n114), .out0(new_n116));
  nor002aa1d32x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nanp02aa1n04x5               g022(.a(\b[7] ), .b(\a[8] ), .o1(new_n118));
  nanp02aa1n04x5               g023(.a(\b[6] ), .b(\a[7] ), .o1(new_n119));
  nor002aa1n12x5               g024(.a(\b[6] ), .b(\a[7] ), .o1(new_n120));
  nona23aa1n09x5               g025(.a(new_n119), .b(new_n118), .c(new_n120), .d(new_n117), .out0(new_n121));
  nano22aa1n03x7               g026(.a(new_n121), .b(new_n116), .c(new_n112), .out0(new_n122));
  oai012aa1n02x7               g027(.a(new_n115), .b(new_n114), .c(new_n113), .o1(new_n123));
  aoi012aa1n12x5               g028(.a(new_n117), .b(new_n120), .c(new_n118), .o1(new_n124));
  tech160nm_fioai012aa1n03p5x5 g029(.a(new_n124), .b(new_n121), .c(new_n123), .o1(new_n125));
  nanp02aa1n09x5               g030(.a(\b[8] ), .b(\a[9] ), .o1(new_n126));
  norb02aa1n02x5               g031(.a(new_n126), .b(new_n97), .out0(new_n127));
  aoai13aa1n02x5               g032(.a(new_n127), .b(new_n125), .c(new_n111), .d(new_n122), .o1(new_n128));
  nor042aa1n06x5               g033(.a(\b[9] ), .b(\a[10] ), .o1(new_n129));
  nand42aa1n20x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  norb02aa1n02x5               g035(.a(new_n130), .b(new_n129), .out0(new_n131));
  xnbna2aa1n03x5               g036(.a(new_n131), .b(new_n128), .c(new_n98), .out0(\s[10] ));
  nor002aa1d32x5               g037(.a(\b[10] ), .b(\a[11] ), .o1(new_n133));
  nand42aa1d28x5               g038(.a(\b[10] ), .b(\a[11] ), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(new_n135));
  nona22aa1n02x4               g040(.a(new_n128), .b(new_n129), .c(new_n97), .out0(new_n136));
  xobna2aa1n03x5               g041(.a(new_n135), .b(new_n136), .c(new_n130), .out0(\s[11] ));
  inv000aa1d42x5               g042(.a(new_n133), .o1(new_n138));
  nanp03aa1n02x5               g043(.a(new_n136), .b(new_n130), .c(new_n135), .o1(new_n139));
  nor002aa1n12x5               g044(.a(\b[11] ), .b(\a[12] ), .o1(new_n140));
  nand42aa1d28x5               g045(.a(\b[11] ), .b(\a[12] ), .o1(new_n141));
  norb02aa1n02x5               g046(.a(new_n141), .b(new_n140), .out0(new_n142));
  xnbna2aa1n03x5               g047(.a(new_n142), .b(new_n139), .c(new_n138), .out0(\s[12] ));
  nano23aa1n09x5               g048(.a(new_n133), .b(new_n140), .c(new_n141), .d(new_n134), .out0(new_n144));
  nano23aa1n09x5               g049(.a(new_n97), .b(new_n129), .c(new_n130), .d(new_n126), .out0(new_n145));
  nand22aa1n09x5               g050(.a(new_n145), .b(new_n144), .o1(new_n146));
  inv000aa1d42x5               g051(.a(new_n146), .o1(new_n147));
  aoai13aa1n02x5               g052(.a(new_n147), .b(new_n125), .c(new_n111), .d(new_n122), .o1(new_n148));
  nona23aa1d18x5               g053(.a(new_n141), .b(new_n134), .c(new_n133), .d(new_n140), .out0(new_n149));
  oaih12aa1n06x5               g054(.a(new_n130), .b(new_n129), .c(new_n97), .o1(new_n150));
  tech160nm_fiaoi012aa1n03p5x5 g055(.a(new_n140), .b(new_n133), .c(new_n141), .o1(new_n151));
  oai012aa1n18x5               g056(.a(new_n151), .b(new_n149), .c(new_n150), .o1(new_n152));
  inv000aa1d42x5               g057(.a(new_n152), .o1(new_n153));
  nor042aa1n04x5               g058(.a(\b[12] ), .b(\a[13] ), .o1(new_n154));
  nand02aa1n06x5               g059(.a(\b[12] ), .b(\a[13] ), .o1(new_n155));
  norb02aa1n03x5               g060(.a(new_n155), .b(new_n154), .out0(new_n156));
  xnbna2aa1n03x5               g061(.a(new_n156), .b(new_n148), .c(new_n153), .out0(\s[13] ));
  nanp02aa1n02x5               g062(.a(new_n148), .b(new_n153), .o1(new_n158));
  aoi012aa1n02x5               g063(.a(new_n154), .b(new_n158), .c(new_n155), .o1(new_n159));
  norp02aa1n04x5               g064(.a(\b[13] ), .b(\a[14] ), .o1(new_n160));
  nand42aa1n06x5               g065(.a(\b[13] ), .b(\a[14] ), .o1(new_n161));
  norb02aa1n02x7               g066(.a(new_n161), .b(new_n160), .out0(new_n162));
  xnrc02aa1n02x5               g067(.a(new_n159), .b(new_n162), .out0(\s[14] ));
  nona23aa1n09x5               g068(.a(new_n161), .b(new_n155), .c(new_n154), .d(new_n160), .out0(new_n164));
  aoi012aa1n03x5               g069(.a(new_n160), .b(new_n154), .c(new_n161), .o1(new_n165));
  aoai13aa1n04x5               g070(.a(new_n165), .b(new_n164), .c(new_n148), .d(new_n153), .o1(new_n166));
  xorb03aa1n02x5               g071(.a(new_n166), .b(\b[14] ), .c(\a[15] ), .out0(\s[15] ));
  nor022aa1n06x5               g072(.a(\b[14] ), .b(\a[15] ), .o1(new_n168));
  tech160nm_finand02aa1n03p5x5 g073(.a(\b[14] ), .b(\a[15] ), .o1(new_n169));
  nor022aa1n06x5               g074(.a(\b[15] ), .b(\a[16] ), .o1(new_n170));
  nand42aa1n03x5               g075(.a(\b[15] ), .b(\a[16] ), .o1(new_n171));
  nanb02aa1n02x5               g076(.a(new_n170), .b(new_n171), .out0(new_n172));
  inv000aa1d42x5               g077(.a(new_n172), .o1(new_n173));
  aoi112aa1n02x5               g078(.a(new_n173), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n174));
  aoai13aa1n02x5               g079(.a(new_n173), .b(new_n168), .c(new_n166), .d(new_n169), .o1(new_n175));
  norb02aa1n02x5               g080(.a(new_n175), .b(new_n174), .out0(\s[16] ));
  nano23aa1n03x5               g081(.a(new_n168), .b(new_n170), .c(new_n171), .d(new_n169), .out0(new_n177));
  nano32aa1n03x7               g082(.a(new_n146), .b(new_n177), .c(new_n156), .d(new_n162), .out0(new_n178));
  aoai13aa1n12x5               g083(.a(new_n178), .b(new_n125), .c(new_n111), .d(new_n122), .o1(new_n179));
  nona23aa1n03x5               g084(.a(new_n171), .b(new_n169), .c(new_n168), .d(new_n170), .out0(new_n180));
  norp02aa1n03x5               g085(.a(new_n180), .b(new_n164), .o1(new_n181));
  norp02aa1n02x5               g086(.a(new_n180), .b(new_n165), .o1(new_n182));
  oa0012aa1n02x5               g087(.a(new_n171), .b(new_n170), .c(new_n168), .o(new_n183));
  aoi112aa1n09x5               g088(.a(new_n183), .b(new_n182), .c(new_n152), .d(new_n181), .o1(new_n184));
  xorc02aa1n02x5               g089(.a(\a[17] ), .b(\b[16] ), .out0(new_n185));
  xnbna2aa1n03x5               g090(.a(new_n185), .b(new_n179), .c(new_n184), .out0(\s[17] ));
  inv040aa1d32x5               g091(.a(\a[18] ), .o1(new_n187));
  nand02aa1d08x5               g092(.a(new_n179), .b(new_n184), .o1(new_n188));
  norp02aa1n02x5               g093(.a(\b[16] ), .b(\a[17] ), .o1(new_n189));
  tech160nm_fiaoi012aa1n05x5   g094(.a(new_n189), .b(new_n188), .c(new_n185), .o1(new_n190));
  xorb03aa1n02x5               g095(.a(new_n190), .b(\b[17] ), .c(new_n187), .out0(\s[18] ));
  inv000aa1d42x5               g096(.a(\a[17] ), .o1(new_n192));
  xroi22aa1d06x4               g097(.a(new_n192), .b(\b[16] ), .c(new_n187), .d(\b[17] ), .out0(new_n193));
  inv000aa1d42x5               g098(.a(new_n193), .o1(new_n194));
  inv000aa1d42x5               g099(.a(\b[17] ), .o1(new_n195));
  oao003aa1n02x5               g100(.a(new_n187), .b(new_n195), .c(new_n189), .carry(new_n196));
  inv000aa1d42x5               g101(.a(new_n196), .o1(new_n197));
  aoai13aa1n06x5               g102(.a(new_n197), .b(new_n194), .c(new_n179), .d(new_n184), .o1(new_n198));
  xorb03aa1n02x5               g103(.a(new_n198), .b(\b[18] ), .c(\a[19] ), .out0(\s[19] ));
  xnrc02aa1n02x5               g104(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nor042aa1n03x5               g105(.a(\b[18] ), .b(\a[19] ), .o1(new_n201));
  nand22aa1n04x5               g106(.a(\b[18] ), .b(\a[19] ), .o1(new_n202));
  nor042aa1n03x5               g107(.a(\b[19] ), .b(\a[20] ), .o1(new_n203));
  nand02aa1n03x5               g108(.a(\b[19] ), .b(\a[20] ), .o1(new_n204));
  norb02aa1n06x4               g109(.a(new_n204), .b(new_n203), .out0(new_n205));
  aoi112aa1n02x5               g110(.a(new_n205), .b(new_n201), .c(new_n198), .d(new_n202), .o1(new_n206));
  aoai13aa1n03x5               g111(.a(new_n205), .b(new_n201), .c(new_n198), .d(new_n202), .o1(new_n207));
  norb02aa1n03x4               g112(.a(new_n207), .b(new_n206), .out0(\s[20] ));
  nano23aa1n02x4               g113(.a(new_n201), .b(new_n203), .c(new_n204), .d(new_n202), .out0(new_n209));
  nand02aa1n02x5               g114(.a(new_n193), .b(new_n209), .o1(new_n210));
  aoi112aa1n02x5               g115(.a(\b[18] ), .b(\a[19] ), .c(\a[20] ), .d(\b[19] ), .o1(new_n211));
  norp02aa1n02x5               g116(.a(\b[17] ), .b(\a[18] ), .o1(new_n212));
  norb02aa1n06x4               g117(.a(new_n202), .b(new_n201), .out0(new_n213));
  aoi112aa1n03x5               g118(.a(\b[16] ), .b(\a[17] ), .c(\a[18] ), .d(\b[17] ), .o1(new_n214));
  oai112aa1n06x5               g119(.a(new_n205), .b(new_n213), .c(new_n214), .d(new_n212), .o1(new_n215));
  nona22aa1n12x5               g120(.a(new_n215), .b(new_n211), .c(new_n203), .out0(new_n216));
  inv000aa1d42x5               g121(.a(new_n216), .o1(new_n217));
  aoai13aa1n04x5               g122(.a(new_n217), .b(new_n210), .c(new_n179), .d(new_n184), .o1(new_n218));
  xorb03aa1n02x5               g123(.a(new_n218), .b(\b[20] ), .c(\a[21] ), .out0(\s[21] ));
  norp02aa1n02x5               g124(.a(\b[20] ), .b(\a[21] ), .o1(new_n220));
  xnrc02aa1n12x5               g125(.a(\b[20] ), .b(\a[21] ), .out0(new_n221));
  inv000aa1d42x5               g126(.a(new_n221), .o1(new_n222));
  xnrc02aa1n12x5               g127(.a(\b[21] ), .b(\a[22] ), .out0(new_n223));
  inv000aa1d42x5               g128(.a(new_n223), .o1(new_n224));
  aoi112aa1n03x5               g129(.a(new_n220), .b(new_n224), .c(new_n218), .d(new_n222), .o1(new_n225));
  aoai13aa1n03x5               g130(.a(new_n224), .b(new_n220), .c(new_n218), .d(new_n222), .o1(new_n226));
  norb02aa1n02x7               g131(.a(new_n226), .b(new_n225), .out0(\s[22] ));
  tech160nm_finor002aa1n03p5x5 g132(.a(new_n223), .b(new_n221), .o1(new_n228));
  nand23aa1n03x5               g133(.a(new_n193), .b(new_n228), .c(new_n209), .o1(new_n229));
  inv000aa1n02x5               g134(.a(new_n220), .o1(new_n230));
  oaoi03aa1n02x5               g135(.a(\a[22] ), .b(\b[21] ), .c(new_n230), .o1(new_n231));
  aoi012aa1n02x5               g136(.a(new_n231), .b(new_n216), .c(new_n228), .o1(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n229), .c(new_n179), .d(new_n184), .o1(new_n233));
  xorb03aa1n02x5               g138(.a(new_n233), .b(\b[22] ), .c(\a[23] ), .out0(\s[23] ));
  nor042aa1n03x5               g139(.a(\b[22] ), .b(\a[23] ), .o1(new_n235));
  nand42aa1n02x5               g140(.a(\b[22] ), .b(\a[23] ), .o1(new_n236));
  nor042aa1n04x5               g141(.a(\b[23] ), .b(\a[24] ), .o1(new_n237));
  nanp02aa1n02x5               g142(.a(\b[23] ), .b(\a[24] ), .o1(new_n238));
  norb02aa1n02x5               g143(.a(new_n238), .b(new_n237), .out0(new_n239));
  aoi112aa1n02x5               g144(.a(new_n235), .b(new_n239), .c(new_n233), .d(new_n236), .o1(new_n240));
  aoai13aa1n03x5               g145(.a(new_n239), .b(new_n235), .c(new_n233), .d(new_n236), .o1(new_n241));
  norb02aa1n02x7               g146(.a(new_n241), .b(new_n240), .out0(\s[24] ));
  nona23aa1n09x5               g147(.a(new_n238), .b(new_n236), .c(new_n235), .d(new_n237), .out0(new_n243));
  inv020aa1n03x5               g148(.a(new_n243), .o1(new_n244));
  nanb03aa1n03x5               g149(.a(new_n210), .b(new_n244), .c(new_n228), .out0(new_n245));
  aoi112aa1n02x5               g150(.a(\b[22] ), .b(\a[23] ), .c(\a[24] ), .d(\b[23] ), .o1(new_n246));
  nanb02aa1n02x5               g151(.a(new_n243), .b(new_n231), .out0(new_n247));
  nona22aa1n02x4               g152(.a(new_n247), .b(new_n246), .c(new_n237), .out0(new_n248));
  aoi013aa1n02x4               g153(.a(new_n248), .b(new_n216), .c(new_n228), .d(new_n244), .o1(new_n249));
  aoai13aa1n04x5               g154(.a(new_n249), .b(new_n245), .c(new_n179), .d(new_n184), .o1(new_n250));
  xorb03aa1n02x5               g155(.a(new_n250), .b(\b[24] ), .c(\a[25] ), .out0(\s[25] ));
  norp02aa1n02x5               g156(.a(\b[24] ), .b(\a[25] ), .o1(new_n252));
  xorc02aa1n02x5               g157(.a(\a[25] ), .b(\b[24] ), .out0(new_n253));
  xorc02aa1n02x5               g158(.a(\a[26] ), .b(\b[25] ), .out0(new_n254));
  aoi112aa1n02x5               g159(.a(new_n252), .b(new_n254), .c(new_n250), .d(new_n253), .o1(new_n255));
  aoai13aa1n03x5               g160(.a(new_n254), .b(new_n252), .c(new_n250), .d(new_n253), .o1(new_n256));
  norb02aa1n02x7               g161(.a(new_n256), .b(new_n255), .out0(\s[26] ));
  nano32aa1d12x5               g162(.a(new_n229), .b(new_n254), .c(new_n244), .d(new_n253), .out0(new_n258));
  nona32aa1n06x5               g163(.a(new_n216), .b(new_n243), .c(new_n223), .d(new_n221), .out0(new_n259));
  aoi112aa1n02x7               g164(.a(new_n246), .b(new_n237), .c(new_n244), .d(new_n231), .o1(new_n260));
  nanp02aa1n02x5               g165(.a(new_n254), .b(new_n253), .o1(new_n261));
  oai022aa1n02x5               g166(.a(\a[25] ), .b(\b[24] ), .c(\b[25] ), .d(\a[26] ), .o1(new_n262));
  aob012aa1n02x5               g167(.a(new_n262), .b(\b[25] ), .c(\a[26] ), .out0(new_n263));
  aoai13aa1n09x5               g168(.a(new_n263), .b(new_n261), .c(new_n259), .d(new_n260), .o1(new_n264));
  xorc02aa1n02x5               g169(.a(\a[27] ), .b(\b[26] ), .out0(new_n265));
  aoai13aa1n06x5               g170(.a(new_n265), .b(new_n264), .c(new_n188), .d(new_n258), .o1(new_n266));
  aoi112aa1n02x5               g171(.a(new_n264), .b(new_n265), .c(new_n188), .d(new_n258), .o1(new_n267));
  norb02aa1n02x5               g172(.a(new_n266), .b(new_n267), .out0(\s[27] ));
  nor042aa1n03x5               g173(.a(\b[26] ), .b(\a[27] ), .o1(new_n269));
  tech160nm_fixorc02aa1n04x5   g174(.a(\a[28] ), .b(\b[27] ), .out0(new_n270));
  nona22aa1n06x5               g175(.a(new_n266), .b(new_n270), .c(new_n269), .out0(new_n271));
  inv000aa1n03x5               g176(.a(new_n269), .o1(new_n272));
  inv000aa1d42x5               g177(.a(new_n270), .o1(new_n273));
  tech160nm_fiaoi012aa1n03p5x5 g178(.a(new_n273), .b(new_n266), .c(new_n272), .o1(new_n274));
  norb02aa1n03x4               g179(.a(new_n271), .b(new_n274), .out0(\s[28] ));
  tech160nm_fixorc02aa1n02p5x5 g180(.a(\a[29] ), .b(\b[28] ), .out0(new_n276));
  inv000aa1d42x5               g181(.a(new_n276), .o1(new_n277));
  and002aa1n02x5               g182(.a(new_n270), .b(new_n265), .o(new_n278));
  aoai13aa1n06x5               g183(.a(new_n278), .b(new_n264), .c(new_n188), .d(new_n258), .o1(new_n279));
  oao003aa1n09x5               g184(.a(\a[28] ), .b(\b[27] ), .c(new_n272), .carry(new_n280));
  aoi012aa1n03x5               g185(.a(new_n277), .b(new_n279), .c(new_n280), .o1(new_n281));
  inv000aa1d42x5               g186(.a(new_n280), .o1(new_n282));
  nona22aa1n02x4               g187(.a(new_n279), .b(new_n282), .c(new_n276), .out0(new_n283));
  norb02aa1n03x4               g188(.a(new_n283), .b(new_n281), .out0(\s[29] ));
  xorb03aa1n02x5               g189(.a(new_n109), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n02x4               g190(.a(new_n277), .b(new_n265), .c(new_n270), .out0(new_n286));
  aoai13aa1n06x5               g191(.a(new_n286), .b(new_n264), .c(new_n188), .d(new_n258), .o1(new_n287));
  oaoi03aa1n02x5               g192(.a(\a[29] ), .b(\b[28] ), .c(new_n280), .o1(new_n288));
  inv000aa1n03x5               g193(.a(new_n288), .o1(new_n289));
  xorc02aa1n02x5               g194(.a(\a[30] ), .b(\b[29] ), .out0(new_n290));
  inv000aa1d42x5               g195(.a(new_n290), .o1(new_n291));
  aoi012aa1n03x5               g196(.a(new_n291), .b(new_n287), .c(new_n289), .o1(new_n292));
  nona22aa1n02x5               g197(.a(new_n287), .b(new_n288), .c(new_n290), .out0(new_n293));
  norb02aa1n02x5               g198(.a(new_n293), .b(new_n292), .out0(\s[30] ));
  nano32aa1n03x7               g199(.a(new_n291), .b(new_n276), .c(new_n270), .d(new_n265), .out0(new_n295));
  aoai13aa1n06x5               g200(.a(new_n295), .b(new_n264), .c(new_n188), .d(new_n258), .o1(new_n296));
  tech160nm_fioaoi03aa1n02p5x5 g201(.a(\a[30] ), .b(\b[29] ), .c(new_n289), .o1(new_n297));
  xorc02aa1n02x5               g202(.a(\a[31] ), .b(\b[30] ), .out0(new_n298));
  nona22aa1n03x5               g203(.a(new_n296), .b(new_n297), .c(new_n298), .out0(new_n299));
  inv000aa1n02x5               g204(.a(new_n297), .o1(new_n300));
  inv000aa1d42x5               g205(.a(new_n298), .o1(new_n301));
  aoi012aa1n06x5               g206(.a(new_n301), .b(new_n296), .c(new_n300), .o1(new_n302));
  norb02aa1n03x4               g207(.a(new_n299), .b(new_n302), .out0(\s[31] ));
  xnbna2aa1n03x5               g208(.a(new_n110), .b(new_n104), .c(new_n105), .out0(\s[3] ));
  xnrc02aa1n02x5               g209(.a(\b[3] ), .b(\a[4] ), .out0(new_n305));
  oai012aa1n02x5               g210(.a(new_n103), .b(new_n110), .c(new_n106), .o1(new_n306));
  oaoi03aa1n02x5               g211(.a(\a[3] ), .b(\b[2] ), .c(new_n110), .o1(new_n307));
  aob012aa1n02x5               g212(.a(new_n306), .b(new_n307), .c(new_n305), .out0(\s[4] ));
  xorb03aa1n02x5               g213(.a(new_n111), .b(\b[4] ), .c(\a[5] ), .out0(\s[5] ));
  nanb02aa1n02x5               g214(.a(new_n114), .b(new_n115), .out0(new_n310));
  aoai13aa1n02x5               g215(.a(new_n310), .b(new_n113), .c(new_n111), .d(new_n112), .o1(new_n311));
  nona23aa1n02x4               g216(.a(new_n306), .b(new_n112), .c(new_n113), .d(new_n99), .out0(new_n312));
  nanp02aa1n02x5               g217(.a(new_n312), .b(new_n116), .o1(new_n313));
  nanp02aa1n02x5               g218(.a(new_n311), .b(new_n313), .o1(\s[6] ));
  aoi022aa1n02x5               g219(.a(new_n312), .b(new_n116), .c(\a[6] ), .d(\b[5] ), .o1(new_n315));
  xorb03aa1n02x5               g220(.a(new_n315), .b(\b[6] ), .c(\a[7] ), .out0(\s[7] ));
  aoi013aa1n02x4               g221(.a(new_n120), .b(new_n313), .c(new_n115), .d(new_n119), .o1(new_n317));
  xnrb03aa1n02x5               g222(.a(new_n317), .b(\b[7] ), .c(\a[8] ), .out0(\s[8] ));
  aoi112aa1n02x5               g223(.a(new_n127), .b(new_n125), .c(new_n111), .d(new_n122), .o1(new_n319));
  norb02aa1n02x5               g224(.a(new_n128), .b(new_n319), .out0(\s[9] ));
endmodule


