// Benchmark "adder" written by ABC on Thu Jul 18 14:48:53 2024

module adder ( 
    \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] , \a[30] ,
    \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] ,
    \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] , \b[23] ,
    \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] , \b[30] ,
    \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] , \s[16] ,
    \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] , \s[23] ,
    \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] , \s[30] ,
    \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] , \s[9]   );
  input  \a[0] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[1] , \a[20] , \a[21] , \a[22] ,
    \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[2] ,
    \a[30] , \a[31] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \b[0] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \b[16] , \b[17] , \b[18] , \b[19] , \b[1] , \b[20] , \b[21] , \b[22] ,
    \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[2] ,
    \b[30] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ;
  output \s[0] , \s[10] , \s[11] , \s[12] , \s[13] , \s[14] , \s[15] ,
    \s[16] , \s[17] , \s[18] , \s[19] , \s[1] , \s[20] , \s[21] , \s[22] ,
    \s[23] , \s[24] , \s[25] , \s[26] , \s[27] , \s[28] , \s[29] , \s[2] ,
    \s[30] , \s[31] , \s[3] , \s[4] , \s[5] , \s[6] , \s[7] , \s[8] ,
    \s[9] ;
  wire new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n201, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n339, new_n341, new_n342, new_n345, new_n346, new_n347,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n355, new_n357,
    new_n358, new_n359;
  inv000aa1d42x5               g000(.a(\a[0] ), .o1(\s[0] ));
  nor002aa1n03x5               g001(.a(\b[1] ), .b(\a[2] ), .o1(new_n97));
  nand42aa1n04x5               g002(.a(\b[1] ), .b(\a[2] ), .o1(new_n98));
  nand22aa1n03x5               g003(.a(\b[0] ), .b(\a[1] ), .o1(new_n99));
  norb03aa1n12x5               g004(.a(new_n98), .b(new_n97), .c(new_n99), .out0(new_n100));
  inv040aa1n02x5               g005(.a(new_n100), .o1(new_n101));
  tech160nm_fioai012aa1n03p5x5 g006(.a(new_n98), .b(\b[3] ), .c(\a[4] ), .o1(new_n102));
  tech160nm_finand02aa1n05x5   g007(.a(\b[2] ), .b(\a[3] ), .o1(new_n103));
  nand02aa1n10x5               g008(.a(\b[3] ), .b(\a[4] ), .o1(new_n104));
  norp02aa1n24x5               g009(.a(\b[2] ), .b(\a[3] ), .o1(new_n105));
  nanb03aa1n02x5               g010(.a(new_n105), .b(new_n103), .c(new_n104), .out0(new_n106));
  nona22aa1n09x5               g011(.a(new_n101), .b(new_n106), .c(new_n102), .out0(new_n107));
  nor042aa1n02x5               g012(.a(\b[3] ), .b(\a[4] ), .o1(new_n108));
  tech160nm_fiaoi012aa1n03p5x5 g013(.a(new_n108), .b(new_n105), .c(new_n104), .o1(new_n109));
  nor042aa1d18x5               g014(.a(\b[6] ), .b(\a[7] ), .o1(new_n110));
  nand42aa1n04x5               g015(.a(\b[6] ), .b(\a[7] ), .o1(new_n111));
  norb02aa1n02x7               g016(.a(new_n111), .b(new_n110), .out0(new_n112));
  tech160nm_fixorc02aa1n03p5x5 g017(.a(\a[5] ), .b(\b[4] ), .out0(new_n113));
  norp02aa1n02x5               g018(.a(\b[5] ), .b(\a[6] ), .o1(new_n114));
  nand02aa1n06x5               g019(.a(\b[5] ), .b(\a[6] ), .o1(new_n115));
  nor022aa1n06x5               g020(.a(\b[7] ), .b(\a[8] ), .o1(new_n116));
  nand02aa1n06x5               g021(.a(\b[7] ), .b(\a[8] ), .o1(new_n117));
  nona23aa1n09x5               g022(.a(new_n117), .b(new_n115), .c(new_n114), .d(new_n116), .out0(new_n118));
  nanb03aa1n03x5               g023(.a(new_n118), .b(new_n112), .c(new_n113), .out0(new_n119));
  tech160nm_fioai012aa1n04x5   g024(.a(new_n117), .b(new_n116), .c(new_n110), .o1(new_n120));
  nanb03aa1n06x5               g025(.a(new_n110), .b(new_n117), .c(new_n111), .out0(new_n121));
  oai022aa1n02x5               g026(.a(\a[5] ), .b(\b[4] ), .c(\b[5] ), .d(\a[6] ), .o1(new_n122));
  oai112aa1n03x5               g027(.a(new_n122), .b(new_n115), .c(\b[7] ), .d(\a[8] ), .o1(new_n123));
  oai012aa1n06x5               g028(.a(new_n120), .b(new_n123), .c(new_n121), .o1(new_n124));
  inv040aa1n03x5               g029(.a(new_n124), .o1(new_n125));
  aoai13aa1n12x5               g030(.a(new_n125), .b(new_n119), .c(new_n107), .d(new_n109), .o1(new_n126));
  nor042aa1n09x5               g031(.a(\b[8] ), .b(\a[9] ), .o1(new_n127));
  nand42aa1n10x5               g032(.a(\b[8] ), .b(\a[9] ), .o1(new_n128));
  norb02aa1n02x5               g033(.a(new_n128), .b(new_n127), .out0(new_n129));
  nor042aa1n04x5               g034(.a(\b[9] ), .b(\a[10] ), .o1(new_n130));
  nand42aa1n08x5               g035(.a(\b[9] ), .b(\a[10] ), .o1(new_n131));
  norb02aa1n02x5               g036(.a(new_n131), .b(new_n130), .out0(new_n132));
  aoi112aa1n02x5               g037(.a(new_n127), .b(new_n132), .c(new_n126), .d(new_n129), .o1(new_n133));
  aoai13aa1n02x5               g038(.a(new_n132), .b(new_n127), .c(new_n126), .d(new_n128), .o1(new_n134));
  norb02aa1n02x5               g039(.a(new_n134), .b(new_n133), .out0(\s[10] ));
  oai012aa1n02x5               g040(.a(new_n131), .b(new_n130), .c(new_n127), .o1(new_n136));
  oai013aa1n03x5               g041(.a(new_n109), .b(new_n100), .c(new_n106), .d(new_n102), .o1(new_n137));
  nano22aa1n03x7               g042(.a(new_n118), .b(new_n113), .c(new_n112), .out0(new_n138));
  nano23aa1d15x5               g043(.a(new_n127), .b(new_n130), .c(new_n131), .d(new_n128), .out0(new_n139));
  aoai13aa1n02x5               g044(.a(new_n139), .b(new_n124), .c(new_n137), .d(new_n138), .o1(new_n140));
  xorc02aa1n12x5               g045(.a(\a[11] ), .b(\b[10] ), .out0(new_n141));
  xnbna2aa1n03x5               g046(.a(new_n141), .b(new_n140), .c(new_n136), .out0(\s[11] ));
  nor042aa1n09x5               g047(.a(\b[10] ), .b(\a[11] ), .o1(new_n143));
  inv000aa1d42x5               g048(.a(new_n143), .o1(new_n144));
  aob012aa1n02x5               g049(.a(new_n141), .b(new_n140), .c(new_n136), .out0(new_n145));
  nor042aa1n02x5               g050(.a(\b[11] ), .b(\a[12] ), .o1(new_n146));
  and002aa1n12x5               g051(.a(\b[11] ), .b(\a[12] ), .o(new_n147));
  nor042aa1n06x5               g052(.a(new_n147), .b(new_n146), .o1(new_n148));
  xnbna2aa1n03x5               g053(.a(new_n148), .b(new_n145), .c(new_n144), .out0(\s[12] ));
  nand23aa1n09x5               g054(.a(new_n139), .b(new_n141), .c(new_n148), .o1(new_n150));
  inv000aa1d42x5               g055(.a(new_n150), .o1(new_n151));
  aoai13aa1n02x5               g056(.a(new_n151), .b(new_n124), .c(new_n137), .d(new_n138), .o1(new_n152));
  aoi112aa1n03x5               g057(.a(new_n147), .b(new_n146), .c(\a[11] ), .d(\b[10] ), .o1(new_n153));
  tech160nm_fioai012aa1n03p5x5 g058(.a(new_n131), .b(\b[10] ), .c(\a[11] ), .o1(new_n154));
  oab012aa1n06x5               g059(.a(new_n154), .b(new_n127), .c(new_n130), .out0(new_n155));
  oaoi03aa1n12x5               g060(.a(\a[12] ), .b(\b[11] ), .c(new_n144), .o1(new_n156));
  aoi012aa1n02x5               g061(.a(new_n156), .b(new_n155), .c(new_n153), .o1(new_n157));
  nanp02aa1n03x5               g062(.a(new_n152), .b(new_n157), .o1(new_n158));
  nor042aa1n04x5               g063(.a(\b[12] ), .b(\a[13] ), .o1(new_n159));
  nand02aa1n06x5               g064(.a(\b[12] ), .b(\a[13] ), .o1(new_n160));
  norb02aa1n02x5               g065(.a(new_n160), .b(new_n159), .out0(new_n161));
  aoi112aa1n02x5               g066(.a(new_n156), .b(new_n161), .c(new_n155), .d(new_n153), .o1(new_n162));
  aoi022aa1n02x5               g067(.a(new_n158), .b(new_n161), .c(new_n152), .d(new_n162), .o1(\s[13] ));
  nor042aa1n04x5               g068(.a(\b[13] ), .b(\a[14] ), .o1(new_n164));
  nand42aa1n06x5               g069(.a(\b[13] ), .b(\a[14] ), .o1(new_n165));
  norb02aa1n02x5               g070(.a(new_n165), .b(new_n164), .out0(new_n166));
  aoi112aa1n02x5               g071(.a(new_n159), .b(new_n166), .c(new_n158), .d(new_n161), .o1(new_n167));
  aoai13aa1n02x5               g072(.a(new_n166), .b(new_n159), .c(new_n158), .d(new_n160), .o1(new_n168));
  norb02aa1n02x5               g073(.a(new_n168), .b(new_n167), .out0(\s[14] ));
  inv000aa1n02x5               g074(.a(new_n157), .o1(new_n170));
  nano23aa1d15x5               g075(.a(new_n159), .b(new_n164), .c(new_n165), .d(new_n160), .out0(new_n171));
  aoai13aa1n06x5               g076(.a(new_n171), .b(new_n170), .c(new_n126), .d(new_n151), .o1(new_n172));
  oai012aa1n18x5               g077(.a(new_n165), .b(new_n164), .c(new_n159), .o1(new_n173));
  xorc02aa1n12x5               g078(.a(\a[15] ), .b(\b[14] ), .out0(new_n174));
  xnbna2aa1n03x5               g079(.a(new_n174), .b(new_n172), .c(new_n173), .out0(\s[15] ));
  inv000aa1d42x5               g080(.a(new_n173), .o1(new_n176));
  aoai13aa1n03x5               g081(.a(new_n174), .b(new_n176), .c(new_n158), .d(new_n171), .o1(new_n177));
  tech160nm_fixorc02aa1n03p5x5 g082(.a(\a[16] ), .b(\b[15] ), .out0(new_n178));
  nor042aa1n06x5               g083(.a(\b[14] ), .b(\a[15] ), .o1(new_n179));
  norp02aa1n02x5               g084(.a(new_n178), .b(new_n179), .o1(new_n180));
  inv000aa1d42x5               g085(.a(new_n179), .o1(new_n181));
  inv000aa1d42x5               g086(.a(new_n174), .o1(new_n182));
  aoai13aa1n03x5               g087(.a(new_n181), .b(new_n182), .c(new_n172), .d(new_n173), .o1(new_n183));
  aoi022aa1n02x5               g088(.a(new_n183), .b(new_n178), .c(new_n177), .d(new_n180), .o1(\s[16] ));
  nano32aa1d12x5               g089(.a(new_n150), .b(new_n178), .c(new_n171), .d(new_n174), .out0(new_n185));
  nanp02aa1n02x5               g090(.a(new_n178), .b(new_n174), .o1(new_n186));
  aoai13aa1n06x5               g091(.a(new_n171), .b(new_n156), .c(new_n155), .d(new_n153), .o1(new_n187));
  oao003aa1n02x5               g092(.a(\a[16] ), .b(\b[15] ), .c(new_n181), .carry(new_n188));
  aoai13aa1n12x5               g093(.a(new_n188), .b(new_n186), .c(new_n187), .d(new_n173), .o1(new_n189));
  xorc02aa1n02x5               g094(.a(\a[17] ), .b(\b[16] ), .out0(new_n190));
  aoai13aa1n06x5               g095(.a(new_n190), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n191));
  aoai13aa1n06x5               g096(.a(new_n185), .b(new_n124), .c(new_n137), .d(new_n138), .o1(new_n192));
  and002aa1n02x5               g097(.a(new_n178), .b(new_n174), .o(new_n193));
  aob012aa1n06x5               g098(.a(new_n193), .b(new_n187), .c(new_n173), .out0(new_n194));
  nano32aa1n02x4               g099(.a(new_n190), .b(new_n194), .c(new_n192), .d(new_n188), .out0(new_n195));
  norb02aa1n02x5               g100(.a(new_n191), .b(new_n195), .out0(\s[17] ));
  nor002aa1d32x5               g101(.a(\b[16] ), .b(\a[17] ), .o1(new_n197));
  inv000aa1d42x5               g102(.a(new_n197), .o1(new_n198));
  nor042aa1n06x5               g103(.a(\b[17] ), .b(\a[18] ), .o1(new_n199));
  nand02aa1n08x5               g104(.a(\b[17] ), .b(\a[18] ), .o1(new_n200));
  norb02aa1n03x5               g105(.a(new_n200), .b(new_n199), .out0(new_n201));
  xnbna2aa1n03x5               g106(.a(new_n201), .b(new_n191), .c(new_n198), .out0(\s[18] ));
  and002aa1n02x5               g107(.a(new_n190), .b(new_n201), .o(new_n203));
  aoai13aa1n03x5               g108(.a(new_n203), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n204));
  oaoi03aa1n02x5               g109(.a(\a[18] ), .b(\b[17] ), .c(new_n198), .o1(new_n205));
  inv000aa1d42x5               g110(.a(new_n205), .o1(new_n206));
  nor002aa1d32x5               g111(.a(\b[18] ), .b(\a[19] ), .o1(new_n207));
  nand02aa1n04x5               g112(.a(\b[18] ), .b(\a[19] ), .o1(new_n208));
  norb02aa1n12x5               g113(.a(new_n208), .b(new_n207), .out0(new_n209));
  xnbna2aa1n03x5               g114(.a(new_n209), .b(new_n204), .c(new_n206), .out0(\s[19] ));
  xnrc02aa1n02x5               g115(.a(\b[0] ), .b(\a[1] ), .out0(\s[1] ));
  nanp03aa1d12x5               g116(.a(new_n194), .b(new_n192), .c(new_n188), .o1(new_n212));
  aoai13aa1n03x5               g117(.a(new_n209), .b(new_n205), .c(new_n212), .d(new_n203), .o1(new_n213));
  nor002aa1n12x5               g118(.a(\b[19] ), .b(\a[20] ), .o1(new_n214));
  nand02aa1d24x5               g119(.a(\b[19] ), .b(\a[20] ), .o1(new_n215));
  norb02aa1n02x5               g120(.a(new_n215), .b(new_n214), .out0(new_n216));
  inv000aa1d42x5               g121(.a(\a[19] ), .o1(new_n217));
  inv000aa1d42x5               g122(.a(\b[18] ), .o1(new_n218));
  aboi22aa1n03x5               g123(.a(new_n214), .b(new_n215), .c(new_n217), .d(new_n218), .out0(new_n219));
  inv000aa1d42x5               g124(.a(new_n207), .o1(new_n220));
  inv000aa1d42x5               g125(.a(new_n209), .o1(new_n221));
  aoai13aa1n02x5               g126(.a(new_n220), .b(new_n221), .c(new_n204), .d(new_n206), .o1(new_n222));
  aoi022aa1n03x5               g127(.a(new_n222), .b(new_n216), .c(new_n213), .d(new_n219), .o1(\s[20] ));
  nano32aa1n03x7               g128(.a(new_n221), .b(new_n190), .c(new_n216), .d(new_n201), .out0(new_n224));
  aoai13aa1n03x5               g129(.a(new_n224), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n225));
  nanb03aa1n12x5               g130(.a(new_n214), .b(new_n215), .c(new_n208), .out0(new_n226));
  oai112aa1n06x5               g131(.a(new_n220), .b(new_n200), .c(new_n199), .d(new_n197), .o1(new_n227));
  aoi012aa1d18x5               g132(.a(new_n214), .b(new_n207), .c(new_n215), .o1(new_n228));
  oai012aa1d24x5               g133(.a(new_n228), .b(new_n227), .c(new_n226), .o1(new_n229));
  nor002aa1d32x5               g134(.a(\b[20] ), .b(\a[21] ), .o1(new_n230));
  nand02aa1n06x5               g135(.a(\b[20] ), .b(\a[21] ), .o1(new_n231));
  norb02aa1n15x5               g136(.a(new_n231), .b(new_n230), .out0(new_n232));
  aoai13aa1n06x5               g137(.a(new_n232), .b(new_n229), .c(new_n212), .d(new_n224), .o1(new_n233));
  nano22aa1n03x7               g138(.a(new_n214), .b(new_n208), .c(new_n215), .out0(new_n234));
  tech160nm_fioai012aa1n04x5   g139(.a(new_n200), .b(\b[18] ), .c(\a[19] ), .o1(new_n235));
  oab012aa1n02x5               g140(.a(new_n235), .b(new_n197), .c(new_n199), .out0(new_n236));
  inv020aa1n02x5               g141(.a(new_n228), .o1(new_n237));
  aoi112aa1n02x5               g142(.a(new_n237), .b(new_n232), .c(new_n236), .d(new_n234), .o1(new_n238));
  aobi12aa1n03x7               g143(.a(new_n233), .b(new_n238), .c(new_n225), .out0(\s[21] ));
  nor042aa1n04x5               g144(.a(\b[21] ), .b(\a[22] ), .o1(new_n240));
  nanp02aa1n12x5               g145(.a(\b[21] ), .b(\a[22] ), .o1(new_n241));
  norb02aa1n02x5               g146(.a(new_n241), .b(new_n240), .out0(new_n242));
  aoib12aa1n02x5               g147(.a(new_n230), .b(new_n241), .c(new_n240), .out0(new_n243));
  inv000aa1d42x5               g148(.a(new_n229), .o1(new_n244));
  inv000aa1d42x5               g149(.a(new_n230), .o1(new_n245));
  inv000aa1d42x5               g150(.a(new_n232), .o1(new_n246));
  aoai13aa1n03x5               g151(.a(new_n245), .b(new_n246), .c(new_n225), .d(new_n244), .o1(new_n247));
  aoi022aa1n03x5               g152(.a(new_n247), .b(new_n242), .c(new_n233), .d(new_n243), .o1(\s[22] ));
  inv000aa1n02x5               g153(.a(new_n224), .o1(new_n249));
  nano22aa1n02x5               g154(.a(new_n249), .b(new_n232), .c(new_n242), .out0(new_n250));
  aoai13aa1n03x5               g155(.a(new_n250), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n251));
  nano23aa1d12x5               g156(.a(new_n230), .b(new_n240), .c(new_n241), .d(new_n231), .out0(new_n252));
  aoi012aa1d18x5               g157(.a(new_n240), .b(new_n230), .c(new_n241), .o1(new_n253));
  inv000aa1n02x5               g158(.a(new_n253), .o1(new_n254));
  aoi012aa1n02x5               g159(.a(new_n254), .b(new_n229), .c(new_n252), .o1(new_n255));
  inv040aa1n03x5               g160(.a(new_n255), .o1(new_n256));
  xorc02aa1n12x5               g161(.a(\a[23] ), .b(\b[22] ), .out0(new_n257));
  aoai13aa1n06x5               g162(.a(new_n257), .b(new_n256), .c(new_n212), .d(new_n250), .o1(new_n258));
  aoi112aa1n02x5               g163(.a(new_n257), .b(new_n254), .c(new_n229), .d(new_n252), .o1(new_n259));
  aobi12aa1n02x7               g164(.a(new_n258), .b(new_n259), .c(new_n251), .out0(\s[23] ));
  tech160nm_fixorc02aa1n02p5x5 g165(.a(\a[24] ), .b(\b[23] ), .out0(new_n261));
  nor042aa1n06x5               g166(.a(\b[22] ), .b(\a[23] ), .o1(new_n262));
  norp02aa1n02x5               g167(.a(new_n261), .b(new_n262), .o1(new_n263));
  inv000aa1d42x5               g168(.a(new_n262), .o1(new_n264));
  inv000aa1d42x5               g169(.a(new_n257), .o1(new_n265));
  aoai13aa1n03x5               g170(.a(new_n264), .b(new_n265), .c(new_n251), .d(new_n255), .o1(new_n266));
  aoi022aa1n03x5               g171(.a(new_n266), .b(new_n261), .c(new_n258), .d(new_n263), .o1(\s[24] ));
  and002aa1n12x5               g172(.a(new_n261), .b(new_n257), .o(new_n268));
  nano22aa1n02x5               g173(.a(new_n249), .b(new_n268), .c(new_n252), .out0(new_n269));
  aoai13aa1n06x5               g174(.a(new_n269), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n270));
  aoai13aa1n04x5               g175(.a(new_n252), .b(new_n237), .c(new_n236), .d(new_n234), .o1(new_n271));
  inv000aa1n06x5               g176(.a(new_n268), .o1(new_n272));
  oao003aa1n02x5               g177(.a(\a[24] ), .b(\b[23] ), .c(new_n264), .carry(new_n273));
  aoai13aa1n12x5               g178(.a(new_n273), .b(new_n272), .c(new_n271), .d(new_n253), .o1(new_n274));
  xorc02aa1n12x5               g179(.a(\a[25] ), .b(\b[24] ), .out0(new_n275));
  aoai13aa1n06x5               g180(.a(new_n275), .b(new_n274), .c(new_n212), .d(new_n269), .o1(new_n276));
  aoai13aa1n06x5               g181(.a(new_n268), .b(new_n254), .c(new_n229), .d(new_n252), .o1(new_n277));
  inv000aa1d42x5               g182(.a(new_n275), .o1(new_n278));
  and003aa1n02x5               g183(.a(new_n277), .b(new_n278), .c(new_n273), .o(new_n279));
  aobi12aa1n03x7               g184(.a(new_n276), .b(new_n279), .c(new_n270), .out0(\s[25] ));
  tech160nm_fixorc02aa1n02p5x5 g185(.a(\a[26] ), .b(\b[25] ), .out0(new_n281));
  nor042aa1n03x5               g186(.a(\b[24] ), .b(\a[25] ), .o1(new_n282));
  norp02aa1n02x5               g187(.a(new_n281), .b(new_n282), .o1(new_n283));
  inv000aa1d42x5               g188(.a(new_n274), .o1(new_n284));
  inv000aa1d42x5               g189(.a(new_n282), .o1(new_n285));
  aoai13aa1n03x5               g190(.a(new_n285), .b(new_n278), .c(new_n270), .d(new_n284), .o1(new_n286));
  aoi022aa1n03x5               g191(.a(new_n286), .b(new_n281), .c(new_n276), .d(new_n283), .o1(\s[26] ));
  and002aa1n12x5               g192(.a(new_n281), .b(new_n275), .o(new_n288));
  nano32aa1n03x7               g193(.a(new_n249), .b(new_n288), .c(new_n252), .d(new_n268), .out0(new_n289));
  aoai13aa1n06x5               g194(.a(new_n289), .b(new_n189), .c(new_n126), .d(new_n185), .o1(new_n290));
  inv000aa1d42x5               g195(.a(new_n288), .o1(new_n291));
  oao003aa1n02x5               g196(.a(\a[26] ), .b(\b[25] ), .c(new_n285), .carry(new_n292));
  aoai13aa1n04x5               g197(.a(new_n292), .b(new_n291), .c(new_n277), .d(new_n273), .o1(new_n293));
  xorc02aa1n12x5               g198(.a(\a[27] ), .b(\b[26] ), .out0(new_n294));
  aoai13aa1n06x5               g199(.a(new_n294), .b(new_n293), .c(new_n212), .d(new_n289), .o1(new_n295));
  inv000aa1d42x5               g200(.a(new_n292), .o1(new_n296));
  aoi112aa1n02x5               g201(.a(new_n294), .b(new_n296), .c(new_n274), .d(new_n288), .o1(new_n297));
  aobi12aa1n02x7               g202(.a(new_n295), .b(new_n297), .c(new_n290), .out0(\s[27] ));
  tech160nm_fixorc02aa1n02p5x5 g203(.a(\a[28] ), .b(\b[27] ), .out0(new_n299));
  norp02aa1n02x5               g204(.a(\b[26] ), .b(\a[27] ), .o1(new_n300));
  norp02aa1n02x5               g205(.a(new_n299), .b(new_n300), .o1(new_n301));
  aoi012aa1n09x5               g206(.a(new_n296), .b(new_n274), .c(new_n288), .o1(new_n302));
  inv000aa1n03x5               g207(.a(new_n300), .o1(new_n303));
  inv000aa1d42x5               g208(.a(new_n294), .o1(new_n304));
  aoai13aa1n03x5               g209(.a(new_n303), .b(new_n304), .c(new_n290), .d(new_n302), .o1(new_n305));
  aoi022aa1n03x5               g210(.a(new_n305), .b(new_n299), .c(new_n295), .d(new_n301), .o1(\s[28] ));
  and002aa1n02x5               g211(.a(new_n299), .b(new_n294), .o(new_n307));
  aoai13aa1n03x5               g212(.a(new_n307), .b(new_n293), .c(new_n212), .d(new_n289), .o1(new_n308));
  xorc02aa1n02x5               g213(.a(\a[29] ), .b(\b[28] ), .out0(new_n309));
  oao003aa1n02x5               g214(.a(\a[28] ), .b(\b[27] ), .c(new_n303), .carry(new_n310));
  norb02aa1n02x5               g215(.a(new_n310), .b(new_n309), .out0(new_n311));
  inv000aa1d42x5               g216(.a(new_n307), .o1(new_n312));
  aoai13aa1n03x5               g217(.a(new_n310), .b(new_n312), .c(new_n290), .d(new_n302), .o1(new_n313));
  aoi022aa1n03x5               g218(.a(new_n313), .b(new_n309), .c(new_n308), .d(new_n311), .o1(\s[29] ));
  xorb03aa1n02x5               g219(.a(new_n99), .b(\b[1] ), .c(\a[2] ), .out0(\s[2] ));
  nano22aa1n06x5               g220(.a(new_n304), .b(new_n299), .c(new_n309), .out0(new_n316));
  aoai13aa1n03x5               g221(.a(new_n316), .b(new_n293), .c(new_n212), .d(new_n289), .o1(new_n317));
  xorc02aa1n02x5               g222(.a(\a[30] ), .b(\b[29] ), .out0(new_n318));
  inv000aa1d42x5               g223(.a(\a[29] ), .o1(new_n319));
  inv000aa1d42x5               g224(.a(\b[28] ), .o1(new_n320));
  oaib12aa1n02x5               g225(.a(new_n310), .b(\b[28] ), .c(new_n319), .out0(new_n321));
  oaoi13aa1n02x5               g226(.a(new_n318), .b(new_n321), .c(new_n319), .d(new_n320), .o1(new_n322));
  inv000aa1d42x5               g227(.a(new_n316), .o1(new_n323));
  oaib12aa1n02x5               g228(.a(new_n321), .b(new_n320), .c(\a[29] ), .out0(new_n324));
  aoai13aa1n03x5               g229(.a(new_n324), .b(new_n323), .c(new_n290), .d(new_n302), .o1(new_n325));
  aoi022aa1n03x5               g230(.a(new_n325), .b(new_n318), .c(new_n317), .d(new_n322), .o1(\s[30] ));
  nano32aa1n06x5               g231(.a(new_n304), .b(new_n318), .c(new_n299), .d(new_n309), .out0(new_n327));
  aoai13aa1n02x5               g232(.a(new_n327), .b(new_n293), .c(new_n212), .d(new_n289), .o1(new_n328));
  aoi022aa1n02x5               g233(.a(\b[29] ), .b(\a[30] ), .c(\a[29] ), .d(\b[28] ), .o1(new_n329));
  norb02aa1n02x5               g234(.a(\b[30] ), .b(\a[31] ), .out0(new_n330));
  obai22aa1n02x7               g235(.a(\a[31] ), .b(\b[30] ), .c(\a[30] ), .d(\b[29] ), .out0(new_n331));
  aoi112aa1n02x5               g236(.a(new_n331), .b(new_n330), .c(new_n321), .d(new_n329), .o1(new_n332));
  xorc02aa1n02x5               g237(.a(\a[31] ), .b(\b[30] ), .out0(new_n333));
  inv000aa1d42x5               g238(.a(new_n327), .o1(new_n334));
  norp02aa1n02x5               g239(.a(\b[29] ), .b(\a[30] ), .o1(new_n335));
  aoi012aa1n02x5               g240(.a(new_n335), .b(new_n321), .c(new_n329), .o1(new_n336));
  aoai13aa1n03x5               g241(.a(new_n336), .b(new_n334), .c(new_n290), .d(new_n302), .o1(new_n337));
  aoi022aa1n03x5               g242(.a(new_n337), .b(new_n333), .c(new_n328), .d(new_n332), .o1(\s[31] ));
  norb02aa1n02x5               g243(.a(new_n103), .b(new_n105), .out0(new_n339));
  xobna2aa1n03x5               g244(.a(new_n339), .b(new_n101), .c(new_n98), .out0(\s[3] ));
  aoai13aa1n02x5               g245(.a(new_n339), .b(new_n100), .c(\a[2] ), .d(\b[1] ), .o1(new_n341));
  nanb02aa1n02x5               g246(.a(new_n108), .b(new_n104), .out0(new_n342));
  xnbna2aa1n03x5               g247(.a(new_n342), .b(new_n341), .c(new_n103), .out0(\s[4] ));
  xnbna2aa1n03x5               g248(.a(new_n113), .b(new_n107), .c(new_n109), .out0(\s[5] ));
  orn002aa1n02x5               g249(.a(\a[5] ), .b(\b[4] ), .o(new_n345));
  norb02aa1n02x5               g250(.a(new_n115), .b(new_n114), .out0(new_n346));
  nanp02aa1n02x5               g251(.a(new_n137), .b(new_n113), .o1(new_n347));
  xnbna2aa1n03x5               g252(.a(new_n346), .b(new_n347), .c(new_n345), .out0(\s[6] ));
  nanp03aa1n02x5               g253(.a(new_n347), .b(new_n345), .c(new_n346), .o1(new_n349));
  nano22aa1n02x4               g254(.a(new_n110), .b(new_n111), .c(new_n115), .out0(new_n350));
  nanp02aa1n02x5               g255(.a(new_n349), .b(new_n350), .o1(new_n351));
  inv000aa1d42x5               g256(.a(new_n110), .o1(new_n352));
  aoi022aa1n02x5               g257(.a(new_n349), .b(new_n115), .c(new_n352), .d(new_n111), .o1(new_n353));
  norb02aa1n02x5               g258(.a(new_n351), .b(new_n353), .out0(\s[7] ));
  norb02aa1n02x5               g259(.a(new_n117), .b(new_n116), .out0(new_n355));
  xnbna2aa1n03x5               g260(.a(new_n355), .b(new_n351), .c(new_n352), .out0(\s[8] ));
  nanp02aa1n02x5               g261(.a(new_n137), .b(new_n138), .o1(new_n357));
  oaib12aa1n02x5               g262(.a(new_n120), .b(new_n127), .c(new_n128), .out0(new_n358));
  oab012aa1n02x4               g263(.a(new_n358), .b(new_n123), .c(new_n121), .out0(new_n359));
  aoi022aa1n02x5               g264(.a(new_n126), .b(new_n129), .c(new_n357), .d(new_n359), .o1(\s[9] ));
endmodule


